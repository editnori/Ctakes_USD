 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|158,166|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Pharmacologic Substance|Allergies|181,186|false|false|false|C0749139|sulfa|Sulfa
Event|Event|Allergies|181,186|false|false|false|||Sulfa
Drug|Antibiotic|Allergies|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Organic Chemical|Allergies|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Pharmacologic Substance|Allergies|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Antibiotic|Allergies|200,211|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|Allergies|200,211|false|false|false|||Antibiotics
Drug|Organic Chemical|Allergies|215,222|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|215,222|false|false|false|C0009214|codeine|Codeine
Drug|Organic Chemical|Allergies|225,232|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|Allergies|225,232|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|Allergies|235,244|false|false|false|||Attending
Finding|Functional Concept|Allergies|235,244|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|270,279|false|false|false|||Shortness
Attribute|Clinical Attribute|Chief Complaint|270,289|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Chief Complaint|270,289|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Chief Complaint|283,289|false|false|false|C0225386|Breath|breath
Finding|Classification|Chief Complaint|292,297|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|298,306|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,306|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|310,328|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|319,328|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|319,328|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|319,328|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|319,328|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|319,328|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|330,342|false|false|false|C1522243|Percutaneous Route of Drug Administration|Percutaneous
Procedure|Diagnostic Procedure|Chief Complaint|330,355|false|false|false|C0558534|Percutaneous liver biopsy|Percutaneous liver biopsy
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|343,348|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Chief Complaint|343,348|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Chief Complaint|343,348|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Chief Complaint|343,348|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Chief Complaint|343,348|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Chief Complaint|343,348|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Chief Complaint|343,348|false|false|false|||liver
Finding|Finding|Chief Complaint|343,348|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Chief Complaint|343,348|false|false|false|C0872387|Procedures on liver|liver
Procedure|Diagnostic Procedure|Chief Complaint|343,355|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Procedure|Health Care Activity|Chief Complaint|343,355|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Event|Event|Chief Complaint|349,355|false|false|false|||biopsy
Finding|Finding|Chief Complaint|349,355|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Chief Complaint|349,355|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Chief Complaint|349,355|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Chief Complaint|349,355|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Finding|Functional Concept|History of Present Illness|408,418|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|History of Present Illness|408,425|false|false|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|History of Present Illness|419,425|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|419,425|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|429,436|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|History of Present Illness|429,436|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|History of Present Illness|429,436|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|History of Present Illness|429,436|false|false|false|||unknown
Finding|Finding|History of Present Illness|429,436|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|History of Present Illness|429,436|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|History of Present Illness|429,436|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|History of Present Illness|429,436|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|History of Present Illness|453,460|false|false|false|||lesions
Finding|Finding|History of Present Illness|453,460|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|464,469|false|false|false|C0024109|Lung|lungs
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|474,479|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|History of Present Illness|474,479|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|History of Present Illness|474,479|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|History of Present Illness|474,479|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|History of Present Illness|474,479|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|History of Present Illness|474,479|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|History of Present Illness|474,479|false|false|false|||liver
Finding|Finding|History of Present Illness|474,479|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|History of Present Illness|474,479|false|false|false|C0872387|Procedures on liver|liver
Event|Event|History of Present Illness|481,491|false|false|false|||presenting
Event|Event|History of Present Illness|497,506|false|false|false|||shortness
Event|Event|History of Present Illness|511,517|false|false|false|||breath
Finding|Body Substance|History of Present Illness|511,517|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|533,542|false|false|false|||presented
Anatomy|Body Location or Region|History of Present Illness|562,571|false|false|false|C0000726|Abdomen|abdominal
Attribute|Clinical Attribute|History of Present Illness|573,577|false|false|false|C2598155||pain
Event|Event|History of Present Illness|573,577|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|573,577|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|573,577|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|582,589|false|false|false|||failure
Finding|Functional Concept|History of Present Illness|582,589|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|582,589|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|582,589|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|History of Present Illness|593,599|false|false|false|||thrive
Event|Event|History of Present Illness|601,611|false|false|false|||Evaluation
Finding|Idea or Concept|History of Present Illness|601,611|false|false|false|C1550157|Processing type - Evaluation|Evaluation
Procedure|Health Care Activity|History of Present Illness|601,611|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|Evaluation
Finding|Finding|History of Present Illness|620,624|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|620,624|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|620,624|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|History of Present Illness|638,647|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|History of Present Illness|638,655|false|false|false|C0412620|CT of abdomen|abdominal CT scan
Procedure|Diagnostic Procedure|History of Present Illness|648,655|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|History of Present Illness|651,655|false|false|false|||scan
Procedure|Diagnostic Procedure|History of Present Illness|651,655|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|History of Present Illness|661,667|false|false|false|||showed
Anatomy|Body Location or Region|History of Present Illness|677,681|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|677,681|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|History of Present Illness|677,681|false|false|false|C0024115|Lung diseases|lung
Event|Event|History of Present Illness|677,681|false|false|false|||lung
Finding|Finding|History of Present Illness|677,681|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Location or Region|History of Present Illness|677,691|false|false|false|C4266618|Lung and Liver|lung and liver
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|686,691|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|History of Present Illness|686,691|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|History of Present Illness|686,691|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|History of Present Illness|686,691|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|History of Present Illness|686,691|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|History of Present Illness|686,691|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|History of Present Illness|686,691|false|false|false|||liver
Finding|Finding|History of Present Illness|686,691|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|History of Present Illness|686,691|false|false|false|C0872387|Procedures on liver|liver
Disorder|Neoplastic Process|History of Present Illness|693,703|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|History of Present Illness|693,703|false|false|false|||metastases
Finding|Finding|History of Present Illness|693,703|false|false|false|C1513183|Metastatic Lesion|metastases
Attribute|Clinical Attribute|History of Present Illness|737,746|false|false|false|C0945731||diagnosis
Event|Event|History of Present Illness|737,746|false|false|false|||diagnosis
Finding|Classification|History of Present Illness|737,746|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|History of Present Illness|737,746|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|737,746|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|History of Present Illness|753,759|false|false|false|||biopsy
Finding|Finding|History of Present Illness|753,759|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|History of Present Illness|753,759|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|History of Present Illness|753,759|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|History of Present Illness|753,759|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Neoplastic Process|History of Present Illness|776,784|false|false|false|C0027651|Neoplasms|oncology
Event|Event|History of Present Illness|776,784|false|false|false|||oncology
Procedure|Health Care Activity|History of Present Illness|776,784|false|false|false|C1555459|oncology services|oncology
Event|Event|History of Present Illness|785,798|false|false|false|||documentation
Finding|Intellectual Product|History of Present Illness|785,798|false|false|false|C0920316|Documentation|documentation
Procedure|Health Care Activity|History of Present Illness|785,798|false|false|false|C0175636|Act of Documentation|documentation
Event|Event|History of Present Illness|805,815|false|false|false|||disengaged
Event|Activity|History of Present Illness|822,826|false|false|false|C1947933|care activity|care
Event|Event|History of Present Illness|822,826|false|false|false|||care
Finding|Finding|History of Present Illness|822,826|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|822,826|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|History of Present Illness|862,867|false|false|false|||state
Finding|Functional Concept|History of Present Illness|862,867|false|false|false|C1442792|State|state
Finding|Finding|History of Present Illness|862,877|false|false|false|C0683314|personal health|state of health
Event|Event|History of Present Illness|871,877|false|false|false|||health
Finding|Idea or Concept|History of Present Illness|871,877|false|false|false|C0018684|Health|health
Event|Event|History of Present Illness|906,915|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|906,915|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|926,935|false|false|false|||developed
Event|Event|History of Present Illness|936,941|false|false|false|||acute
Finding|Intellectual Product|History of Present Illness|936,941|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|945,952|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|945,952|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|945,952|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|History of Present Illness|954,963|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|954,973|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|954,973|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|History of Present Illness|967,973|false|false|false|||breath
Finding|Body Substance|History of Present Illness|967,973|false|false|false|C0225386|Breath|breath
Finding|Functional Concept|History of Present Illness|980,987|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|983,987|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|983,987|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|History of Present Illness|983,987|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|983,987|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|983,987|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|History of Present Illness|993,1001|false|false|false|||reported
Anatomy|Body Location or Region|History of Present Illness|1013,1018|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1013,1018|false|false|false|C0741025|Chest problem|chest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1020,1024|false|false|false|C0001044;C2932864|ACHE protein, human;acetylcholinesterase|ache
Drug|Enzyme|History of Present Illness|1020,1024|false|false|false|C0001044;C2932864|ACHE protein, human;acetylcholinesterase|ache
Event|Event|History of Present Illness|1020,1024|false|false|false|||ache
Finding|Gene or Genome|History of Present Illness|1020,1024|false|false|false|C0030193;C0234238;C1412122|ACHE Gene;Ache;Pain|ache
Finding|Sign or Symptom|History of Present Illness|1020,1024|false|false|false|C0030193;C0234238;C1412122|ACHE Gene;Ache;Pain|ache
Event|Event|History of Present Illness|1046,1055|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|1046,1065|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1046,1065|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1059,1065|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|History of Present Illness|1067,1071|false|false|false|C2598155||Pain
Finding|Functional Concept|History of Present Illness|1067,1071|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|History of Present Illness|1067,1071|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|History of Present Illness|1076,1087|false|false|false|||exacerbated
Finding|Intellectual Product|History of Present Illness|1091,1097|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|direct
Event|Event|History of Present Illness|1098,1106|false|false|false|||pressure
Finding|Finding|History of Present Illness|1098,1106|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|1098,1106|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|1098,1106|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|1098,1106|false|false|false|C0033095||pressure
Event|Event|History of Present Illness|1108,1115|false|false|false|||nothing
Attribute|Clinical Attribute|History of Present Illness|1135,1139|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1135,1139|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1135,1139|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1135,1139|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1146,1152|true|false|false|||denied
Event|Event|History of Present Illness|1170,1180|true|false|false|||exertional
Finding|Sign or Symptom|History of Present Illness|1170,1180|true|false|false|C0239313|exercise induced|exertional
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1181,1190|true|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|History of Present Illness|1181,1190|true|false|false|C1179435|Protein Component|component
Event|Event|History of Present Illness|1181,1190|true|false|false|||component
Finding|Conceptual Entity|History of Present Illness|1181,1190|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|History of Present Illness|1181,1190|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|History of Present Illness|1181,1190|true|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Anatomy|Body Location or Region|History of Present Illness|1198,1203|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1198,1203|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1205,1209|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1205,1209|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1205,1209|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1205,1209|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1213,1222|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|1213,1232|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1213,1232|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1226,1232|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1238,1243|false|false|false|||feels
Event|Event|History of Present Illness|1249,1257|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1249,1257|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1249,1257|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Neoplastic Process|History of Present Illness|1263,1272|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|History of Present Illness|1263,1272|false|false|false|||secondary
Finding|Functional Concept|History of Present Illness|1263,1272|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Neoplastic Process|History of Present Illness|1281,1287|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|1281,1287|false|false|false|||cancer
Event|Event|History of Present Illness|1294,1299|false|false|false|||feels
Disorder|Neoplastic Process|History of Present Illness|1310,1316|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|1310,1316|false|false|false|||cancer
Event|Activity|History of Present Illness|1322,1328|false|false|false|C1947932|Smear - instruction imperative|spread
Event|Event|History of Present Illness|1322,1328|false|false|false|||spread
Event|Event|History of Present Illness|1335,1342|false|false|false|||reports
Event|Event|History of Present Illness|1343,1349|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1343,1349|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|History of Present Illness|1351,1358|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|1351,1358|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|1351,1358|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Organic Chemical|History of Present Illness|1373,1378|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1373,1378|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1373,1378|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1373,1378|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1396,1403|false|false|false|||present
Finding|Finding|History of Present Illness|1396,1403|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|History of Present Illness|1396,1403|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|History of Present Illness|1441,1445|false|false|false|||seen
Event|Event|History of Present Illness|1469,1479|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|1469,1479|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|1469,1479|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Functional Concept|History of Present Illness|1483,1487|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|History of Present Illness|1502,1507|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1502,1523|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|1508,1513|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|1508,1513|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1508,1523|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|History of Present Illness|1508,1529|false|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1514,1523|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|History of Present Illness|1514,1529|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|History of Present Illness|1524,1529|false|true|false|C1717255||edema
Event|Event|History of Present Illness|1524,1529|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|1524,1529|false|true|false|C0013604|Edema|edema
Anatomy|Body Location or Region|History of Present Illness|1535,1540|true|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|1535,1540|true|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1535,1550|true|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1541,1550|true|false|false|C0015385|Limb structure|extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1551,1557|true|false|false|C0042449|Veins|venous
Event|Event|History of Present Illness|1559,1570|true|false|false|||ultrasounds
Procedure|Diagnostic Procedure|History of Present Illness|1559,1570|true|false|false|C0041618|Ultrasonography|ultrasounds
Event|Event|History of Present Illness|1571,1579|true|false|false|||negative
Finding|Classification|History of Present Illness|1571,1579|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1571,1579|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1571,1579|true|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|1589,1595|true|false|false|||change
Finding|Functional Concept|History of Present Illness|1589,1595|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1589,1595|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|History of Present Illness|1589,1598|true|false|false|C0392747|Changing|change in
Attribute|Clinical Attribute|History of Present Illness|1599,1604|true|false|false|C1717255||edema
Event|Event|History of Present Illness|1599,1604|true|false|false|||edema
Finding|Pathologic Function|History of Present Illness|1599,1604|true|false|false|C0013604|Edema|edema
Event|Event|History of Present Illness|1623,1628|false|false|false|||visit
Finding|Social Behavior|History of Present Illness|1623,1628|false|false|false|C0545082|Visit|visit
Event|Event|History of Present Illness|1634,1640|false|false|false|||denies
Event|Event|History of Present Illness|1652,1657|true|false|false|||fever
Finding|Finding|History of Present Illness|1652,1657|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1652,1657|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1659,1665|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1659,1665|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|1667,1673|true|false|false|||sweats
Finding|Body Substance|History of Present Illness|1667,1673|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|1667,1673|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Disorder|Disease or Syndrome|History of Present Illness|1675,1678|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|History of Present Illness|1675,1678|false|false|false|||PND
Finding|Gene or Genome|History of Present Illness|1675,1678|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|History of Present Illness|1681,1690|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|1681,1690|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1681,1690|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|History of Present Illness|1695,1705|false|false|false|||positional
Finding|Finding|History of Present Illness|1695,1705|false|false|false|C0240795|positional|positional
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1706,1715|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|History of Present Illness|1706,1715|false|false|false|C1179435|Protein Component|component
Event|Event|History of Present Illness|1706,1715|false|false|false|||component
Finding|Conceptual Entity|History of Present Illness|1706,1715|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|History of Present Illness|1706,1715|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|History of Present Illness|1706,1715|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Attribute|Clinical Attribute|History of Present Illness|1719,1723|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1719,1723|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1719,1723|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1719,1723|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|1737,1744|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1745,1750|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1745,1756|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1745,1756|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|1751,1756|false|false|false|||signs
Finding|Finding|History of Present Illness|1751,1756|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1751,1756|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Lab|Laboratory or Test Result|History of Present Illness|1791,1795|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1796,1803|false|false|false|||notable
Disorder|Disease or Syndrome|History of Present Illness|1808,1820|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|History of Present Illness|1808,1820|false|false|false|||leukocytosis
Finding|Finding|History of Present Illness|1808,1820|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Attribute|Clinical Attribute|History of Present Illness|1830,1840|false|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|History of Present Illness|1830,1840|false|false|false|||hematocrit
Finding|Finding|History of Present Illness|1830,1840|false|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|History of Present Illness|1830,1840|false|false|false|C0018935|Hematocrit Measurement|hematocrit
Drug|Organic Chemical|History of Present Illness|1853,1860|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|History of Present Illness|1853,1860|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|History of Present Illness|1853,1860|false|false|false|||lactate
Procedure|Laboratory Procedure|History of Present Illness|1853,1860|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|History of Present Illness|1869,1879|false|false|false|||Urinalysis
Procedure|Laboratory Procedure|History of Present Illness|1869,1879|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|Urinalysis
Disorder|Cell or Molecular Dysfunction|History of Present Illness|1884,1892|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|History of Present Illness|1884,1892|false|false|false|||positive
Finding|Classification|History of Present Illness|1884,1892|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|History of Present Illness|1884,1892|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Anatomy|Cell|History of Present Illness|1918,1923|false|false|false|C0007634|Cells|cells
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1925,1928|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|History of Present Illness|1925,1928|true|false|false|||CTA
Finding|Gene or Genome|History of Present Illness|1925,1928|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|1925,1928|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|History of Present Illness|1933,1941|false|false|false|||negative
Finding|Classification|History of Present Illness|1933,1941|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1933,1941|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1933,1941|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|History of Present Illness|1933,1945|false|false|false|C0205160|Negative|negative for
Drug|Pharmacologic Substance|History of Present Illness|1946,1953|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|History of Present Illness|1946,1953|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|History of Present Illness|1946,1953|true|false|false|||central
Procedure|Laboratory Procedure|History of Present Illness|1946,1953|true|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1954,1963|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|1954,1963|true|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|1954,1963|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|1954,1971|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolus
Event|Event|History of Present Illness|1964,1971|true|false|false|||embolus
Finding|Finding|History of Present Illness|1964,1971|true|false|false|C1704212;C2046122|Embolus|embolus
Event|Event|History of Present Illness|1973,1978|true|false|false|||focal
Disorder|Disease or Syndrome|History of Present Illness|1980,1993|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|History of Present Illness|1980,1993|false|false|false|||consolidation
Anatomy|Tissue|History of Present Illness|1998,2005|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|History of Present Illness|1998,2005|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|History of Present Illness|1998,2014|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|History of Present Illness|1998,2014|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|History of Present Illness|1998,2014|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|History of Present Illness|2006,2014|false|false|false|||effusion
Finding|Body Substance|History of Present Illness|2006,2014|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|History of Present Illness|2006,2014|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|History of Present Illness|2006,2014|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|History of Present Illness|2027,2033|false|false|false|||reveal
Finding|Intellectual Product|History of Present Illness|2027,2033|false|false|false|C5444168|Registry to Evaluate Early and Long-Term Pulmonary Arterial (PAH) Hypertension Disease Management (REVEAL)|reveal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2047,2056|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|2047,2056|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|2047,2056|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|History of Present Illness|2047,2064|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|History of Present Illness|2057,2064|false|false|false|||nodules
Finding|Finding|History of Present Illness|2069,2073|false|false|false|C5575035|Well (answer to question)|well
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2077,2085|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Finding|History of Present Illness|2077,2091|false|false|false|C0019209|Hepatomegaly|enlarged liver
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2086,2091|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|History of Present Illness|2086,2091|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|History of Present Illness|2086,2091|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|History of Present Illness|2086,2091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|History of Present Illness|2086,2091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|History of Present Illness|2086,2091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|History of Present Illness|2086,2091|false|false|false|||liver
Finding|Finding|History of Present Illness|2086,2091|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|History of Present Illness|2086,2091|false|false|false|C0872387|Procedures on liver|liver
Event|Event|History of Present Illness|2098,2104|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|2098,2104|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Neoplastic Process|History of Present Illness|2105,2115|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|History of Present Illness|2105,2115|false|false|false|||metastases
Finding|Finding|History of Present Illness|2105,2115|false|false|false|C1513183|Metastatic Lesion|metastases
Event|Event|History of Present Illness|2117,2120|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|2117,2120|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|2117,2120|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|History of Present Illness|2125,2136|false|false|false|||interpreted
Anatomy|Body Space or Junction|History of Present Illness|2140,2145|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|2140,2145|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|2140,2145|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|2140,2145|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Disorder|Disease or Syndrome|History of Present Illness|2140,2157|false|false|false|C0039239|Sinus Tachycardia|sinus tachycardia
Finding|Finding|History of Present Illness|2140,2157|false|false|false|C2108109;C5235163|Sinus Tachycardia by ECG Finding;continuous electrocardiogram sinus tachycardia|sinus tachycardia
Event|Event|History of Present Illness|2146,2157|false|false|false|||tachycardia
Finding|Finding|History of Present Illness|2146,2157|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Intellectual Product|History of Present Illness|2167,2174|false|false|false|C0282416|Overall Publication Type|overall
Event|Event|History of Present Illness|2175,2185|false|false|false|||consistent
Finding|Idea or Concept|History of Present Illness|2175,2185|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|History of Present Illness|2175,2190|false|false|false|C0332290|Consistent with|consistent with
Drug|Antibiotic|History of Present Illness|2198,2209|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Drug|Organic Chemical|History of Present Illness|2198,2209|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Event|Event|History of Present Illness|2198,2209|false|false|false|||Ceftriaxone
Drug|Antibiotic|History of Present Illness|2210,2222|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|2210,2222|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|2210,2222|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|2210,2222|false|false|false|||azithromycin
Event|Event|History of Present Illness|2229,2238|false|false|false|||initiated
Finding|Finding|History of Present Illness|2243,2251|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|History of Present Illness|2252,2261|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|History of Present Illness|2252,2261|false|false|false|||pneumonia
Drug|Food|History of Present Illness|2263,2268|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|History of Present Illness|2263,2274|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|History of Present Illness|2263,2274|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|History of Present Illness|2269,2274|false|false|false|||signs
Finding|Finding|History of Present Illness|2269,2274|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|2269,2274|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|History of Present Illness|2279,2287|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|2279,2287|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2279,2287|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2279,2287|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|2337,2344|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|2337,2344|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|2337,2344|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2352,2357|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|2364,2371|false|false|false|||reports
Event|Event|History of Present Illness|2377,2386|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|2377,2396|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|2377,2396|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|2390,2396|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|2401,2409|false|false|false|||improved
Anatomy|Body Location or Region|History of Present Illness|2427,2432|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2427,2432|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2427,2437|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2427,2437|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2433,2437|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2433,2437|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2433,2437|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2433,2437|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|2433,2442|false|false|false|C0908489|Pain-Free|pain free
Event|Event|History of Present Illness|2438,2442|false|false|false|||free
Finding|Functional Concept|History of Present Illness|2438,2442|false|false|false|C0332296|Free of (attribute)|free
Event|Event|Past Medical History|2472,2475|false|false|false|||OMR
Finding|Gene or Genome|Past Medical History|2472,2475|false|false|false|C1412647|ATP5F1A gene|OMR
Finding|Functional Concept|Past Medical History|2479,2489|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Past Medical History|2479,2496|false|false|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|Past Medical History|2490,2496|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|2490,2496|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2500,2507|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Past Medical History|2500,2507|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Past Medical History|2500,2507|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Past Medical History|2500,2507|false|false|false|||unknown
Finding|Finding|Past Medical History|2500,2507|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Past Medical History|2500,2507|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Past Medical History|2500,2507|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Past Medical History|2500,2507|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Finding|Past Medical History|2518,2522|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Past Medical History|2518,2522|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Past Medical History|2518,2522|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Past Medical History|2518,2528|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|Past Medical History|2518,2528|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|Past Medical History|2523,2528|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Past Medical History|2523,2528|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Event|Event|Past Medical History|2529,2532|false|false|false|||SBO
Procedure|Diagnostic Procedure|Past Medical History|2541,2563|false|false|false|C0085704|Exploratory laparotomy|exploratory laparotomy
Event|Event|Past Medical History|2553,2563|false|false|false|||laparotomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2553,2563|false|false|false|C0023038|Laparotomy|laparotomy
Event|Event|Past Medical History|2565,2570|false|false|false|||lysis
Finding|Cell Function|Past Medical History|2565,2570|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Finding|Pathologic Function|Past Medical History|2565,2570|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Event|Event|Past Medical History|2575,2584|false|false|false|||adhesions
Finding|Pathologic Function|Past Medical History|2575,2584|false|false|false|C0001511|Tissue Adhesions|adhesions
Anatomy|Body Location or Region|Past Medical History|2590,2601|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2590,2601|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2590,2611|false|false|false|C0192601|Small intestine excision|small bowel resection
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2596,2601|false|false|false|C0021853|Intestines|bowel
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2596,2611|false|false|false|C0741614|Bowel resection|bowel resection
Event|Event|Past Medical History|2602,2611|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2602,2611|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|Past Medical History|2617,2634|false|false|false|||enteroenterostomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2617,2634|false|false|false|C0192711;C0192741|Anastomosis of intestine;Anastomosis of small intestine to small intestine|enteroenterostomy
Disorder|Neoplastic Process|Past Medical History|2638,2647|false|false|false|C0007095|Carcinoid Tumor|carcinoid
Event|Event|Past Medical History|2638,2647|false|false|false|||carcinoid
Disorder|Disease or Syndrome|Past Medical History|2650,2664|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Past Medical History|2650,2664|false|false|false|||hyperlipidemia
Finding|Finding|Past Medical History|2650,2664|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Drug|Organic Chemical|Past Medical History|2667,2674|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Past Medical History|2667,2674|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Past Medical History|2667,2674|false|false|false|C0042890|Vitamins|vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Past Medical History|2667,2678|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Organic Chemical|Past Medical History|2667,2678|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Pharmacologic Substance|Past Medical History|2667,2678|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Vitamin|Past Medical History|2667,2678|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Procedure|Laboratory Procedure|Past Medical History|2667,2678|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|vitamin B12
Disorder|Disease or Syndrome|Past Medical History|2667,2689|false|false|false|C0042847|Vitamin B 12 Deficiency|vitamin B12 deficiency
Finding|Finding|Past Medical History|2667,2689|false|false|false|C5886863|Decreased circulating vitamin B12 concentration|vitamin B12 deficiency
Event|Event|Past Medical History|2675,2678|false|false|false|||B12
Finding|Gene or Genome|Past Medical History|2675,2678|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Disorder|Disease or Syndrome|Past Medical History|2679,2689|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Past Medical History|2679,2689|false|false|false|||deficiency
Finding|Functional Concept|Past Medical History|2679,2689|false|false|false|C0011155|Deficiency|deficiency
Anatomy|Body Location or Region|Past Medical History|2692,2700|false|false|false|C0027530|Neck|cervical
Disorder|Disease or Syndrome|Past Medical History|2701,2704|false|false|false|C0029408|Degenerative polyarthritis|DJD
Event|Event|Past Medical History|2701,2704|false|false|false|||DJD
Disorder|Disease or Syndrome|Past Medical History|2707,2721|false|false|false|C0029408|Degenerative polyarthritis|osteoarthritis
Event|Event|Past Medical History|2707,2721|false|false|false|||osteoarthritis
Anatomy|Body Location or Region|Past Medical History|2730,2734|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2730,2734|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Past Medical History|2730,2734|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Past Medical History|2730,2734|false|false|false|C0740941|Lung Problem|lung
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2730,2744|false|false|false|C0396565|Lung excision|lung resection
Event|Event|Past Medical History|2735,2744|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2735,2744|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|Past Medical History|2763,2775|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|2763,2775|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2763,2775|false|false|false|C0020699|Hysterectomy|hysterectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2787,2792|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2789,2792|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Past Medical History|2789,2792|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Past Medical History|2789,2792|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Past Medical History|2789,2792|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Past Medical History|2789,2792|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2789,2792|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|Past Medical History|2793,2800|false|false|false|||surgery
Finding|Finding|Past Medical History|2793,2800|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Past Medical History|2793,2800|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Past Medical History|2793,2800|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2793,2800|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Family Medical History|2844,2847|false|false|false|||OMR
Finding|Gene or Genome|Family Medical History|2844,2847|false|false|false|C1412647|ATP5F1A gene|OMR
Event|Event|Family Medical History|2849,2855|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|2849,2855|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|Family Medical History|2858,2862|false|false|false|||Died
Finding|Finding|Family Medical History|2858,2862|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|Died
Finding|Organism Function|Family Medical History|2858,2862|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|Died
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2866,2876|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2866,2876|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|Family Medical History|2866,2876|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|Family Medical History|2866,2876|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Disorder|Neoplastic Process|Family Medical History|2866,2883|false|false|false|C0235974;C0346647|Malignant neoplasm of pancreas;Pancreatic carcinoma|pancreatic cancer
Disorder|Neoplastic Process|Family Medical History|2877,2883|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|2877,2883|false|false|false|||cancer
Attribute|Clinical Attribute|Family Medical History|2887,2890|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|2887,2890|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|2887,2890|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|2887,2890|false|false|false|||age
Finding|Conceptual Entity|Family Medical History|2898,2904|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2898,2904|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|2907,2911|false|false|false|||Died
Finding|Finding|Family Medical History|2907,2911|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|Died
Finding|Organism Function|Family Medical History|2907,2911|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|Died
Disorder|Disease or Syndrome|Family Medical History|2919,2926|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|2919,2926|false|false|false|||disease
Attribute|Clinical Attribute|Family Medical History|2930,2933|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|2930,2933|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|2930,2933|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|General Exam|2960,2969|false|false|false|||admission
Procedure|Health Care Activity|General Exam|2960,2969|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Space or Junction|General Exam|2991,2996|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|2991,2996|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|2991,2996|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|2991,2996|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|General Exam|3008,3015|false|false|false|||GENERAL
Finding|Classification|General Exam|3008,3015|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3008,3015|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|3027,3036|false|false|false|||appearing
Event|Event|General Exam|3038,3046|false|false|false|||speaking
Event|Event|General Exam|3055,3064|false|false|false|||sentences
Finding|Intellectual Product|General Exam|3055,3064|false|false|false|C0876929|Sentence|sentences
Anatomy|Body Location or Region|General Exam|3067,3072|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3081,3087|false|false|false|||PERRLA
Finding|Finding|General Exam|3081,3087|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|General Exam|3089,3093|false|false|false|||EOMI
Event|Event|General Exam|3103,3112|false|false|false|||anicteric
Finding|Finding|General Exam|3103,3112|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3114,3117|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3114,3117|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3120,3124|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3120,3124|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3120,3124|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|3126,3132|true|false|false|||supple
Finding|Functional Concept|General Exam|3126,3132|true|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3137,3140|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3137,3140|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3137,3140|true|false|false|||LAD
Finding|Gene or Genome|General Exam|3137,3140|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|3145,3148|true|false|false|||JVD
Finding|Finding|General Exam|3145,3148|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|General Exam|3151,3156|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|General Exam|3151,3156|true|false|false|C0741025|Chest problem|CHEST
Finding|Intellectual Product|General Exam|3158,3162|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|General Exam|3176,3180|false|false|false|C2598155||pain
Event|Event|General Exam|3176,3180|false|false|false|||pain
Finding|Functional Concept|General Exam|3176,3180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|3176,3180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|3184,3188|false|false|false|||palp
Finding|Conceptual Entity|General Exam|3184,3188|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Finding|Gene or Genome|General Exam|3184,3188|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Event|Event|General Exam|3217,3221|true|false|false|||mass
Finding|Finding|General Exam|3217,3221|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|3217,3221|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3217,3221|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|General Exam|3224,3229|true|false|false|C0024109|Lung|LUNGS
Finding|Intellectual Product|General Exam|3231,3235|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|General Exam|3236,3244|false|false|false|||aeration
Procedure|Therapeutic or Preventive Procedure|General Exam|3236,3244|false|false|false|C2215609|aeration|aeration
Drug|Amino Acid, Peptide, or Protein|General Exam|3260,3263|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|3260,3263|true|false|false|||CTA
Finding|Gene or Genome|General Exam|3260,3263|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|3260,3263|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Attribute|Clinical Attribute|General Exam|3283,3287|true|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|General Exam|3283,3287|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|General Exam|3283,3287|true|false|false|||resp
Event|Event|General Exam|3289,3298|true|false|false|||unlabored
Finding|Functional Concept|General Exam|3289,3298|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|General Exam|3303,3319|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|3303,3323|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|3313,3319|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|3313,3319|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|3320,3323|true|false|false|||use
Finding|Functional Concept|General Exam|3320,3323|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|3320,3323|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|General Exam|3326,3331|true|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|General Exam|3326,3331|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|General Exam|3326,3331|true|false|false|||HEART
Finding|Sign or Symptom|General Exam|3326,3331|true|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|General Exam|3333,3338|false|false|false|||clear
Finding|Idea or Concept|General Exam|3333,3338|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|General Exam|3351,3356|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|3351,3356|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|3351,3356|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|General Exam|3351,3363|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|General Exam|3351,3363|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|General Exam|3351,3363|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Event|Event|General Exam|3357,3363|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3357,3363|false|false|false|C0037709||sounds
Event|Event|General Exam|3365,3377|false|false|false|||tachycardiac
Event|Event|General Exam|3382,3389|false|false|false|||regular
Event|Event|General Exam|3391,3397|false|false|false|||rhythm
Finding|Finding|General Exam|3391,3397|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3391,3397|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|3404,3407|false|false|false|||SEM
Finding|Finding|General Exam|3404,3407|false|false|false|C0694547|SYSTOLIC EJECTION MURMUR|SEM
Anatomy|Body Location or Region|General Exam|3420,3427|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3420,3427|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3420,3427|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3420,3427|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|3436,3441|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3436,3448|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3442,3448|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3442,3448|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|General Exam|3450,3454|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3450,3454|false|false|false|||soft
Finding|Intellectual Product|General Exam|3456,3460|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|General Exam|3461,3471|false|false|false|||tenderness
Finding|Mental Process|General Exam|3461,3471|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3461,3471|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|General Exam|3475,3479|false|false|false|||palp
Finding|Conceptual Entity|General Exam|3475,3479|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Finding|Gene or Genome|General Exam|3475,3479|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Event|Event|General Exam|3501,3511|true|false|false|||pronounced
Anatomy|Body Location or Region|General Exam|3519,3522|true|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|General Exam|3543,3550|true|false|false|||rebound
Event|Event|General Exam|3554,3562|true|false|false|||guarding
Finding|Finding|General Exam|3554,3562|true|false|false|C0427198|Protective muscle spasm|guarding
Finding|Finding|General Exam|3564,3578|true|false|false|C0577045|Liver palpable|palpable liver
Anatomy|Body Part, Organ, or Organ Component|General Exam|3573,3578|true|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|3573,3578|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|3573,3578|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|3573,3578|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|3573,3578|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|3573,3578|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|3573,3578|true|false|false|||liver
Finding|Finding|General Exam|3573,3578|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|3573,3578|true|false|false|C0872387|Procedures on liver|liver
Finding|Finding|General Exam|3573,3583|true|false|false|C0426689|Liver edge|liver edge
Event|Event|General Exam|3579,3583|false|false|false|||edge
Finding|Conceptual Entity|General Exam|3579,3583|false|false|false|C2697523|Graph Edge|edge
Anatomy|Body Part, Organ, or Organ Component|General Exam|3586,3597|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|3599,3603|false|false|false|||left
Finding|Functional Concept|General Exam|3599,3603|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|General Exam|3606,3611|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|General Exam|3612,3628|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|3615,3622|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|3615,3628|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|3623,3628|false|false|false|C1717255||edema
Event|Event|General Exam|3623,3628|false|false|false|||edema
Finding|Pathologic Function|General Exam|3623,3628|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|3636,3640|false|false|false|C0230444|Shin|shin
Drug|Food|General Exam|3646,3652|false|false|false|C5890763||pulses
Event|Event|General Exam|3646,3652|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3646,3652|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3646,3652|false|false|false|C0034107|Pulse taking|pulses
Finding|Organ or Tissue Function|General Exam|3646,3659|false|false|false|C0232142||pulses radial
Event|Event|General Exam|3653,3659|false|false|false|||radial
Finding|Conceptual Entity|General Exam|3653,3659|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Event|Event|General Exam|3676,3681|false|false|false|||awake
Finding|Finding|General Exam|3676,3681|false|false|false|C0234422|Awake (finding)|awake
Event|Event|General Exam|3683,3684|false|false|false|||A
Anatomy|Body System|General Exam|3690,3693|false|false|false|C3714787|Central Nervous System|CNs
Finding|Finding|General Exam|3709,3715|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|3717,3723|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|3717,3723|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Attribute|Clinical Attribute|General Exam|3717,3732|false|false|false|C4050373||muscle strength
Finding|Organ or Tissue Function|General Exam|3717,3732|false|false|false|C0517349|Muscle Strength|muscle strength
Event|Event|General Exam|3724,3732|false|false|false|||strength
Finding|Idea or Concept|General Exam|3724,3732|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|3750,3759|false|false|false|||sensation
Finding|Finding|General Exam|3750,3759|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3750,3759|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3750,3759|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|3768,3774|false|false|false|||intact
Finding|Finding|General Exam|3768,3774|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3779,3788|false|false|false|||discharge
Finding|Body Substance|General Exam|3779,3788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|3779,3788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|3779,3788|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|3779,3788|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|General Exam|3828,3835|false|false|false|||GENERAL
Finding|Classification|General Exam|3828,3835|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3828,3835|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|3837,3842|false|false|false|C0028754|Obesity|obese
Event|Event|General Exam|3837,3842|false|false|false|||obese
Disorder|Disease or Syndrome|General Exam|3844,3847|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3844,3847|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3844,3847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3844,3847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3844,3847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|3844,3847|false|false|false|||NAD
Finding|Finding|General Exam|3844,3847|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|3849,3854|false|false|false|||lying
Disorder|Disease or Syndrome|General Exam|3858,3861|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|3858,3861|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|General Exam|3875,3886|false|false|false|C0233471|Flat affect|flat affect
Event|Event|General Exam|3880,3886|false|false|false|||affect
Finding|Mental Process|General Exam|3880,3886|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|3880,3886|false|false|false|C2237113|assessment of affect|affect
Finding|Intellectual Product|General Exam|3892,3896|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Finding|General Exam|3892,3908|false|false|false|C1445953|Poor eye contact|poor eye contact
Anatomy|Body Location or Region|General Exam|3897,3900|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|General Exam|3897,3900|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|General Exam|3897,3900|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|General Exam|3897,3900|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|General Exam|3897,3900|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|General Exam|3897,3900|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|General Exam|3897,3900|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Social Behavior|General Exam|3897,3908|false|false|false|C0870532|eye contact|eye contact
Event|Activity|General Exam|3901,3908|false|false|false|C3812666|Personal Contact|contact
Event|Event|General Exam|3901,3908|false|false|false|||contact
Finding|Functional Concept|General Exam|3901,3908|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|General Exam|3901,3908|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|General Exam|3901,3908|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|General Exam|3901,3908|false|false|false|C0392367|Physical contact|contact
Anatomy|Body Location or Region|General Exam|3909,3914|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3916,3920|false|false|false|||NCAT
Event|Event|General Exam|3922,3926|false|false|false|||EOMI
Finding|Intellectual Product|General Exam|3928,3932|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|3933,3940|false|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|3933,3948|false|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|General Exam|3941,3948|false|false|false|C0022346|Icterus|icterus
Anatomy|Body Part, Organ, or Organ Component|General Exam|3955,3966|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|General Exam|3955,3966|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|General Exam|3955,3966|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|General Exam|3955,3966|false|false|false|||conjunctiva
Finding|Body Substance|General Exam|3955,3966|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|General Exam|3955,3966|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|General Exam|3955,3966|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|General Exam|3968,3971|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3968,3971|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Intellectual Product|General Exam|3974,3978|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Sign or Symptom|General Exam|3974,3988|false|false|false|C0149758|Poor dentition|poor dentition
Anatomy|Body Part, Organ, or Organ Component|General Exam|3979,3988|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Finding|Intellectual Product|General Exam|3990,3994|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|4004,4015|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|General Exam|4004,4015|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|General Exam|4004,4015|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|General Exam|4004,4015|false|false|false|||conjunctiva
Finding|Body Substance|General Exam|4004,4015|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|General Exam|4004,4015|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|General Exam|4004,4015|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Location or Region|General Exam|4017,4021|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|4017,4021|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|4017,4021|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|4023,4029|true|false|false|||supple
Finding|Functional Concept|General Exam|4023,4029|true|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|4034,4037|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|4034,4037|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|4034,4037|true|false|false|||LAD
Finding|Gene or Genome|General Exam|4034,4037|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|4040,4047|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4040,4047|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|4049,4060|false|false|false|||tachycardic
Event|Event|General Exam|4065,4072|true|false|false|||regular
Anatomy|Body Location or Region|General Exam|4090,4094|true|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|General Exam|4090,4094|true|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|General Exam|4090,4094|true|false|false|C0024115|Lung diseases|LUNG
Event|Event|General Exam|4090,4094|true|false|false|||LUNG
Finding|Finding|General Exam|4090,4094|true|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|General Exam|4096,4100|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|4096,4100|false|false|false|||CTAB
Disorder|Disease or Syndrome|General Exam|4104,4112|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Finding|General Exam|4121,4144|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|General Exam|4131,4137|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|General Exam|4131,4144|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|General Exam|4138,4144|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4138,4144|false|false|false|C0037709||sounds
Finding|Functional Concept|General Exam|4148,4153|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|4155,4159|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|4155,4159|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|4155,4159|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4155,4159|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|4155,4159|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|4155,4159|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Event|Event|General Exam|4161,4165|false|false|false|||exam
Finding|Functional Concept|General Exam|4161,4165|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4161,4165|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|4166,4173|false|false|false|||limited
Disorder|Neoplastic Process|General Exam|4174,4183|true|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|General Exam|4174,4183|true|false|false|||secondary
Finding|Functional Concept|General Exam|4174,4183|true|false|false|C1522484|metastatic qualifier|secondary
Anatomy|Anatomical Structure|General Exam|4187,4191|true|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|4187,4191|true|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|4187,4191|true|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|General Exam|4187,4199|true|false|false|C1318474|Assessment of body build|body habitus
Event|Event|General Exam|4192,4199|true|false|false|||habitus
Attribute|Clinical Attribute|General Exam|4204,4212|true|false|false|C0080078|Range of Motion, Articular|mobility
Event|Event|General Exam|4204,4212|true|false|false|||mobility
Finding|Finding|General Exam|4204,4212|true|false|false|C0425245|Mobility finding|mobility
Event|Event|General Exam|4222,4223|true|false|false|||r
Disorder|Congenital Abnormality|General Exam|4228,4244|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|4228,4248|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|4238,4244|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|4238,4244|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|4245,4248|true|false|false|||use
Finding|Functional Concept|General Exam|4245,4248|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|4245,4248|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Location or Region|General Exam|4249,4256|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4249,4256|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4249,4256|true|false|false|||ABDOMEN
Finding|Finding|General Exam|4249,4256|true|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4258,4263|true|false|false|C0028754|Obesity|obese
Event|Event|General Exam|4258,4263|true|false|false|||obese
Event|Event|General Exam|4285,4293|true|false|false|||guarding
Finding|Finding|General Exam|4285,4293|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Governmental or Regulatory Activity|General Exam|4305,4309|true|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|General Exam|4314,4322|false|false|false|||firmness
Anatomy|Body Location or Region|General Exam|4336,4343|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|4336,4343|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|4336,4343|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|General Exam|4336,4347|false|false|false|C0000726|Abdomen|abdomen and
Event|Event|General Exam|4348,4354|false|false|false|||tender
Event|Event|General Exam|4358,4367|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|4358,4367|false|false|false|C0030247|Palpation|palpation
Event|Governmental or Regulatory Activity|General Exam|4379,4383|false|false|false|C1510751|Academic Research Enhancement Awards|area
Anatomy|Body Part, Organ, or Organ Component|General Exam|4385,4396|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Drug|Food|General Exam|4409,4415|false|false|false|C5890763||pulses
Event|Event|General Exam|4409,4415|false|false|false|||pulses
Finding|Physiologic Function|General Exam|4409,4415|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4409,4415|false|false|false|C0034107|Pulse taking|pulses
Finding|Finding|General Exam|4429,4445|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|4432,4439|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4432,4445|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4440,4445|false|false|false|C1717255||edema
Event|Event|General Exam|4440,4445|false|false|false|||edema
Finding|Pathologic Function|General Exam|4440,4445|false|false|false|C0013604|Edema|edema
Event|Event|General Exam|4478,4487|true|false|false|||asterixis
Finding|Sign or Symptom|General Exam|4478,4487|true|false|false|C0232766|Asterixis|asterixis
Event|Event|General Exam|4489,4495|true|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|4505,4516|true|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|4527,4535|false|false|false|||movement
Finding|Organism Function|General Exam|4527,4535|false|false|false|C0026649|Movement|movement
Phenomenon|Natural Phenomenon or Process|General Exam|4543,4550|false|false|false|C0282189|Gravity (physical force)|gravity
Attribute|Clinical Attribute|General Exam|4555,4561|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|General Exam|4562,4569|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|General Exam|4562,4569|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Finding|Idea or Concept|General Exam|4576,4580|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|General Exam|4581,4585|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|General Exam|4581,4585|false|false|false|C0741992|Hand problem|hand
Disorder|Disease or Syndrome|General Exam|4587,4591|false|false|false|C0021400|Influenza|grip
Event|Event|General Exam|4587,4591|false|false|false|||grip
Finding|Organism Function|General Exam|4587,4591|false|false|false|C0220843|grasp|grip
Attribute|Clinical Attribute|General Exam|4587,4600|false|false|false|C2598165||grip strength
Event|Event|General Exam|4592,4600|false|false|false|||strength
Finding|Idea or Concept|General Exam|4592,4600|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|4631,4640|false|false|false|||admission
Procedure|Health Care Activity|General Exam|4631,4640|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|General Exam|4654,4659|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4654,4659|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4654,4659|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4660,4663|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4670,4673|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4670,4673|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4670,4673|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4680,4683|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4680,4683|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4680,4683|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4680,4683|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4689,4692|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4689,4692|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4700,4703|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4700,4703|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4700,4703|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4700,4703|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4700,4703|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4707,4710|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4707,4710|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4707,4710|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4707,4710|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4707,4710|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4707,4710|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4717,4721|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4738,4741|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4758,4763|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4758,4763|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4758,4763|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|4776,4782|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4789,4794|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4789,4794|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4789,4794|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4800,4803|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|4800,4803|false|false|false|||Eos
Finding|Gene or Genome|General Exam|4800,4803|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4829,4834|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4829,4834|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4829,4834|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4839,4842|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4839,4842|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4839,4842|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4864,4869|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4864,4869|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4864,4869|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4864,4877|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4864,4877|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4864,4877|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4870,4877|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4870,4877|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4870,4877|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4870,4877|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4870,4877|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4870,4877|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|4951,4956|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4951,4956|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4951,4956|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4957,4960|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4957,4960|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4957,4960|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4957,4960|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4957,4960|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4957,4960|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4957,4960|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4957,4960|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4964,4967|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4964,4967|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4964,4967|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4964,4967|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4964,4967|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|4964,4967|false|false|false|||AST
Finding|Gene or Genome|General Exam|4964,4967|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4988,4991|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|4988,4991|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|4988,4991|false|false|false|||CPK
Finding|Gene or Genome|General Exam|4988,4991|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|4988,4991|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|4999,5006|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4999,5006|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|5062,5067|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5062,5067|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5062,5067|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5068,5073|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|5068,5073|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|5068,5073|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|5068,5073|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|General Exam|5071,5073|false|false|false|||MB
Finding|Gene or Genome|General Exam|5071,5075|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|MB-1
Disorder|Disease or Syndrome|General Exam|5102,5107|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5102,5107|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5102,5107|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5102,5115|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|5108,5115|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|5108,5115|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|5108,5115|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|5108,5115|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|5108,5115|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|5108,5115|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|5108,5115|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|General Exam|5140,5145|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5140,5145|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5140,5145|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|5169,5174|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5169,5174|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5169,5174|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5169,5182|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|5175,5182|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|5175,5182|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|5175,5182|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|General Exam|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|5201,5212|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|5207,5212|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5207,5212|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Finding|Body Substance|General Exam|5253,5258|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5253,5258|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5253,5258|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|5253,5264|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|5259,5264|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|5259,5264|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|5265,5268|false|false|false|||NEG
Finding|Finding|General Exam|5265,5268|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|5269,5276|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|5269,5276|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|5269,5276|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|General Exam|5277,5280|false|false|false|||NEG
Finding|Finding|General Exam|5277,5280|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|5281,5288|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|5281,5288|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|5281,5288|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|5281,5288|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|5281,5288|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|General Exam|5293,5300|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5293,5300|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5293,5300|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5293,5300|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5293,5300|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5293,5300|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|5301,5304|false|false|false|||NEG
Finding|Finding|General Exam|5301,5304|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|5305,5311|false|false|false|C0022634|Ketones|Ketone
Disorder|Disease or Syndrome|General Exam|5351,5354|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|General Exam|5351,5354|false|false|false|||MOD
Finding|Body Substance|General Exam|5367,5372|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5367,5372|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5367,5372|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|5367,5376|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|General Exam|5373,5376|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5373,5376|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5373,5376|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|5379,5382|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|General Exam|5399,5404|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|General Exam|5399,5404|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5399,5404|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|General Exam|5399,5404|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|General Exam|5405,5409|false|false|false|||NONE
Disorder|Disease or Syndrome|General Exam|5411,5414|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|General Exam|5411,5414|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|General Exam|5411,5414|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|General Exam|5411,5414|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|General Exam|5411,5414|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|General Exam|5411,5414|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|General Exam|5411,5414|true|false|false|||Epi
Finding|Gene or Genome|General Exam|5411,5414|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|General Exam|5411,5414|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|General Exam|5411,5414|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|General Exam|5430,5435|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5430,5435|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5430,5435|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|5450,5459|false|false|false|||discharge
Finding|Body Substance|General Exam|5450,5459|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|5450,5459|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|5450,5459|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|5450,5459|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|General Exam|5473,5478|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5473,5478|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5473,5478|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|5479,5482|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|5489,5492|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5489,5492|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5489,5492|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5499,5502|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|5499,5502|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|5499,5502|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|5499,5502|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|5508,5511|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|5508,5511|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|5519,5522|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|5519,5522|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|5519,5522|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5519,5522|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5519,5522|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5526,5529|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5526,5529|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|5526,5529|false|false|false|||MCH
Finding|Gene or Genome|General Exam|5526,5529|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5526,5529|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5526,5529|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|5535,5539|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|5535,5539|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|5556,5559|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|5576,5581|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5576,5581|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5576,5581|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|5576,5589|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|5576,5589|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|5576,5589|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5582,5589|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5582,5589|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5582,5589|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5582,5589|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5582,5589|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5582,5589|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|5664,5669|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5664,5669|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5664,5669|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5664,5677|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|5670,5677|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5670,5677|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5670,5677|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5670,5677|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5670,5677|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|5670,5677|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|5670,5677|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5670,5677|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|General Exam|5701,5713|false|false|false|||Microbiology
Finding|Functional Concept|General Exam|5701,5713|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Finding|Intellectual Product|General Exam|5701,5713|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Procedure|Laboratory Procedure|General Exam|5701,5713|false|false|false|C0085672|Microbiology procedure|Microbiology
Disorder|Disease or Syndrome|General Exam|5715,5720|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|5715,5720|false|false|false|||Blood
Finding|Body Substance|General Exam|5715,5720|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|5734,5740|true|false|false|||growth
Finding|Finding|General Exam|5734,5740|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|General Exam|5734,5740|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|General Exam|5734,5740|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|General Exam|5734,5740|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|General Exam|5734,5740|true|false|false|C2911660|Growth action|growth
Finding|Body Substance|General Exam|5741,5746|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|General Exam|5741,5746|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|General Exam|5741,5746|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|General Exam|5757,5763|true|false|false|||growth
Finding|Finding|General Exam|5757,5763|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|General Exam|5757,5763|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|General Exam|5757,5763|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|General Exam|5757,5763|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|General Exam|5757,5763|true|false|false|C2911660|Growth action|growth
Disorder|Disease or Syndrome|General Exam|5764,5769|true|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|5764,5769|true|false|false|||Blood
Finding|Body Substance|General Exam|5764,5769|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|5783,5789|true|false|false|||growth
Finding|Finding|General Exam|5783,5789|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|General Exam|5783,5789|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|General Exam|5783,5789|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|General Exam|5783,5789|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|General Exam|5783,5789|true|false|false|C2911660|Growth action|growth
Event|Event|General Exam|5791,5800|true|false|false|||Pathology
Finding|Functional Concept|General Exam|5791,5800|true|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|Pathology
Finding|Pathologic Function|General Exam|5791,5800|true|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|Pathology
Procedure|Laboratory Procedure|General Exam|5791,5800|true|false|false|C0919386|Pathology procedure|Pathology
Anatomy|Body Part, Organ, or Organ Component|General Exam|5802,5807|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|General Exam|5802,5807|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|General Exam|5802,5807|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|General Exam|5802,5807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|General Exam|5802,5807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|General Exam|5802,5807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Event|Event|General Exam|5802,5807|false|false|false|||Liver
Finding|Finding|General Exam|5802,5807|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|General Exam|5802,5807|false|false|false|C0872387|Procedures on liver|Liver
Procedure|Diagnostic Procedure|General Exam|5802,5814|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|Liver biopsy
Procedure|Health Care Activity|General Exam|5802,5814|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|Liver biopsy
Event|Event|General Exam|5808,5814|false|false|false|||biopsy
Finding|Finding|General Exam|5808,5814|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|General Exam|5808,5814|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|General Exam|5808,5814|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|General Exam|5808,5814|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Anatomy|Body Part, Organ, or Organ Component|General Exam|5822,5827|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|General Exam|5822,5827|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|General Exam|5822,5827|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|General Exam|5822,5827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|General Exam|5822,5827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|General Exam|5822,5827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Event|Event|General Exam|5822,5827|false|false|false|||Liver
Finding|Finding|General Exam|5822,5827|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|General Exam|5822,5827|false|false|false|C0872387|Procedures on liver|Liver
Anatomy|Cell Component|General Exam|5829,5833|false|false|false|C1167518|viral nucleocapsid location|core
Finding|Body Substance|General Exam|5829,5833|false|false|false|C3274653|Core Specimen|core
Procedure|Diagnostic Procedure|General Exam|5829,5847|false|false|false|C1318309|Core needle biopsy|core needle biopsy
Finding|Intellectual Product|General Exam|5834,5840|false|false|false|C1546717||needle
Procedure|Diagnostic Procedure|General Exam|5834,5847|false|false|false|C0005560;C0936232;C1548887|Consent Type - Needle Biopsy;Needle biopsy (procedure);Puncture biopsy|needle biopsy
Procedure|Health Care Activity|General Exam|5834,5847|false|false|false|C0005560;C0936232;C1548887|Consent Type - Needle Biopsy;Needle biopsy (procedure);Puncture biopsy|needle biopsy
Event|Event|General Exam|5841,5847|false|false|false|||biopsy
Finding|Finding|General Exam|5841,5847|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|General Exam|5841,5847|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|General Exam|5841,5847|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|General Exam|5841,5847|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Neoplastic Process|General Exam|5853,5867|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|Adenocarcinoma
Event|Event|General Exam|5853,5867|false|false|false|||Adenocarcinoma
Event|Event|General Exam|5869,5878|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|General Exam|5883,5888|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|5883,5888|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|5883,5888|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|5883,5888|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|5883,5888|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|5883,5888|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|5883,5888|false|false|false|||liver
Finding|Finding|General Exam|5883,5888|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|5883,5888|false|false|false|C0872387|Procedures on liver|liver
Event|Event|General Exam|5890,5893|false|false|false|||see
Event|Event|General Exam|5901,5905|false|false|false|||Note
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5907,5933|false|false|false|C4317108|immunohistochemical stains|Immunohistochemical stains
Procedure|Laboratory Procedure|General Exam|5907,5933|false|false|false|C1508788|immunohistochemical stains procedure|Immunohistochemical stains
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5927,5933|false|false|false|C0038128|Stains|stains
Event|Event|General Exam|5927,5933|false|false|false|||stains
Finding|Molecular Function|General Exam|5927,5933|false|false|false|C2757062|Dyes [MoA]|stains
Procedure|Laboratory Procedure|General Exam|5927,5933|false|false|false|C0487602|Staining method|stains
Disorder|Neoplastic Process|General Exam|5954,5959|false|false|false|C0027651|Neoplasms|tumor
Finding|Finding|General Exam|5954,5959|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|General Exam|5954,5959|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Anatomy|Cell|General Exam|5954,5965|false|false|false|C0431085;C5551176|Tumor cells;Tumor cells, uncertain whether benign or malignant|tumor cells
Anatomy|Cell|General Exam|5960,5965|false|false|false|C0007634|Cells|cells
Disorder|Cell or Molecular Dysfunction|General Exam|5971,5979|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|General Exam|5971,5979|false|false|false|||positive
Finding|Classification|General Exam|5971,5979|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|5971,5979|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|5971,5983|false|false|false|C1446409|Positive|positive for
Event|Event|General Exam|5984,5988|false|false|false|||CK20
Finding|Gene or Genome|General Exam|5984,5988|false|false|false|C1426926;C3272788|KRT20 gene;KRT20 wt Allele|CK20
Drug|Antibiotic|General Exam|5993,5996|true|false|false|C0007538;C0285590|bicalutamide;cefadroxil|CDX
Drug|Organic Chemical|General Exam|5993,5996|true|false|false|C0007538;C0285590|bicalutamide;cefadroxil|CDX
Drug|Pharmacologic Substance|General Exam|5993,5996|true|false|false|C0007538;C0285590|bicalutamide;cefadroxil|CDX
Event|Event|General Exam|5993,5996|true|false|false|||CDX
Finding|Body Substance|General Exam|5993,5996|true|false|false|C4722223|Cell Line-Derived Xenograft|CDX
Procedure|Laboratory Procedure|General Exam|5993,5996|true|false|false|C5963431|Companion Diagnostic Test|CDX
Event|Event|General Exam|6004,6012|false|false|false|||negative
Finding|Classification|General Exam|6004,6012|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|6004,6012|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|6004,6012|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|General Exam|6004,6016|false|false|false|C0205160|Negative|negative for
Lab|Laboratory or Test Result|General Exam|6004,6030|false|false|false|C4698687|Negative for CK7 and TTF-1|negative for CK7 and TTF-1
Event|Event|General Exam|6017,6020|true|false|false|||CK7
Finding|Gene or Genome|General Exam|6017,6020|true|false|false|C1416745;C3272782|KRT7 gene;KRT7 wt Allele|CK7
Event|Event|General Exam|6025,6028|true|false|false|||TTF
Finding|Gene or Genome|General Exam|6025,6028|true|false|false|C1332112;C1705840|RHOH gene;RHOH wt Allele|TTF
Procedure|Therapeutic or Preventive Procedure|General Exam|6025,6028|true|false|false|C4087167|Tumour treating fields therapy|TTF
Drug|Amino Acid, Peptide, or Protein|General Exam|6025,6030|true|false|false|C0084785;C1452466;C1610981|NKX2-1 protein, human;TTF1 protein, human;thyroid transcription factor 1|TTF-1
Drug|Biologically Active Substance|General Exam|6025,6030|true|false|false|C0084785;C1452466;C1610981|NKX2-1 protein, human;TTF1 protein, human;thyroid transcription factor 1|TTF-1
Finding|Gene or Genome|General Exam|6025,6030|true|false|false|C1384616;C2347318;C3811254|NKX2-1 gene;NKX2-1 wt Allele;TTF1 wt Allele|TTF-1
Event|Event|General Exam|6040,6047|false|false|false|||results
Event|Event|General Exam|6052,6062|false|false|false|||consistent
Finding|Idea or Concept|General Exam|6052,6062|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|6052,6067|false|false|false|C0332290|Consistent with|consistent with
Disorder|Neoplastic Process|General Exam|6068,6078|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastasis
Event|Event|General Exam|6068,6078|false|false|false|||metastasis
Finding|Finding|General Exam|6068,6078|false|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Finding|Pathologic Function|General Exam|6068,6078|false|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Event|Event|General Exam|6108,6115|false|false|false|||Imaging
Finding|Finding|General Exam|6108,6115|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|6108,6115|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|General Exam|6117,6120|false|false|false|||EKG
Finding|Intellectual Product|General Exam|6117,6120|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|6117,6120|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|General Exam|6128,6133|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|General Exam|6128,6133|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|General Exam|6128,6133|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|General Exam|6128,6133|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Disorder|Disease or Syndrome|General Exam|6128,6145|false|false|false|C0039239|Sinus Tachycardia|Sinus tachycardia
Finding|Finding|General Exam|6128,6145|false|false|false|C2108109;C5235163|Sinus Tachycardia by ECG Finding;continuous electrocardiogram sinus tachycardia|Sinus tachycardia
Event|Event|General Exam|6134,6145|false|false|false|||tachycardia
Finding|Finding|General Exam|6134,6145|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Finding|General Exam|6147,6150|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|General Exam|6147,6150|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Event|Event|General Exam|6151,6158|false|false|false|||voltage
Disorder|Congenital Abnormality|General Exam|6197,6210|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|6197,6210|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|6197,6210|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|6237,6244|false|false|false|||tracing
Disorder|Congenital Abnormality|General Exam|6268,6281|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|6268,6281|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|6268,6281|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|6300,6309|false|false|false|||prominent
Procedure|Diagnostic Procedure|General Exam|6320,6332|false|false|false|C2318073|portable x-ray of chest|Portable CXR
Event|Event|General Exam|6329,6332|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|6329,6332|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Body Part, Organ, or Organ Component|General Exam|6352,6361|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|6352,6361|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|6352,6361|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Neoplastic Process|General Exam|6352,6372|false|false|false|C0153676|Secondary malignant neoplasm of lung|pulmonary metastases
Disorder|Neoplastic Process|General Exam|6362,6372|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|General Exam|6362,6372|false|false|false|||metastases
Finding|Finding|General Exam|6362,6372|false|false|false|C1513183|Metastatic Lesion|metastases
Finding|Finding|General Exam|6375,6383|false|false|false|C0332149|Possible|Possible
Finding|Intellectual Product|General Exam|6384,6388|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|6389,6398|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|6389,6398|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|6389,6398|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|6400,6408|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|General Exam|6409,6419|false|false|false|||congestion
Finding|Pathologic Function|General Exam|6409,6419|false|false|false|C0700148|Congestion|congestion
Finding|Finding|General Exam|6422,6425|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|General Exam|6422,6425|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Anatomy|Body Location or Region|General Exam|6426,6430|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|6426,6430|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|6426,6430|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|6426,6430|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|General Exam|6426,6438|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|General Exam|6431,6438|false|false|false|||volumes
Drug|Amino Acid, Peptide, or Protein|General Exam|6441,6444|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|6441,6444|false|false|false|||CTA
Finding|Gene or Genome|General Exam|6441,6444|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|6441,6444|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Drug|Pharmacologic Substance|General Exam|6459,6466|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|General Exam|6459,6466|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|General Exam|6459,6466|true|false|false|||central
Procedure|Laboratory Procedure|General Exam|6459,6466|true|false|false|C1879652|Central Minus|central
Finding|Functional Concept|General Exam|6480,6494|true|false|false|C0332555|Filling defect|filling defect
Disorder|Disease or Syndrome|General Exam|6488,6494|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|General Exam|6488,6494|true|false|false|||defect
Finding|Functional Concept|General Exam|6488,6494|true|false|false|C1457869|Defect|defect
Anatomy|Body Part, Organ, or Organ Component|General Exam|6502,6511|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|6502,6511|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|6502,6511|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|6513,6521|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|General Exam|6513,6521|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|General Exam|6513,6521|false|false|false|||arteries
Procedure|Health Care Activity|General Exam|6513,6521|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|General Exam|6523,6533|false|false|false|||Evaluation
Finding|Idea or Concept|General Exam|6523,6533|false|false|false|C1550157|Processing type - Evaluation|Evaluation
Procedure|Health Care Activity|General Exam|6523,6533|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|Evaluation
Finding|Finding|General Exam|6537,6553|false|false|false|C3829283|Limited a Little|slightly limited
Event|Event|General Exam|6546,6553|false|false|false|||limited
Finding|Functional Concept|General Exam|6546,6553|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|General Exam|6546,6553|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Functional Concept|General Exam|6572,6580|false|false|false|C1522229|Intravenous Bolus|IV bolus
Event|Event|General Exam|6575,6580|false|false|false|||bolus
Finding|Body Substance|General Exam|6575,6580|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|General Exam|6575,6580|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|General Exam|6575,6580|false|false|false|C1511237|bolus infusion|bolus
Anatomy|Body Part, Organ, or Organ Component|General Exam|6609,6618|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|6609,6618|true|false|false|C2707265||pulmonary
Finding|Finding|General Exam|6609,6618|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|General Exam|6609,6626|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|General Exam|6619,6626|false|false|false|||nodules
Event|Event|General Exam|6634,6638|false|false|false|||seen
Attribute|Clinical Attribute|General Exam|6653,6661|false|false|false|C5886017||CT study
Event|Event|General Exam|6656,6661|false|false|false|||study
Finding|Intellectual Product|General Exam|6656,6661|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|6656,6661|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|General Exam|6679,6688|false|false|false|||increased
Disorder|Disease or Syndrome|General Exam|6701,6714|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|6701,6714|true|false|false|||consolidation
Anatomy|Tissue|General Exam|6718,6725|true|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|6718,6725|true|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|General Exam|6718,6734|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|General Exam|6718,6734|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|General Exam|6718,6734|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|General Exam|6726,6734|true|false|false|||effusion
Finding|Body Substance|General Exam|6726,6734|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|6726,6734|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|6726,6734|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Procedure|Therapeutic or Preventive Procedure|General Exam|6742,6750|false|false|false|C1293134|Enlargement procedure|Enlarged
Finding|Finding|General Exam|6742,6756|false|false|false|C0019209|Hepatomegaly|Enlarged liver
Anatomy|Body Part, Organ, or Organ Component|General Exam|6751,6756|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|6751,6756|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|6751,6756|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|6751,6756|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|6751,6756|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|6751,6756|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|6751,6756|false|false|false|||liver
Finding|Finding|General Exam|6751,6756|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|6751,6756|false|false|false|C0872387|Procedures on liver|liver
Event|Event|General Exam|6781,6788|false|false|false|||lesions
Finding|Finding|General Exam|6781,6788|false|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|6796,6806|false|false|false|||suggestion
Finding|Idea or Concept|General Exam|6796,6806|false|false|false|C0038659;C1705535|suggestion;therapeutic suggestion|suggestion
Event|Event|General Exam|6810,6819|false|false|false|||increased
Event|Event|General Exam|6820,6826|false|false|false|||burden
Finding|Idea or Concept|General Exam|6820,6826|false|false|false|C2828008|Burden|burden
Disorder|Disease or Syndrome|General Exam|6830,6837|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|6830,6837|false|false|false|||disease
Finding|Functional Concept|General Exam|6840,6845|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|General Exam|6840,6860|false|false|false|C0230177|Structure of right upper quadrant of abdomen|Right upper quadrant
Event|Event|General Exam|6861,6871|false|false|false|||ultrasound
Finding|Functional Concept|General Exam|6861,6871|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|6861,6871|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|6861,6871|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Location or Region|General Exam|6897,6904|false|false|false|C0205054|Hepatic|hepatic
Finding|Functional Concept|General Exam|6905,6915|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|General Exam|6905,6923|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|General Exam|6905,6923|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|General Exam|6916,6923|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|6916,6923|false|false|false|||disease
Event|Event|General Exam|6929,6937|true|false|false|||evidence
Finding|Idea or Concept|General Exam|6929,6937|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|6929,6940|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|General Exam|6942,6949|true|false|false|C0521378|Biliary|biliary
Anatomy|Body Part, Organ, or Organ Component|General Exam|6942,6954|true|false|false|C0005400|Bile duct structure|biliary duct
Anatomy|Body Part, Organ, or Organ Component|General Exam|6950,6954|true|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Event|Event|General Exam|6955,6966|true|false|false|||obstruction
Finding|Finding|General Exam|6955,6966|true|false|false|C0028778|Obstruction|obstruction
Procedure|Diagnostic Procedure|General Exam|6969,6981|false|false|false|C2318073|portable x-ray of chest|Portable CXR
Event|Event|General Exam|6978,6981|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|6978,6981|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|General Exam|6992,6995|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|General Exam|6992,6995|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Anatomy|Body Location or Region|General Exam|6996,7000|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|6996,7000|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|6996,7000|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|6996,7000|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|General Exam|6996,7008|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|General Exam|7001,7008|false|false|false|||volumes
Finding|Intellectual Product|General Exam|7013,7017|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|7018,7027|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7018,7027|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7018,7027|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|General Exam|7018,7047|false|false|false|C5849517|Pulmonary vascular congestion|pulmonary vascular congestion
Anatomy|Body Part, Organ, or Organ Component|General Exam|7028,7036|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|General Exam|7037,7047|false|false|false|||congestion
Finding|Pathologic Function|General Exam|7037,7047|false|false|false|C0700148|Congestion|congestion
Event|Event|General Exam|7052,7061|false|false|false|||unchanged
Finding|Finding|General Exam|7052,7061|false|false|false|C0442739||unchanged
Finding|Finding|General Exam|7067,7070|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|General Exam|7067,7070|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Functional Concept|General Exam|7077,7082|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|General Exam|7092,7099|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|7092,7099|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|General Exam|7092,7108|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|General Exam|7092,7108|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|General Exam|7092,7108|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|General Exam|7100,7108|false|false|false|||effusion
Finding|Body Substance|General Exam|7100,7108|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|7100,7108|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|7100,7108|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Finding|General Exam|7116,7119|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|7116,7119|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|General Exam|7126,7135|true|false|false|||opacities
Finding|Finding|General Exam|7126,7135|true|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|General Exam|7126,7135|true|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Event|Event|General Exam|7139,7146|true|false|false|||suggest
Disorder|Disease or Syndrome|General Exam|7147,7156|true|true|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|7147,7156|true|false|false|||pneumonia
Anatomy|Body Location or Region|General Exam|7173,7177|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|7173,7177|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|General Exam|7173,7177|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|General Exam|7173,7177|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|General Exam|7173,7180|false|false|false|C0202691|CAT scan of head|head CT
Event|Event|General Exam|7178,7180|false|false|false|||CT
Finding|Intellectual Product|General Exam|7191,7196|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|General Exam|7197,7209|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|General Exam|7197,7209|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|7210,7217|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|7210,7217|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|General Exam|7210,7217|true|false|false|||process
Finding|Functional Concept|General Exam|7210,7217|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|7210,7217|true|false|false|C1522240|Process|process
Event|Event|General Exam|7223,7227|true|false|false|||mass
Finding|Finding|General Exam|7223,7227|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|7223,7227|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|7223,7227|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|General Exam|7231,7241|true|false|false|||identified
Event|Event|General Exam|7244,7247|false|false|false|||MRI
Finding|Gene or Genome|General Exam|7244,7247|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|General Exam|7244,7247|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|General Exam|7244,7247|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|General Exam|7257,7266|false|false|false|||sensitive
Finding|Functional Concept|General Exam|7257,7266|false|false|false|C0332324|Sensitive|sensitive
Event|Event|General Exam|7271,7281|false|false|false|||evaluation
Finding|Idea or Concept|General Exam|7271,7281|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|General Exam|7271,7281|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Disorder|Neoplastic Process|General Exam|7285,7295|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|General Exam|7285,7295|false|false|false|||metastases
Finding|Finding|General Exam|7285,7295|false|false|false|C1513183|Metastatic Lesion|metastases
Finding|Functional Concept|General Exam|7298,7302|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|General Exam|7298,7306|false|false|false|C0524471|Left hip region structure|Left hip
Anatomy|Body Part, Organ, or Organ Component|General Exam|7303,7306|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|7303,7306|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|7303,7306|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|7303,7306|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|7303,7306|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|7303,7306|false|false|false|C1292890|Procedure on hip|hip
Event|Event|General Exam|7307,7309|false|false|false|||XR
Finding|Pathologic Function|General Exam|7329,7334|true|false|false|C0024348|Lysis|lytic
Finding|Finding|General Exam|7329,7341|true|true|false|C0221204;C2021200|Lytic lesion|lytic lesion
Finding|Pathologic Function|General Exam|7329,7341|true|true|false|C0221204;C2021200|Lytic lesion|lytic lesion
Event|Event|General Exam|7335,7341|true|false|false|||lesion
Finding|Finding|General Exam|7335,7341|true|true|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|7335,7341|true|true|false|C0221198;C1546698|Lesion|lesion
Event|Event|General Exam|7355,7358|false|false|false|||MRI
Finding|Gene or Genome|General Exam|7355,7358|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|General Exam|7355,7358|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|General Exam|7355,7358|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|General Exam|7380,7388|false|false|false|||evaluate
Anatomy|Body Part, Organ, or Organ Component|General Exam|7396,7403|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|General Exam|7396,7403|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|General Exam|7404,7410|false|false|false|||lesion
Finding|Finding|General Exam|7404,7410|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|7404,7410|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|General Exam|7414,7423|false|false|false|||indicated
Anatomy|Body Location or Region|General Exam|7435,7442|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|7435,7442|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|General Exam|7435,7442|false|false|false|||abdomen
Finding|Finding|General Exam|7435,7442|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|General Exam|7450,7461|false|false|false|||Radiographs
Procedure|Diagnostic Procedure|General Exam|7450,7461|false|false|false|C1306645|Plain x-ray|Radiographs
Anatomy|Body Location or Region|General Exam|7469,7476|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|7469,7476|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|7469,7476|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|General Exam|7469,7480|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|General Exam|7469,7487|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|General Exam|7481,7487|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|7481,7487|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|7481,7487|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|7481,7487|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|General Exam|7488,7499|false|false|false|||demonstrate
Anatomy|Body Part, Organ, or Organ Component|General Exam|7517,7522|false|false|false|C0021853|Intestines|bowel
Drug|Biomedical or Dental Material|General Exam|7523,7526|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|General Exam|7523,7526|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|General Exam|7523,7526|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Event|Event|General Exam|7523,7526|false|false|false|||gas
Finding|Gene or Genome|General Exam|7523,7526|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|General Exam|7523,7526|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|General Exam|7523,7526|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|General Exam|7523,7526|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Event|Event|General Exam|7527,7534|false|false|false|||pattern
Attribute|Clinical Attribute|General Exam|7539,7547|false|false|false|C3172260||relative
Finding|Idea or Concept|General Exam|7539,7547|false|false|false|C1546849|Living Arrangement - Relative|relative
Event|Event|General Exam|7548,7555|false|false|false|||paucity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7559,7564|false|false|false|C0021853|Intestines|bowel
Drug|Biomedical or Dental Material|General Exam|7565,7568|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|General Exam|7565,7568|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|General Exam|7565,7568|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Event|Event|General Exam|7565,7568|false|false|false|||gas
Finding|Gene or Genome|General Exam|7565,7568|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|General Exam|7565,7568|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|General Exam|7565,7568|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|General Exam|7565,7568|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Event|Event|General Exam|7572,7579|false|false|false|||present
Finding|Finding|General Exam|7572,7579|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|7572,7579|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Location or Region|General Exam|7598,7609|false|false|false|C0230167|Structure of mid abdomen (surface region)|mid abdomen
Anatomy|Body Location or Region|General Exam|7602,7609|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|7602,7609|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|7602,7609|false|false|false|C0941288|Abdomen problem|abdomen
Finding|Finding|General Exam|7611,7617|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|7611,7617|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Anatomical Abnormality|General Exam|7632,7643|false|false|false|C2711450|Enlargement (morphologic abnormality)|enlargement
Event|Event|General Exam|7632,7643|false|false|false|||enlargement
Finding|Pathologic Function|General Exam|7632,7643|false|false|false|C0020564|Hypertrophy|enlargement
Procedure|Therapeutic or Preventive Procedure|General Exam|7632,7643|false|false|false|C1293134|Enlargement procedure|enlargement
Anatomy|Body Part, Organ, or Organ Component|General Exam|7652,7657|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|7652,7657|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|7652,7657|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|7652,7657|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|7652,7657|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|7652,7657|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|7652,7657|false|false|false|||liver
Finding|Finding|General Exam|7652,7657|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|7652,7657|false|false|false|C0872387|Procedures on liver|liver
Event|Event|General Exam|7659,7669|false|false|false|||displacing
Anatomy|Body Part, Organ, or Organ Component|General Exam|7670,7675|false|false|false|C0021853|Intestines|bowel
Event|Event|General Exam|7676,7681|false|false|false|||loops
Event|Event|General Exam|7684,7688|false|false|false|||Note
Finding|Intellectual Product|General Exam|7698,7705|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|General Exam|7698,7705|false|false|false|C1550585|Entity Handling - upright|upright
Event|Event|General Exam|7707,7711|false|false|false|||view
Event|Event|General Exam|7727,7737|false|false|false|||suboptimal
Event|Event|General Exam|7743,7749|false|false|false|||limits
Finding|Functional Concept|General Exam|7743,7749|false|false|false|C0439801|Limited (extensiveness)|limits
Event|Event|General Exam|7750,7760|false|false|false|||evaluation
Finding|Idea or Concept|General Exam|7750,7760|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|General Exam|7750,7760|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|General Exam|7765,7769|false|false|false|||free
Finding|Functional Concept|General Exam|7765,7769|false|false|false|C0332296|Free of (attribute)|free
Event|Event|General Exam|7771,7786|false|false|false|||intraperitoneal
Finding|Finding|General Exam|7771,7786|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Finding|Functional Concept|General Exam|7771,7786|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Drug|Inorganic Chemical|General Exam|7787,7790|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|7787,7790|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|7787,7790|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|General Exam|7787,7790|false|false|false|||air
Finding|Finding|General Exam|7787,7790|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|7787,7790|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|7787,7790|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Functional Concept|General Exam|7796,7800|false|false|false|C0332296|Free of (attribute)|free
Finding|Finding|General Exam|7801,7816|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Finding|Functional Concept|General Exam|7801,7816|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Drug|Inorganic Chemical|General Exam|7817,7820|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|7817,7820|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|7817,7820|false|true|false|C0001861;C3536832|Air (substance);air|air
Event|Event|General Exam|7817,7820|false|false|false|||air
Finding|Finding|General Exam|7817,7820|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|7817,7820|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|7817,7820|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|General Exam|7824,7833|false|false|false|||suspected
Finding|Functional Concept|General Exam|7849,7853|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|General Exam|7862,7871|false|false|false|C4554531|Pressure injury|decubitus
Event|Event|General Exam|7862,7871|false|false|false|||decubitus
Anatomy|Body Location or Region|General Exam|7884,7891|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|7884,7891|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|7884,7891|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|General Exam|7902,7913|false|false|false|||recommended
Finding|Functional Concept|Hospital Course|7962,7972|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Hospital Course|7962,7979|false|false|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|Hospital Course|7973,7979|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|7973,7979|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7983,7990|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Hospital Course|7983,7990|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Hospital Course|7983,7990|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Hospital Course|7983,7990|false|false|false|||unknown
Finding|Finding|Hospital Course|7983,7990|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Hospital Course|7983,7990|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Hospital Course|7983,7990|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Hospital Course|7983,7990|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|Hospital Course|8011,8018|false|false|false|||lesions
Finding|Finding|Hospital Course|8011,8018|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8026,8031|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8026,8031|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8026,8031|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8026,8031|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8026,8031|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8026,8031|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|8026,8031|false|false|false|||liver
Finding|Finding|Hospital Course|8026,8031|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8026,8031|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8036,8041|false|false|false|C0024109|Lung|lungs
Event|Event|Hospital Course|8058,8067|false|false|false|||presented
Event|Event|Hospital Course|8073,8082|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|8073,8092|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|8073,8092|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|Hospital Course|8086,8092|false|false|false|||breath
Finding|Body Substance|Hospital Course|8086,8092|false|false|false|C0225386|Breath|breath
Finding|Finding|Hospital Course|8094,8100|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8094,8100|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|8108,8117|false|false|false|||worsening
Finding|Idea or Concept|Hospital Course|8108,8117|false|true|false|C1546960|Patient Outcome - Worsening|worsening
Finding|Functional Concept|Hospital Course|8119,8133|false|false|false|C1522224|Intrapulmonary Route of Administration|intrapulmonary
Disorder|Neoplastic Process|Hospital Course|8134,8139|false|false|false|C0027651|Neoplasms|tumor
Event|Event|Hospital Course|8134,8139|false|false|false|||tumor
Finding|Finding|Hospital Course|8134,8139|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|Hospital Course|8134,8139|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Procedure|Diagnostic Procedure|Hospital Course|8134,8146|false|false|false|C1449699|Tumor Burden|tumor burden
Event|Event|Hospital Course|8140,8146|false|false|false|||burden
Finding|Idea or Concept|Hospital Course|8140,8146|false|false|false|C2828008|Burden|burden
Event|Event|Hospital Course|8168,8180|false|false|false|||percutaneous
Finding|Functional Concept|Hospital Course|8168,8180|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8182,8187|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8182,8187|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8182,8187|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8182,8187|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8182,8187|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8182,8187|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|8182,8187|false|false|false|||liver
Finding|Finding|Hospital Course|8182,8187|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8182,8187|false|false|false|C0872387|Procedures on liver|liver
Procedure|Diagnostic Procedure|Hospital Course|8182,8194|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Procedure|Health Care Activity|Hospital Course|8182,8194|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Event|Event|Hospital Course|8188,8194|false|false|false|||biopsy
Finding|Finding|Hospital Course|8188,8194|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|8188,8194|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|8188,8194|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|8188,8194|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|8200,8209|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|8200,8209|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|8200,8209|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|8200,8209|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|8210,8220|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|8210,8220|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|8210,8225|false|false|false|C0332290|Consistent with|consistent with
Finding|Functional Concept|Hospital Course|8226,8236|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8237,8242|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Hospital Course|8237,8242|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Hospital Course|8237,8242|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|Hospital Course|8237,8242|false|false|false|||colon
Finding|Finding|Hospital Course|8237,8242|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Hospital Course|8244,8250|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|8244,8250|false|false|false|||cancer
Event|Event|Hospital Course|8252,8261|false|false|false|||prompting
Event|Event|Hospital Course|8262,8270|false|false|false|||transfer
Finding|Functional Concept|Hospital Course|8262,8270|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|Hospital Course|8262,8270|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|Hospital Course|8262,8270|false|false|false|C4706767|Transfer (immobility management)|transfer
Disorder|Neoplastic Process|Hospital Course|8278,8286|false|false|false|C0027651|Neoplasms|oncology
Event|Event|Hospital Course|8278,8286|false|false|false|||oncology
Procedure|Health Care Activity|Hospital Course|8278,8286|false|false|false|C1555459|oncology services|oncology
Procedure|Health Care Activity|Hospital Course|8278,8294|false|false|false|C1555459|oncology services|oncology service
Event|Occupational Activity|Hospital Course|8287,8294|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|8287,8294|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|8311,8321|false|false|false|||discharged
Event|Event|Hospital Course|8322,8326|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8322,8326|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8322,8326|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8322,8326|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8332,8339|false|false|false|||hospice
Procedure|Health Care Activity|Hospital Course|8332,8339|false|false|false|C0085555|Hospice Care|hospice
Finding|Functional Concept|Hospital Course|8361,8371|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|Hospital Course|8361,8392|false|false|false|C4324497|Adenocarcinoma of colon metastatic|Metastatic colon adenocarcinoma
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8372,8377|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Hospital Course|8372,8377|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Hospital Course|8372,8377|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Hospital Course|8372,8377|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Hospital Course|8372,8392|false|false|false|C0338106|Adenocarcinoma of colon|colon adenocarcinoma
Disorder|Neoplastic Process|Hospital Course|8378,8392|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|8378,8392|false|false|false|||adenocarcinoma
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8394,8397|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|8394,8397|true|false|false|||CTA
Finding|Gene or Genome|Hospital Course|8394,8397|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|8394,8397|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|8401,8408|false|false|false|||exclude
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8409,8418|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|8409,8418|true|true|false|C2707265||pulmonary
Finding|Finding|Hospital Course|8409,8418|true|true|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Hospital Course|8420,8427|true|false|false|||embolus
Finding|Finding|Hospital Course|8420,8427|true|false|false|C1704212;C2046122|Embolus|embolus
Finding|Functional Concept|Hospital Course|8432,8437|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|8432,8452|true|false|false|C0230177|Structure of right upper quadrant of abdomen|right upper quadrant
Event|Event|Hospital Course|8453,8463|false|false|false|||ultrasound
Finding|Functional Concept|Hospital Course|8453,8463|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Hospital Course|8453,8463|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Hospital Course|8453,8463|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|Hospital Course|8467,8476|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8467,8476|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|8478,8490|false|false|false|||demonstrated
Event|Event|Hospital Course|8491,8502|false|false|false|||progression
Finding|Functional Concept|Hospital Course|8491,8502|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|8491,8502|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Event|Event|Hospital Course|8528,8538|false|false|false|||metastatic
Finding|Functional Concept|Hospital Course|8528,8538|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Hospital Course|8540,8546|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|8540,8546|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8550,8557|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Hospital Course|8550,8557|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Hospital Course|8550,8557|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Hospital Course|8550,8557|false|false|false|||unknown
Finding|Finding|Hospital Course|8550,8557|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Hospital Course|8550,8557|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Hospital Course|8550,8557|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Hospital Course|8550,8557|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|Hospital Course|8566,8575|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8580,8585|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8580,8585|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8580,8585|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8580,8585|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8580,8585|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8580,8585|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|8580,8585|false|false|false|||liver
Finding|Finding|Hospital Course|8580,8585|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8580,8585|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8590,8595|false|false|false|C0024109|Lung|lungs
Attribute|Clinical Attribute|Hospital Course|8615,8624|false|false|false|C0945731||diagnosis
Event|Event|Hospital Course|8615,8624|false|false|false|||diagnosis
Finding|Classification|Hospital Course|8615,8624|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|8615,8624|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8615,8624|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Classification|Hospital Course|8632,8642|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8632,8642|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|8643,8650|false|false|false|||setting
Finding|Mental Process|Hospital Course|8643,8650|false|false|false|C0542559|contextual factors|setting
Finding|Body Substance|Hospital Course|8658,8665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8658,8665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8658,8665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|8667,8677|false|false|false|||reluctance
Finding|Mental Process|Hospital Course|8667,8677|false|false|false|C2347948|Reluctance|reluctance
Event|Event|Hospital Course|8681,8687|false|false|false|||engage
Event|Activity|Hospital Course|8693,8697|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|8693,8697|false|false|false|||care
Finding|Finding|Hospital Course|8693,8697|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8693,8697|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Hospital Course|8699,8711|false|false|false|C1522243|Percutaneous Route of Drug Administration|Percutaneous
Procedure|Diagnostic Procedure|Hospital Course|8699,8724|false|false|false|C0558534|Percutaneous liver biopsy|Percutaneous liver biopsy
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8712,8717|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8712,8717|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8712,8717|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8712,8717|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8712,8717|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8712,8717|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|8712,8717|false|false|false|||liver
Finding|Finding|Hospital Course|8712,8717|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8712,8717|false|false|false|C0872387|Procedures on liver|liver
Procedure|Diagnostic Procedure|Hospital Course|8712,8724|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Procedure|Health Care Activity|Hospital Course|8712,8724|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Event|Event|Hospital Course|8718,8724|false|false|false|||biopsy
Finding|Finding|Hospital Course|8718,8724|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|8718,8724|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|8718,8724|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|8718,8724|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|8737,8745|false|false|false|||revealed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8754,8761|false|false|false|C0009368|Colon structure (body structure)|colonic
Disorder|Neoplastic Process|Hospital Course|8754,8776|false|false|false|C0338106|Adenocarcinoma of colon|colonic adenocarcinoma
Disorder|Neoplastic Process|Hospital Course|8762,8776|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|8762,8776|false|false|false|||adenocarcinoma
Event|Event|Hospital Course|8789,8799|false|false|false|||discussion
Finding|Social Behavior|Hospital Course|8789,8799|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8789,8799|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|Hospital Course|8809,8819|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8809,8819|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Neoplastic Process|Hospital Course|8820,8828|false|false|false|C0027651|Neoplasms|oncology
Event|Event|Hospital Course|8820,8828|false|false|false|||oncology
Procedure|Health Care Activity|Hospital Course|8820,8828|false|false|false|C1555459|oncology services|oncology
Event|Event|Hospital Course|8829,8838|false|false|false|||providers
Finding|Functional Concept|Hospital Course|8829,8838|false|false|false|C1138603|Provider|providers
Event|Event|Hospital Course|8849,8860|false|false|false|||transferred
Finding|Idea or Concept|Hospital Course|8868,8877|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|8868,8877|false|false|false|C1555324|inpatient encounter|inpatient
Disorder|Neoplastic Process|Hospital Course|8878,8886|false|false|false|C0027651|Neoplasms|oncology
Event|Event|Hospital Course|8878,8886|false|false|false|||oncology
Procedure|Health Care Activity|Hospital Course|8878,8886|false|false|false|C1555459|oncology services|oncology
Procedure|Health Care Activity|Hospital Course|8878,8894|false|false|false|C1555459|oncology services|oncology service
Event|Event|Hospital Course|8887,8894|false|false|false|||service
Event|Occupational Activity|Hospital Course|8887,8894|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|8887,8894|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|8910,8915|false|false|false|||trial
Procedure|Research Activity|Hospital Course|8910,8915|false|false|false|C0008976|Clinical Trials|trial
Event|Event|Hospital Course|8919,8923|false|false|false|||FLOX
Finding|Body Substance|Hospital Course|8944,8951|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8944,8951|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8944,8951|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|8954,8963|false|false|false|C3641766|Very Poor|very poor
Finding|Intellectual Product|Hospital Course|8959,8963|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|Hospital Course|8964,8974|false|false|false|||functional
Finding|Conceptual Entity|Hospital Course|8964,8974|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|Hospital Course|8964,8974|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Attribute|Clinical Attribute|Hospital Course|8980,8991|false|false|false|C2707262||nutritional
Finding|Finding|Hospital Course|8980,8998|false|false|false|C0392209|Nutritional status|nutritional status
Attribute|Clinical Attribute|Hospital Course|8992,8998|false|false|false|C5889824||status
Event|Event|Hospital Course|8992,8998|false|false|false|||status
Finding|Idea or Concept|Hospital Course|8992,8998|false|false|false|C1546481|What subject filter - Status|status
Attribute|Clinical Attribute|Hospital Course|9001,9006|false|false|false|C2979882||goals
Event|Event|Hospital Course|9001,9006|false|false|false|||goals
Finding|Idea or Concept|Hospital Course|9001,9006|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|Hospital Course|9001,9006|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|Hospital Course|9001,9014|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|Hospital Course|9010,9014|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|9010,9014|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|9010,9014|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Hospital Course|9015,9025|false|false|false|||discussion
Finding|Social Behavior|Hospital Course|9015,9025|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9015,9025|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|Hospital Course|9030,9034|false|false|false|||held
Finding|Body Substance|Hospital Course|9045,9052|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9045,9052|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9045,9052|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|9055,9058|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|9055,9058|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|9055,9058|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Event|Event|Hospital Course|9075,9082|false|false|false|||decided
Event|Event|Hospital Course|9086,9091|false|false|false|||focus
Finding|Functional Concept|Hospital Course|9086,9091|false|false|false|C1285542|Has focus|focus
Attribute|Clinical Attribute|Hospital Course|9093,9098|false|false|false|C2979882||goals
Event|Event|Hospital Course|9093,9098|false|false|false|||goals
Finding|Idea or Concept|Hospital Course|9093,9098|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|Hospital Course|9093,9098|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|Hospital Course|9093,9106|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|Hospital Course|9102,9106|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|9102,9106|false|false|false|||care
Finding|Finding|Hospital Course|9102,9106|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|9102,9106|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|9102,9109|false|false|false|C1555558|care of - AddressPartType|care of
Drug|Organic Chemical|Hospital Course|9110,9117|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|9110,9117|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|Hospital Course|9110,9117|false|false|false|||comfort
Finding|Mental Process|Hospital Course|9110,9117|false|false|false|C1331418|Comfort|comfort
Attribute|Clinical Attribute|Hospital Course|9122,9129|false|false|false|C3854129||symptom
Event|Event|Hospital Course|9122,9129|false|false|false|||symptom
Finding|Sign or Symptom|Hospital Course|9122,9129|false|false|false|C1457887|Symptoms|symptom
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9122,9140|false|false|false|C0030231;C1536570|Palliative Care;Symptom Management|symptom management
Event|Event|Hospital Course|9130,9140|false|false|false|||management
Event|Occupational Activity|Hospital Course|9130,9140|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|9130,9140|false|false|false|C0376636|Disease Management|management
Finding|Body Substance|Hospital Course|9149,9156|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9149,9156|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9149,9156|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|9162,9172|false|false|false|||discharged
Event|Event|Hospital Course|9173,9177|false|false|false|||home
Finding|Idea or Concept|Hospital Course|9173,9177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9173,9177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9173,9177|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|9183,9187|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9183,9187|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9183,9187|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|Hospital Course|9183,9195|false|false|false|C3275086|Home Hospice|home hospice
Event|Event|Hospital Course|9188,9195|false|false|false|||hospice
Procedure|Health Care Activity|Hospital Course|9188,9195|false|false|false|C0085555|Hospice Care|hospice
Finding|Functional Concept|Hospital Course|9203,9207|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9203,9213|false|false|false|C0230426|Structure of left thigh|Left thigh
Anatomy|Body Location or Region|Hospital Course|9208,9213|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Finding|Finding|Hospital Course|9208,9222|false|false|false|C2083469|thigh weakness|thigh weakness
Event|Event|Hospital Course|9214,9222|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|9214,9222|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Hospital Course|9231,9241|false|false|false|||tenderness
Finding|Mental Process|Hospital Course|9231,9241|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Hospital Course|9231,9241|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Hospital Course|9251,9256|false|false|false|||found
Finding|Functional Concept|Hospital Course|9272,9276|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9272,9282|false|false|false|C0230426|Structure of left thigh|left thigh
Anatomy|Body Location or Region|Hospital Course|9277,9282|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Finding|Finding|Hospital Course|9277,9291|false|false|false|C2083469|thigh weakness|thigh weakness
Event|Event|Hospital Course|9283,9291|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|9283,9291|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Hospital Course|9295,9306|false|false|false|||association
Finding|Conceptual Entity|Hospital Course|9295,9306|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Mental Process|Hospital Course|9295,9306|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Social Behavior|Hospital Course|9295,9306|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Phenomenon|Phenomenon or Process|Hospital Course|9295,9306|false|false|false|C0596306|Chemical Association|association
Event|Event|Hospital Course|9329,9339|false|false|false|||tenderness
Finding|Mental Process|Hospital Course|9329,9339|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Hospital Course|9329,9339|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Hospital Course|9351,9361|false|false|false|||chronicity
Finding|Mental Process|Hospital Course|9369,9376|true|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|9381,9390|true|false|false|||preserved
Drug|Biomedical or Dental Material|Hospital Course|9391,9397|true|false|false|C1272938|Rectal Dosage Form|rectal
Finding|Finding|Hospital Course|9391,9397|true|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Finding|Functional Concept|Hospital Course|9391,9397|true|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Event|Event|Hospital Course|9398,9402|true|false|false|||tone
Finding|Sign or Symptom|Hospital Course|9411,9428|true|false|false|C3266098|Numbness of saddle area|saddle anesthesia
Attribute|Clinical Attribute|Hospital Course|9418,9428|true|false|false|C2926599||anesthesia
Drug|Pharmacologic Substance|Hospital Course|9418,9428|true|false|false|C4049933|Anesthesia substance|anesthesia
Event|Event|Hospital Course|9418,9428|true|false|false|||anesthesia
Finding|Finding|Hospital Course|9418,9428|true|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Finding|Sign or Symptom|Hospital Course|9418,9428|true|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9418,9428|true|false|false|C0002903;C0002912|Anesthesia procedures;Dental anesthesia|anesthesia
Event|Event|Hospital Course|9438,9443|false|false|false|||noted
Event|Event|Hospital Course|9451,9462|false|false|false|||incontinent
Finding|Functional Concept|Hospital Course|9451,9462|false|false|false|C0231238|Incontinent|incontinent
Finding|Finding|Hospital Course|9451,9471|false|false|false|C0042024;C2048804|Urinary Incontinence;incontinent of urine on urethra exam|incontinent of urine
Finding|Pathologic Function|Hospital Course|9451,9471|false|false|false|C0042024;C2048804|Urinary Incontinence;incontinent of urine on urethra exam|incontinent of urine
Event|Event|Hospital Course|9466,9471|false|false|false|||urine
Finding|Body Substance|Hospital Course|9466,9471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|9466,9471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|9466,9471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|Hospital Course|9481,9486|true|false|false|||feces
Finding|Body Substance|Hospital Course|9481,9486|true|false|false|C0015733|Feces|feces
Event|Event|Hospital Course|9494,9504|false|false|false|||underlying
Finding|Finding|Hospital Course|9494,9504|false|false|false|C4722602|Underlying|underlying
Disorder|Neoplastic Process|Hospital Course|9506,9516|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|9506,9516|false|false|false|||malignancy
Event|Event|Hospital Course|9528,9535|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|9528,9535|false|false|false|C2699424|Concern|concern
Finding|Functional Concept|Hospital Course|9540,9544|false|false|false|C0443157|Bony|bony
Disorder|Neoplastic Process|Hospital Course|9540,9555|false|false|false|C0153690|Metastatic malignant neoplasm to bone|bony metastases
Disorder|Neoplastic Process|Hospital Course|9545,9555|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|Hospital Course|9545,9555|false|false|false|||metastases
Finding|Finding|Hospital Course|9545,9555|false|false|false|C1513183|Metastatic Lesion|metastases
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9559,9563|false|false|false|C1550235|Cord - Body Parts|cord
Disorder|Disease or Syndrome|Hospital Course|9559,9563|false|true|false|C3489532|Cone-Rod Dystrophy 2|cord
Event|Event|Hospital Course|9559,9563|false|false|false|||cord
Event|Event|Hospital Course|9565,9576|false|false|false|||involvement
Finding|Functional Concept|Hospital Course|9565,9576|false|false|false|C1314939|Involvement with|involvement
Event|Event|Hospital Course|9595,9608|false|false|false|||consideration
Finding|Finding|Hospital Course|9595,9608|false|false|false|C0518609|Consideration|consideration
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9618,9626|false|false|false|C1550254|Body Parts - Epidural|epidural
Finding|Functional Concept|Hospital Course|9618,9626|false|false|false|C0592511|Epidural Route of Administration|epidural
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9618,9626|false|false|false|C0812144||epidural
Disorder|Disease or Syndrome|Hospital Course|9628,9635|false|false|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|9628,9635|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|9628,9635|false|false|false|C1546533||abscess
Event|Event|Hospital Course|9637,9646|false|false|false|||prompting
Finding|Finding|Hospital Course|9647,9656|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Event|Event|Hospital Course|9657,9667|false|false|false|||initiation
Finding|Functional Concept|Hospital Course|9657,9667|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|Hospital Course|9657,9667|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|Hospital Course|9657,9667|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Antibiotic|Hospital Course|9679,9689|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|Hospital Course|9679,9689|false|false|false|||antibiotic
Event|Event|Hospital Course|9691,9699|false|false|false|||coverage
Finding|Functional Concept|Hospital Course|9691,9699|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Idea or Concept|Hospital Course|9691,9699|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Intellectual Product|Hospital Course|9691,9699|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9705,9715|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|9705,9715|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|Hospital Course|9705,9715|false|false|false|||vancomycin
Procedure|Laboratory Procedure|Hospital Course|9705,9715|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|Hospital Course|9716,9723|false|false|false|C0055003|cefepime|cefepim
Drug|Organic Chemical|Hospital Course|9716,9723|false|false|false|C0055003|cefepime|cefepim
Event|Event|Hospital Course|9716,9723|false|false|false|||cefepim
Event|Event|Hospital Course|9765,9772|false|false|false|||efforts
Event|Event|Hospital Course|9778,9786|false|false|false|||declined
Event|Event|Hospital Course|9796,9804|true|false|false|||attempts
Event|Event|Hospital Course|9821,9824|true|false|false|||MRI
Finding|Gene or Genome|Hospital Course|9821,9824|true|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|9821,9824|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|9821,9824|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Drug|Organic Chemical|Hospital Course|9841,9850|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|9841,9850|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|9851,9864|false|false|false|||premedication
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9851,9864|false|false|false|C0033045|Premedication|premedication
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9874,9888|false|false|false|C0008909|Claustrophobia|claustrophobia
Event|Event|Hospital Course|9874,9888|false|false|false|||claustrophobia
Procedure|Diagnostic Procedure|Hospital Course|9890,9900|false|false|false|C0027853|Neurologic Examination|Neuro exam
Event|Event|Hospital Course|9896,9900|false|false|false|||exam
Finding|Functional Concept|Hospital Course|9896,9900|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|9896,9900|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|9905,9914|false|false|false|||monitored
Event|Event|Hospital Course|9919,9927|false|false|false|||remained
Event|Event|Hospital Course|9928,9934|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|9928,9934|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Location or Region|Hospital Course|9941,9950|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Hospital Course|9941,9955|false|false|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Hospital Course|9951,9955|false|false|false|C2598155||pain
Event|Event|Hospital Course|9951,9955|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9951,9955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9951,9955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9973,10000|true|false|false|C0262527|Intermittent abdominal pain|intermittent abdominal pain
Anatomy|Body Location or Region|Hospital Course|9986,9995|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|9986,10000|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|9996,10000|true|false|false|C2598155||pain
Event|Event|Hospital Course|9996,10000|true|false|false|||pain
Finding|Functional Concept|Hospital Course|9996,10000|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9996,10000|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|10006,10016|true|false|false|||tenderness
Finding|Mental Process|Hospital Course|10006,10016|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Hospital Course|10006,10016|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|Hospital Course|10025,10035|true|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|Hospital Course|10025,10035|true|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Event|Event|Hospital Course|10036,10041|true|false|false|||signs
Finding|Finding|Hospital Course|10036,10041|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|10036,10041|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|10059,10070|true|false|false|||obstruction
Finding|Finding|Hospital Course|10059,10070|true|false|false|C0028778|Obstruction|obstruction
Finding|Mental Process|Hospital Course|10078,10085|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Location or Region|Hospital Course|10089,10103|false|false|false|C0230168|Abdominal Cavity|intraabdominal
Disorder|Neoplastic Process|Hospital Course|10104,10114|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|10104,10114|false|false|false|||malignancy
Event|Event|Hospital Course|10136,10144|false|false|false|||episodes
Event|Event|Hospital Course|10148,10154|false|false|false|||emesis
Finding|Body Substance|Hospital Course|10148,10154|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|10148,10154|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|10148,10154|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Event|Event|Hospital Course|10155,10166|false|false|false|||hematemesis
Finding|Sign or Symptom|Hospital Course|10155,10166|false|false|false|C0018926|Hematemesis|hematemesis
Event|Event|Hospital Course|10193,10197|true|false|false|||KUBs
Event|Event|Hospital Course|10203,10211|false|false|false|||negative
Finding|Classification|Hospital Course|10203,10211|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|10203,10211|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|10203,10211|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|10203,10215|false|false|false|C0205160|Negative|negative for
Event|Event|Hospital Course|10216,10227|true|false|false|||obstruction
Finding|Finding|Hospital Course|10216,10227|true|false|false|C0028778|Obstruction|obstruction
Attribute|Clinical Attribute|Hospital Course|10229,10239|true|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|Hospital Course|10229,10239|true|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|Hospital Course|10232,10239|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|10232,10239|true|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|Hospital Course|10232,10239|true|false|false|||abdomen
Finding|Finding|Hospital Course|10232,10239|true|false|false|C0941288|Abdomen problem|abdomen
Event|Event|Hospital Course|10245,10252|false|false|false|||planned
Event|Event|Hospital Course|10256,10264|false|false|false|||evaluate
Event|Event|Hospital Course|10281,10288|false|false|false|||sources
Finding|Finding|Hospital Course|10281,10288|false|false|false|C0449416|Source|sources
Anatomy|Body Location or Region|Hospital Course|10293,10307|false|false|false|C0230168|Abdominal Cavity|intraabdominal
Event|Event|Hospital Course|10308,10317|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|10308,10317|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|10308,10317|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|10308,10317|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|10327,10335|false|false|false|||declined
Event|Event|Hospital Course|10349,10358|true|false|false|||occasions
Attribute|Clinical Attribute|Hospital Course|10360,10364|false|false|false|C2598155||Pain
Event|Event|Hospital Course|10360,10364|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|10360,10364|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|10360,10364|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|Hospital Course|10369,10379|false|false|false|||controlled
Drug|Organic Chemical|Hospital Course|10385,10398|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|10385,10398|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|10385,10398|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|10385,10398|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Organic Chemical|Hospital Course|10403,10411|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|10403,10411|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|10403,10411|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|10403,10411|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Event|Event|Hospital Course|10416,10422|false|false|false|||needed
Finding|Sign or Symptom|Hospital Course|10431,10442|false|false|false|C0018926|Hematemesis|Hematemesis
Finding|Finding|Hospital Course|10462,10468|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Event|Event|Hospital Course|10469,10476|false|false|false|||episode
Finding|Intellectual Product|Hospital Course|10487,10493|false|false|false|C1705102|Volume (publication)|volume
Event|Event|Hospital Course|10494,10500|false|false|false|||emesis
Finding|Body Substance|Hospital Course|10494,10500|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|10494,10500|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|10494,10500|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Disorder|Disease or Syndrome|Hospital Course|10549,10554|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|10549,10554|false|false|false|||blood
Finding|Body Substance|Hospital Course|10549,10554|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Hospital Course|10559,10564|false|false|false|||found
Disorder|Cell or Molecular Dysfunction|Hospital Course|10577,10585|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|10577,10585|false|false|false|||positive
Finding|Classification|Hospital Course|10577,10585|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|10577,10585|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Drug|Food|Hospital Course|10587,10592|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|Hospital Course|10587,10598|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|Hospital Course|10587,10598|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|Hospital Course|10593,10598|false|false|false|||signs
Finding|Finding|Hospital Course|10593,10598|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|10593,10598|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Attribute|Clinical Attribute|Hospital Course|10603,10613|false|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|Hospital Course|10603,10613|false|false|false|||hematocrit
Finding|Finding|Hospital Course|10603,10613|false|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|Hospital Course|10603,10613|false|false|false|C0018935|Hematocrit Measurement|hematocrit
Event|Event|Hospital Course|10615,10623|false|false|false|||remained
Event|Event|Hospital Course|10624,10630|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|10624,10630|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Organic Chemical|Hospital Course|10635,10647|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|Hospital Course|10635,10647|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|Hospital Course|10635,10647|false|false|false|||pantoprazole
Event|Event|Hospital Course|10652,10661|false|false|false|||initiated
Finding|Intellectual Product|Hospital Course|10667,10683|false|false|false|C1314977|Gastrointestinal attachment|gastrointestinal
Event|Event|Hospital Course|10684,10695|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10684,10695|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|10713,10728|true|false|false|||discontinuation
Finding|Finding|Hospital Course|10713,10728|true|false|false|C0457454;C1444662|Discontinuation (procedure);Discontinued|discontinuation
Finding|Functional Concept|Hospital Course|10713,10728|true|false|false|C0457454;C1444662|Discontinuation (procedure);Discontinued|discontinuation
Drug|Pharmacologic Substance|Hospital Course|10733,10736|true|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|Hospital Course|10733,10736|true|false|false|||PPI
Finding|Physiologic Function|Hospital Course|10733,10736|true|false|false|C0871125|Prepulse Inhibition|PPI
Disorder|Neoplastic Process|Hospital Course|10746,10756|true|false|false|C1458156|Recurrent Malignant Neoplasm|recurrence
Event|Event|Hospital Course|10746,10756|true|false|false|||recurrence
Finding|Pathologic Function|Hospital Course|10746,10756|true|false|false|C2825055|Recurrence (disease attribute)|recurrence
Phenomenon|Phenomenon or Process|Hospital Course|10746,10756|true|false|false|C0034897|Recurrence|recurrence
Event|Event|Hospital Course|10761,10773|true|false|false|||questionable
Event|Event|Hospital Course|10783,10790|false|false|false|||episode
Disorder|Disease or Syndrome|Hospital Course|10801,10806|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|10801,10806|false|false|false|||blood
Finding|Body Substance|Hospital Course|10801,10806|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|10811,10814|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|Hospital Course|10811,10814|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Drug|Food|Hospital Course|10815,10823|false|false|false|C3853215|Popsicle|popsicle
Event|Event|Hospital Course|10815,10823|false|false|false|||popsicle
Event|Event|Hospital Course|10828,10834|false|false|false|||eating
Finding|Finding|Hospital Course|10838,10842|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|10838,10842|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|10838,10842|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|10845,10871|false|false|false|||Esophagogastroduodenoscopy
Procedure|Diagnostic Procedure|Hospital Course|10845,10871|false|false|false|C0079304|Esophagogastroduodenoscopy|Esophagogastroduodenoscopy
Event|Event|Hospital Course|10876,10884|false|false|false|||deferred
Disorder|Anatomical Abnormality|Hospital Course|10892,10899|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|Hospital Course|10892,10899|false|false|false|||absence
Finding|Functional Concept|Hospital Course|10892,10899|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|Hospital Course|10892,10902|false|false|false|C0332197|Absent|absence of
Event|Event|Hospital Course|10914,10925|false|false|false|||hematemesis
Finding|Sign or Symptom|Hospital Course|10914,10925|false|false|false|C0018926|Hematemesis|hematemesis
Event|Event|Hospital Course|10936,10940|true|false|false|||EGDs
Procedure|Diagnostic Procedure|Hospital Course|10936,10940|true|false|false|C0079304|Esophagogastroduodenoscopy|EGDs
Event|Event|Hospital Course|10946,10955|true|false|false|||available
Finding|Functional Concept|Hospital Course|10946,10955|true|false|false|C0470187|Availability of|available
Event|Event|Hospital Course|10959,10962|true|false|false|||OMR
Finding|Gene or Genome|Hospital Course|10959,10962|true|false|false|C1412647|ATP5F1A gene|OMR
Finding|Mental Process|Hospital Course|10978,10984|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Hospital Course|10978,10991|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Hospital Course|10978,10991|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Hospital Course|10985,10991|false|false|false|C5889824||status
Event|Event|Hospital Course|10985,10991|false|false|false|||status
Finding|Idea or Concept|Hospital Course|10985,10991|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|11016,11023|true|false|false|||altered
Event|Event|Hospital Course|11036,11045|true|false|false|||admission
Procedure|Health Care Activity|Hospital Course|11036,11045|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|11053,11061|true|false|false|||oriented
Attribute|Clinical Attribute|Hospital Course|11075,11081|true|false|false|C5890614||person
Finding|Intellectual Product|Hospital Course|11075,11081|true|false|false|C1522390|Person Info|person
Event|Activity|Hospital Course|11087,11092|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Hospital Course|11087,11092|false|false|false|||place
Finding|Functional Concept|Hospital Course|11087,11092|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|11087,11092|false|false|false|C1533810||place
Event|Event|Hospital Course|11110,11120|false|false|false|||difficulty
Finding|Finding|Hospital Course|11110,11120|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Gene or Genome|Hospital Course|11131,11137|false|false|false|C1424587|LITAF gene|simple
Event|Event|Hospital Course|11138,11146|false|false|false|||commands
Event|Event|Hospital Course|11151,11159|false|false|false|||compared
Finding|Finding|Hospital Course|11166,11175|false|false|false|C0087130|Uncertainty|uncertain
Drug|Biomedical or Dental Material|Hospital Course|11176,11184|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|11176,11184|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|11176,11184|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Hospital Course|11186,11196|false|false|false|C0009450|Communicable Diseases|Infectious
Event|Event|Hospital Course|11186,11196|false|false|false|||Infectious
Event|Occupational Activity|Hospital Course|11197,11201|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|11197,11204|false|false|false|C0750430|Work-up|work up
Event|Event|Hospital Course|11202,11204|false|false|false|||up
Disorder|Disease or Syndrome|Hospital Course|11217,11222|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|11217,11222|false|false|false|||blood
Finding|Body Substance|Hospital Course|11217,11222|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Hospital Course|11227,11232|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|11227,11232|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|11227,11232|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|Hospital Course|11233,11241|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|11233,11241|false|false|false|C0010453|Culture (Anthropological)|cultures
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11246,11249|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|11246,11249|false|false|false|||CTA
Finding|Gene or Genome|Hospital Course|11246,11249|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|11246,11249|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|11253,11262|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|11253,11262|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|11268,11278|false|false|false|||subsequent
Event|Event|Hospital Course|11280,11284|false|false|false|||CXRs
Event|Event|Hospital Course|11290,11301|false|false|false|||unrevealing
Anatomy|Body Location or Region|Hospital Course|11315,11319|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11315,11319|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|11315,11319|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11315,11319|true|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|Hospital Course|11315,11322|true|false|false|C0202691|CAT scan of head|head CT
Event|Event|Hospital Course|11320,11322|true|false|false|||CT
Event|Event|Hospital Course|11327,11335|false|false|false|||negative
Finding|Classification|Hospital Course|11327,11335|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|11327,11335|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|11327,11335|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|11327,11339|false|false|false|C0205160|Negative|negative for
Finding|Intellectual Product|Hospital Course|11341,11346|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Hospital Course|11347,11359|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Hospital Course|11347,11359|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11360,11367|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|11360,11367|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|11360,11367|true|false|false|||process
Finding|Functional Concept|Hospital Course|11360,11367|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|11360,11367|true|false|false|C1522240|Process|process
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11369,11374|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|Hospital Course|11369,11374|false|false|false|C0006111|Brain Diseases|Brain
Procedure|Diagnostic Procedure|Hospital Course|11369,11378|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|Brain MRI
Event|Event|Hospital Course|11375,11378|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|11375,11378|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|11375,11378|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|11375,11378|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Activity|Hospital Course|11394,11403|true|false|false|C2828389|Exclusion|exclusion
Event|Event|Hospital Course|11394,11403|true|false|false|||exclusion
Finding|Functional Concept|Hospital Course|11394,11403|true|false|false|C0680251|Exclusion Criteria|exclusion
Disorder|Neoplastic Process|Hospital Course|11408,11418|true|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|Hospital Course|11408,11418|true|false|false|||metastases
Finding|Finding|Hospital Course|11408,11418|true|false|false|C1513183|Metastatic Lesion|metastases
Event|Event|Hospital Course|11432,11440|true|false|false|||obtained
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11448,11462|true|false|false|C0008909|Claustrophobia|claustrophobia
Event|Event|Hospital Course|11448,11462|true|false|false|||claustrophobia
Event|Event|Hospital Course|11463,11466|true|false|false|||MRI
Finding|Gene or Genome|Hospital Course|11463,11466|true|true|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|11463,11466|true|true|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|11463,11466|true|true|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Drug|Organic Chemical|Hospital Course|11468,11476|false|false|false|C2825146|Aversion|aversion
Drug|Pharmacologic Substance|Hospital Course|11468,11476|false|false|false|C2825146|Aversion|aversion
Event|Event|Hospital Course|11468,11476|false|false|false|||aversion
Finding|Mental Process|Hospital Course|11468,11476|false|false|false|C0233496|Aversion (finding)|aversion
Finding|Idea or Concept|Hospital Course|11480,11485|false|false|false|C1552828|Table Frame - above|above
Event|Event|Hospital Course|11488,11491|true|false|false|||ABG
Finding|Gene or Genome|Hospital Course|11488,11491|true|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|Hospital Course|11488,11491|true|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Event|Event|Hospital Course|11507,11512|true|false|false|||signs
Finding|Finding|Hospital Course|11507,11512|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|11507,11512|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Drug|Biologically Active Substance|Hospital Course|11516,11519|true|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|Hospital Course|11516,11519|true|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|Hospital Course|11516,11519|true|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|Hospital Course|11516,11519|true|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Finding|Hospital Course|11516,11529|true|false|false|C0020440|Hypercapnia|CO2 retention
Attribute|Clinical Attribute|Hospital Course|11520,11529|true|false|false|C1318143|Retention - dental|retention
Event|Event|Hospital Course|11520,11529|true|false|false|||retention
Finding|Cell Function|Hospital Course|11520,11529|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|Hospital Course|11520,11529|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|Hospital Course|11520,11529|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Event|Event|Hospital Course|11532,11539|false|false|false|||History
Finding|Conceptual Entity|Hospital Course|11532,11539|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|11532,11539|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|11532,11539|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|11532,11542|false|false|false|C0262926|Medical History|History of
Drug|Hazardous or Poisonous Substance|Hospital Course|11543,11550|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Organic Chemical|Hospital Course|11543,11550|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Pharmacologic Substance|Hospital Course|11543,11550|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Event|Event|Hospital Course|11543,11550|false|false|false|||opiates
Procedure|Laboratory Procedure|Hospital Course|11543,11550|false|false|false|C0242401|Opiate Measurement|opiates
Event|Event|Hospital Course|11551,11557|false|false|false|||making
Finding|Body Substance|Hospital Course|11558,11565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11558,11565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11558,11565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|11566,11572|false|false|false|||sleepy
Finding|Finding|Hospital Course|11566,11572|false|false|false|C0013144|Drowsiness|sleepy
Disorder|Disease or Syndrome|Hospital Course|11577,11580|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|11577,11580|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|11577,11580|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Event|Event|Hospital Course|11584,11592|false|false|false|||possible
Finding|Finding|Hospital Course|11584,11592|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|11607,11613|false|false|false|||factor
Finding|Conceptual Entity|Hospital Course|11607,11613|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|Hospital Course|11607,11613|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Intellectual Product|Hospital Course|11607,11613|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Event|Event|Hospital Course|11639,11651|false|false|false|||discontinued
Anatomy|Body Location or Region|Hospital Course|11654,11661|false|false|false|C0205054|Hepatic|Hepatic
Disorder|Disease or Syndrome|Hospital Course|11654,11676|false|false|false|C0019151|Hepatic Encephalopathy|Hepatic encephalopathy
Disorder|Disease or Syndrome|Hospital Course|11662,11676|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|Hospital Course|11662,11676|false|false|false|||encephalopathy
Event|Event|Hospital Course|11685,11697|false|false|false|||differential
Finding|Idea or Concept|Hospital Course|11685,11697|false|false|false|C1549478|Amount type - Differential|differential
Event|Event|Hospital Course|11704,11714|false|false|false|||metastatic
Finding|Functional Concept|Hospital Course|11704,11714|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Event|Event|Hospital Course|11716,11723|false|false|false|||lesions
Finding|Finding|Hospital Course|11716,11723|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11727,11732|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|11727,11732|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|11727,11732|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|11727,11732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|11727,11732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|11727,11732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|11727,11732|false|false|false|||liver
Finding|Finding|Hospital Course|11727,11732|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|11727,11732|false|false|false|C0872387|Procedures on liver|liver
Event|Event|Hospital Course|11737,11746|false|false|false|||asterixis
Finding|Sign or Symptom|Hospital Course|11737,11746|false|false|false|C0232766|Asterixis|asterixis
Event|Event|Hospital Course|11750,11754|false|false|false|||exam
Finding|Functional Concept|Hospital Course|11750,11754|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|11750,11754|false|false|false|C0582103|Medical Examination|exam
Disorder|Disease or Syndrome|Hospital Course|11757,11760|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Event|Event|Hospital Course|11757,11760|false|false|false|||AMS
Finding|Gene or Genome|Hospital Course|11757,11760|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|Hospital Course|11757,11760|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Finding|Finding|Hospital Course|11783,11789|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|11783,11789|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11783,11800|false|false|false|C0588008|Severe depression|severe depression
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11790,11800|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|11790,11800|false|false|false|||depression
Finding|Functional Concept|Hospital Course|11790,11800|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|11790,11800|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Mental Process|Hospital Course|11802,11808|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Hospital Course|11802,11815|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|Hospital Course|11802,11815|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|Hospital Course|11809,11815|false|false|false|C5889824||status
Event|Event|Hospital Course|11809,11815|false|false|false|||status
Finding|Idea or Concept|Hospital Course|11809,11815|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|11816,11825|false|false|false|||monitored
Event|Event|Hospital Course|11830,11838|false|false|false|||remained
Event|Event|Hospital Course|11840,11846|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|11840,11846|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Body Substance|Hospital Course|11851,11858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11851,11858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11851,11858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Biomedical or Dental Material|Hospital Course|11862,11870|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|11862,11870|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|11862,11870|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Hospital Course|11875,11878|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|11875,11878|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|11875,11878|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Event|Event|Hospital Course|11882,11891|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11882,11891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11882,11891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11882,11891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11882,11891|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|11898,11907|false|false|false|||Shortness
Attribute|Clinical Attribute|Hospital Course|11898,11917|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Hospital Course|11898,11917|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Hospital Course|11911,11917|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|11923,11932|false|false|false|||presented
Finding|Intellectual Product|Hospital Course|11938,11943|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|11938,11949|true|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|Hospital Course|11944,11949|true|false|false|||onset
Event|Event|Hospital Course|11951,11960|true|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|11951,11970|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|11951,11970|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|11964,11970|true|false|false|C0225386|Breath|breath
Disorder|Disease or Syndrome|Hospital Course|11979,11984|true|false|false|C0398650|Immune thrombocytopenic purpura|frank
Event|Event|Hospital Course|11985,11992|true|false|false|||hypoxia
Finding|Finding|Hospital Course|11985,11992|true|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|Hospital Course|11985,11992|true|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11994,11997|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|11994,11997|true|false|false|||CTA
Finding|Gene or Genome|Hospital Course|11994,11997|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|11994,11997|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|12001,12010|true|false|false|||admission
Procedure|Health Care Activity|Hospital Course|12001,12010|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|12016,12024|false|false|false|||negative
Finding|Classification|Hospital Course|12016,12024|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|12016,12024|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|12016,12024|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|12016,12028|false|false|false|C0205160|Negative|negative for
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12029,12038|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|12029,12038|true|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|12029,12038|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|12029,12046|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolus
Event|Event|Hospital Course|12039,12046|true|false|false|||embolus
Finding|Finding|Hospital Course|12039,12046|true|false|false|C1704212;C2046122|Embolus|embolus
Drug|Organic Chemical|Hospital Course|12069,12073|true|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Hospital Course|12069,12073|true|false|false|C0009074|clotrimazole|clot
Event|Event|Hospital Course|12069,12073|true|false|false|||clot
Finding|Pathologic Function|Hospital Course|12069,12073|true|false|false|C0302148|Blood Clot|clot
Event|Event|Hospital Course|12088,12096|true|false|false|||excluded
Anatomy|Tissue|Hospital Course|12112,12119|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|12112,12119|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|Hospital Course|12112,12128|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|Hospital Course|12112,12128|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|Hospital Course|12112,12128|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|Hospital Course|12120,12128|false|false|false|||effusion
Finding|Body Substance|Hospital Course|12120,12128|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Hospital Course|12120,12128|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Hospital Course|12120,12128|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|Hospital Course|12133,12138|false|false|false|||focal
Event|Event|Hospital Course|12140,12150|false|false|false|||infiltrate
Finding|Functional Concept|Hospital Course|12140,12150|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Hospital Course|12140,12150|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Hospital Course|12140,12150|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|Hospital Course|12152,12155|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|12152,12155|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|12152,12155|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12160,12167|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|12160,12167|false|false|false|C1314974|Cardiac attachment|cardiac
Attribute|Clinical Attribute|Hospital Course|12160,12175|false|false|false|C2926589||cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12160,12175|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Drug|Enzyme|Hospital Course|12160,12175|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Procedure|Laboratory Procedure|Hospital Course|12160,12175|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12168,12175|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|Hospital Course|12168,12175|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|Hospital Course|12168,12175|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Event|Event|Hospital Course|12168,12175|false|false|false|||enzymes
Finding|Functional Concept|Hospital Course|12168,12175|false|false|false|C0014445|enzymology|enzymes
Event|Event|Hospital Course|12181,12191|false|false|false|||reassuring
Finding|Intellectual Product|Hospital Course|12201,12206|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|12201,12224|false|false|false|C0948089|Acute Coronary Syndrome|acute coronary syndrome
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12207,12215|false|false|false|C0018787|Heart|coronary
Disorder|Disease or Syndrome|Hospital Course|12216,12224|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|12216,12224|false|false|false|||syndrome
Finding|Finding|Hospital Course|12227,12230|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Hospital Course|12227,12230|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Event|Event|Hospital Course|12231,12239|false|false|false|||voltages
Event|Event|Hospital Course|12243,12246|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|12243,12246|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|12243,12246|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|12252,12262|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|12252,12262|false|false|false|C0332290|Consistent with|consistent
Event|Event|Hospital Course|12282,12289|false|false|false|||limited
Finding|Functional Concept|Hospital Course|12282,12289|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|Hospital Course|12282,12289|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Event|Event|Hospital Course|12290,12299|false|false|false|||suspicion
Finding|Mental Process|Hospital Course|12290,12299|false|false|false|C0242114|Suspicion|suspicion
Anatomy|Body Location or Region|Hospital Course|12304,12315|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12304,12315|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Hospital Course|12304,12324|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Hospital Course|12304,12324|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|Hospital Course|12316,12324|false|false|false|||effusion
Finding|Body Substance|Hospital Course|12316,12324|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Hospital Course|12316,12324|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Hospital Course|12316,12324|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|Hospital Course|12327,12336|false|false|false|||Shortness
Attribute|Clinical Attribute|Hospital Course|12327,12346|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Hospital Course|12327,12346|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Hospital Course|12340,12346|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|12347,12355|true|false|false|||resolved
Event|Event|Hospital Course|12375,12384|true|false|false|||admission
Procedure|Health Care Activity|Hospital Course|12375,12384|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|12404,12413|true|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|12404,12413|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|12404,12413|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|12404,12413|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12404,12413|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|12424,12433|true|false|false|||exception
Finding|Conceptual Entity|Hospital Course|12424,12433|true|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Idea or Concept|Hospital Course|12424,12433|true|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Drug|Pharmacologic Substance|Hospital Course|12437,12447|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Hospital Course|12437,12447|false|false|false|||nebulizers
Disorder|Injury or Poisoning|Hospital Course|12453,12465|false|false|false|C0161635;C0851326;C2880043|Expectorants causing adverse effects in therapeutic use;Poisoning by expectorant;Poisoning by, adverse effect of and underdosing of expectorants|expectorants
Drug|Pharmacologic Substance|Hospital Course|12453,12465|false|false|false|C0015314|Expectorants|expectorants
Event|Event|Hospital Course|12453,12465|false|false|false|||expectorants
Event|Event|Hospital Course|12469,12475|false|false|false|||needed
Disorder|Disease or Syndrome|Hospital Course|12482,12494|false|false|false|C0023518|Leukocytosis|Leukocytosis
Event|Event|Hospital Course|12482,12494|false|false|false|||Leukocytosis
Finding|Finding|Hospital Course|12482,12494|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Anatomy|Cell|Hospital Course|12496,12512|false|false|false|C0023516|Leukocytes|White blood cell
Lab|Laboratory or Test Result|Hospital Course|12496,12518|false|false|false|C0427512||White blood cell count
Procedure|Laboratory Procedure|Hospital Course|12496,12518|false|false|false|C0023508|White Blood Cell Count procedure|White blood cell count
Disorder|Disease or Syndrome|Hospital Course|12502,12507|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|12502,12507|false|false|false|||blood
Finding|Body Substance|Hospital Course|12502,12507|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|Hospital Course|12502,12512|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|Hospital Course|12502,12518|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|Hospital Course|12508,12512|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|12508,12512|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|Hospital Course|12508,12518|false|false|false|C0007584|Cell Count|cell count
Event|Event|Hospital Course|12513,12518|false|false|false|||count
Event|Event|Hospital Course|12523,12531|false|false|false|||elevated
Event|Event|Hospital Course|12536,12542|false|false|false|||peaked
Event|Event|Hospital Course|12553,12563|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|12553,12563|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|12553,12568|false|false|false|C0332290|Consistent with|consistent with
Drug|Biomedical or Dental Material|Hospital Course|12576,12584|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|12576,12584|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|12576,12584|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|12586,12592|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|12586,12592|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|12593,12603|false|false|false|||reflecting
Disorder|Neoplastic Process|Hospital Course|12616,12626|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|12616,12626|false|false|false|||malignancy
Event|Event|Hospital Course|12631,12636|false|false|false|||noted
Finding|Idea or Concept|Hospital Course|12637,12642|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|Hospital Course|12644,12654|false|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Hospital Course|12644,12654|false|false|false|||infectious
Event|Occupational Activity|Hospital Course|12655,12659|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|12655,12662|false|false|false|C0750430|Work-up|work up
Event|Event|Hospital Course|12660,12662|false|false|false|||up
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12674,12677|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|12674,12677|false|false|false|||CTA
Finding|Gene or Genome|Hospital Course|12674,12677|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|12674,12677|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|12679,12684|false|false|false|||urine
Finding|Body Substance|Hospital Course|12679,12684|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|12679,12684|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|12679,12684|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Disorder|Disease or Syndrome|Hospital Course|12689,12694|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|12689,12694|false|false|false|||blood
Finding|Body Substance|Hospital Course|12689,12694|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Hospital Course|12689,12703|false|false|false|C0200949|Blood culture|blood cultures
Event|Event|Hospital Course|12695,12703|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|12695,12703|false|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|Hospital Course|12709,12713|false|false|false|||CXRs
Event|Event|Hospital Course|12720,12731|false|false|false|||unrevealing
Event|Event|Hospital Course|12737,12745|false|false|false|||remained
Event|Event|Hospital Course|12746,12754|false|false|false|||afebrile
Finding|Finding|Hospital Course|12746,12754|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|12765,12774|false|false|false|||exception
Finding|Conceptual Entity|Hospital Course|12765,12774|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Idea or Concept|Hospital Course|12765,12774|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Event|Event|Hospital Course|12779,12787|false|false|false|||isolated
Finding|Functional Concept|Hospital Course|12779,12787|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Hospital Course|12779,12787|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Finding|Hospital Course|12788,12797|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Event|Event|Hospital Course|12798,12803|false|false|false|||fever
Finding|Finding|Hospital Course|12798,12803|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|12798,12803|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Hospital Course|12817,12823|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|12817,12823|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|Hospital Course|12824,12829|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|12824,12835|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|12824,12835|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|12830,12835|false|false|false|||signs
Finding|Finding|Hospital Course|12830,12835|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|12830,12835|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12843,12848|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|Hospital Course|12843,12848|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|Hospital Course|12843,12848|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|Hospital Course|12843,12848|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|Hospital Course|12843,12848|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|Hospital Course|12843,12848|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Finding|Finding|Hospital Course|12843,12848|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|Hospital Course|12843,12848|false|false|false|C0872387|Procedures on liver|Liver
Finding|Organ or Tissue Function|Hospital Course|12843,12857|false|false|false|C0232741|Liver function|Liver function
Procedure|Laboratory Procedure|Hospital Course|12843,12862|false|false|false|C0023901|Liver Function Tests|Liver function test
Event|Event|Hospital Course|12849,12857|false|false|false|||function
Finding|Finding|Hospital Course|12849,12857|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|12849,12857|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|12849,12857|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|12849,12857|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Procedure|Diagnostic Procedure|Hospital Course|12849,12862|false|false|false|C5670437|Function Test|function test
Anatomy|Body Location or Region|Hospital Course|12858,12862|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Hospital Course|12858,12862|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|12858,12862|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|12858,12862|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|12858,12862|false|false|false|C0022885|Laboratory Procedures|test
Disorder|Congenital Abnormality|Hospital Course|12863,12876|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Hospital Course|12863,12876|false|false|false|||abnormalities
Finding|Functional Concept|Hospital Course|12863,12876|false|false|false|C0000769|teratologic|abnormalities
Anatomy|Body Space or Junction|Hospital Course|12878,12881|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|Hospital Course|12878,12881|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12878,12881|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|Hospital Course|12878,12881|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|Hospital Course|12878,12881|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|Hospital Course|12878,12881|false|false|false|||AST
Finding|Gene or Genome|Hospital Course|12878,12881|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Event|Event|Hospital Course|12882,12890|false|false|false|||remained
Event|Event|Hospital Course|12891,12899|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12913,12933|false|false|false|C0002059|Alkaline Phosphatase|alkaline phosphatase
Drug|Enzyme|Hospital Course|12913,12933|false|false|false|C0002059|Alkaline Phosphatase|alkaline phosphatase
Finding|Physiologic Function|Hospital Course|12913,12933|false|false|false|C4553029|Alkaline phosphatase metabolic function|alkaline phosphatase
Procedure|Laboratory Procedure|Hospital Course|12913,12933|false|false|false|C0201850|Alkaline phosphatase measurement|alkaline phosphatase
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12922,12933|false|false|false|C0031678|Phosphoric Monoester Hydrolases|phosphatase
Drug|Enzyme|Hospital Course|12922,12933|false|false|false|C0031678|Phosphoric Monoester Hydrolases|phosphatase
Event|Event|Hospital Course|12922,12933|false|false|false|||phosphatase
Finding|Molecular Function|Hospital Course|12922,12933|false|false|false|C1149880|phosphoric monoester hydrolase activity|phosphatase
Event|Event|Hospital Course|12934,12938|false|false|false|||260s
Drug|Biologically Active Substance|Hospital Course|12952,12967|false|false|false|C0005437|Bilirubin|total bilirubin
Drug|Organic Chemical|Hospital Course|12952,12967|false|false|false|C0005437|Bilirubin|total bilirubin
Finding|Physiologic Function|Hospital Course|12952,12967|false|false|false|C4553024|Total bilirubin metabolic function|total bilirubin
Lab|Laboratory or Test Result|Hospital Course|12952,12967|false|false|false|C0368753|Total bilirubin level|total bilirubin
Procedure|Laboratory Procedure|Hospital Course|12952,12967|false|false|false|C0201913|Bilirubin, total measurement|total bilirubin
Drug|Biologically Active Substance|Hospital Course|12958,12967|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Organic Chemical|Hospital Course|12958,12967|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Pharmacologic Substance|Hospital Course|12958,12967|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Event|Event|Hospital Course|12958,12967|false|false|false|||bilirubin
Procedure|Laboratory Procedure|Hospital Course|12958,12967|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|bilirubin
Finding|Finding|Hospital Course|12981,12987|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|12981,12987|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Location or Region|Hospital Course|12995,13002|false|false|false|C0205054|Hepatic|hepatic
Event|Event|Hospital Course|13003,13015|false|false|false|||infiltration
Finding|Functional Concept|Hospital Course|13003,13015|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|Hospital Course|13003,13015|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13003,13015|false|false|false|C0702249|Infiltration (procedure)|infiltration
Disorder|Neoplastic Process|Hospital Course|13019,13029|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|13019,13029|false|false|false|||malignancy
Finding|Functional Concept|Hospital Course|13032,13037|true|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|Hospital Course|13032,13052|true|false|false|C0230177|Structure of right upper quadrant of abdomen|Right upper quadrant
Event|Event|Hospital Course|13053,13063|true|false|false|||ultrasound
Finding|Functional Concept|Hospital Course|13053,13063|true|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Hospital Course|13053,13063|true|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Hospital Course|13053,13063|true|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|Hospital Course|13068,13076|false|false|false|||negative
Finding|Classification|Hospital Course|13068,13076|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|13068,13076|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|13068,13076|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|13068,13080|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|Hospital Course|13081,13094|true|false|false|C0008325|Cholecystitis|cholecystitis
Event|Event|Hospital Course|13081,13094|true|false|false|||cholecystitis
Event|Event|Hospital Course|13099,13110|true|false|false|||obstructive
Finding|Functional Concept|Hospital Course|13099,13110|true|false|false|C0549186|Obstructed|obstructive
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13111,13118|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|13111,13118|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|13111,13118|true|false|false|||process
Finding|Functional Concept|Hospital Course|13111,13118|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|13111,13118|true|false|false|C1522240|Process|process
Event|Event|Hospital Course|13139,13151|false|false|false|||superimposed
Anatomy|Body Location or Region|Hospital Course|13153,13167|false|false|false|C0230168|Abdominal Cavity|intraabdominal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13168,13175|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|13168,13175|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|13168,13175|true|false|false|||process
Finding|Functional Concept|Hospital Course|13168,13175|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|13168,13175|true|false|false|C1522240|Process|process
Disorder|Disease or Syndrome|Hospital Course|13185,13194|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|13185,13194|true|false|false|||infection
Finding|Pathologic Function|Hospital Course|13185,13194|true|false|false|C3714514|Infection|infection
Event|Event|Hospital Course|13209,13217|true|false|false|||excluded
Finding|Mental Process|Hospital Course|13226,13233|true|false|false|C0542559|contextual factors|setting
Anatomy|Body Location or Region|Hospital Course|13237,13246|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|13237,13251|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|13247,13251|true|false|false|C2598155||pain
Event|Event|Hospital Course|13247,13251|true|false|false|||pain
Finding|Functional Concept|Hospital Course|13247,13251|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|13247,13251|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|13257,13263|false|false|false|||emesis
Finding|Body Substance|Hospital Course|13257,13263|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|13257,13263|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|13257,13263|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Idea or Concept|Hospital Course|13267,13272|false|false|false|C1552828|Table Frame - above|above
Event|Event|Hospital Course|13283,13291|false|false|false|||declined
Event|Event|Hospital Course|13292,13294|true|false|false|||CT
Event|Event|Hospital Course|13307,13317|true|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|13307,13317|true|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|13307,13317|true|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|Hospital Course|13324,13340|false|false|false|C4054756|Elevated lactate level|Elevated lactate
Drug|Organic Chemical|Hospital Course|13333,13340|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|Hospital Course|13333,13340|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|Hospital Course|13333,13340|false|false|false|||lactate
Procedure|Laboratory Procedure|Hospital Course|13333,13340|false|false|false|C0202115|Lactic acid measurement|lactate
Drug|Organic Chemical|Hospital Course|13342,13349|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|Hospital Course|13342,13349|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|Hospital Course|13342,13349|false|false|false|||Lactate
Procedure|Laboratory Procedure|Hospital Course|13342,13349|false|false|false|C0202115|Lactic acid measurement|Lactate
Event|Event|Hospital Course|13354,13359|false|false|false|||found
Event|Event|Hospital Course|13386,13395|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|13386,13395|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|13404,13411|false|false|false|C3845930|Copious|copious
Drug|Substance|Hospital Course|13415,13421|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|13415,13421|false|false|false|||fluids
Finding|Body Substance|Hospital Course|13415,13421|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13415,13421|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Finding|Hospital Course|13423,13429|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|13423,13429|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|13430,13440|false|false|false|||reflecting
Finding|Mental Process|Hospital Course|13430,13440|false|true|false|C0558058|Reflecting|reflecting
Event|Event|Hospital Course|13442,13453|false|false|false|||compromised
Anatomy|Body Location or Region|Hospital Course|13454,13461|false|false|false|C0205054|Hepatic|hepatic
Attribute|Clinical Attribute|Hospital Course|13462,13471|false|false|false|C1382187|Clearance of substance|clearance
Event|Event|Hospital Course|13462,13471|false|false|false|||clearance
Phenomenon|Natural Phenomenon or Process|Hospital Course|13462,13471|false|false|false|C2825073|Clearance [PK]|clearance
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13462,13471|false|false|false|C4554548|Clearance procedure|clearance
Finding|Mental Process|Hospital Course|13479,13486|false|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|13501,13513|false|false|false|||infiltration
Finding|Functional Concept|Hospital Course|13501,13513|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|Hospital Course|13501,13513|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13501,13513|false|false|false|C0702249|Infiltration (procedure)|infiltration
Anatomy|Body Space or Junction|Hospital Course|13522,13527|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|Hospital Course|13522,13527|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|Hospital Course|13522,13527|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|Hospital Course|13522,13527|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Disorder|Disease or Syndrome|Hospital Course|13522,13539|false|false|false|C0039239|Sinus Tachycardia|Sinus tachycardia
Finding|Finding|Hospital Course|13522,13539|false|false|false|C2108109;C5235163|Sinus Tachycardia by ECG Finding;continuous electrocardiogram sinus tachycardia|Sinus tachycardia
Event|Event|Hospital Course|13528,13539|false|false|false|||tachycardia
Finding|Finding|Hospital Course|13528,13539|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Hospital Course|13545,13553|false|false|false|||remained
Finding|Idea or Concept|Hospital Course|13554,13566|false|false|false|C0750508|persistently|persistently
Event|Event|Hospital Course|13567,13578|false|false|false|||tachycardic
Event|Event|Hospital Course|13604,13613|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|13604,13613|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Mental Process|Hospital Course|13621,13628|false|false|false|C0542559|contextual factors|setting
Finding|Intellectual Product|Hospital Course|13632,13636|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|Hospital Course|13637,13639|false|false|false|||PO
Event|Event|Hospital Course|13641,13647|false|false|false|||intake
Finding|Functional Concept|Hospital Course|13641,13647|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|13641,13647|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|Hospital Course|13666,13676|false|false|false|||responsive
Finding|Functional Concept|Hospital Course|13666,13676|false|false|false|C0205342|Responsive|responsive
Finding|Finding|Hospital Course|13680,13687|false|false|false|C3845930|Copious|copious
Drug|Substance|Hospital Course|13691,13697|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|13691,13697|false|false|false|||fluids
Finding|Body Substance|Hospital Course|13691,13697|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13691,13697|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Hospital Course|13700,13711|false|false|false|||Tachycardia
Finding|Finding|Hospital Course|13700,13711|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|Tachycardia
Event|Event|Hospital Course|13721,13728|false|false|false|||present
Finding|Finding|Hospital Course|13721,13728|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Hospital Course|13721,13728|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Disease or Syndrome|Hospital Course|13769,13781|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Hospital Course|13769,13781|true|false|false|||leukocytosis
Finding|Finding|Hospital Course|13769,13781|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Finding|Hospital Course|13786,13802|true|false|false|C4054756|Elevated lactate level|elevated lactate
Drug|Organic Chemical|Hospital Course|13795,13802|true|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|Hospital Course|13795,13802|true|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|Hospital Course|13795,13802|true|false|false|||lactate
Procedure|Laboratory Procedure|Hospital Course|13795,13802|true|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|Hospital Course|13817,13822|true|false|false|||clear
Finding|Idea or Concept|Hospital Course|13817,13822|true|false|false|C1550016|Remote control command - Clear|clear
Disorder|Disease or Syndrome|Hospital Course|13824,13834|true|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Hospital Course|13835,13841|true|false|false|||source
Finding|Finding|Hospital Course|13835,13841|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|Hospital Course|13835,13841|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|Hospital Course|13835,13841|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Finding|Hospital Course|13849,13852|true|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|13849,13852|true|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Hospital Course|13853,13862|false|false|false|||suspicion
Finding|Mental Process|Hospital Course|13853,13862|false|false|false|C0242114|Suspicion|suspicion
Disorder|Disease or Syndrome|Hospital Course|13867,13873|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|Hospital Course|13867,13873|false|false|false|||sepsis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13889,13898|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|13889,13898|true|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|13889,13898|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|13889,13906|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolus
Event|Event|Hospital Course|13899,13906|true|false|false|||embolus
Finding|Finding|Hospital Course|13899,13906|true|false|false|C1704212;C2046122|Embolus|embolus
Event|Event|Hospital Course|13920,13928|true|false|false|||excluded
Drug|Pharmacologic Substance|Hospital Course|13936,13941|true|false|false|C1874451|Basis|basis
Finding|Functional Concept|Hospital Course|13936,13941|true|false|false|C1527178|Basis - conceptual entity|basis
Event|Event|Hospital Course|13946,13955|true|false|false|||admission
Procedure|Health Care Activity|Hospital Course|13946,13955|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13956,13959|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|13956,13959|true|false|false|||CTA
Finding|Gene or Genome|Hospital Course|13956,13959|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|13956,13959|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|13965,13974|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|13965,13984|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|13965,13984|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|13978,13984|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|13995,14000|false|false|false|||lived
Event|Event|Hospital Course|14021,14028|true|false|false|||hypoxic
Finding|Pathologic Function|Hospital Course|14021,14028|true|false|false|C0242184|Hypoxia|hypoxic
Attribute|Clinical Attribute|Hospital Course|14030,14040|true|false|false|C1542366|hematocrit attribute|Hematocrit
Event|Event|Hospital Course|14030,14040|true|false|false|||Hematocrit
Finding|Finding|Hospital Course|14030,14040|true|false|false|C0518014|Hematocrit level|Hematocrit
Procedure|Laboratory Procedure|Hospital Course|14030,14040|true|false|false|C0018935|Hematocrit Measurement|Hematocrit
Event|Event|Hospital Course|14050,14056|true|false|false|||stable
Finding|Intellectual Product|Hospital Course|14050,14056|true|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|14065,14070|true|false|false|||signs
Finding|Finding|Hospital Course|14065,14070|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|14065,14070|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|14082,14090|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|14082,14090|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|14101,14110|false|false|false|||exception
Finding|Conceptual Entity|Hospital Course|14101,14110|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Idea or Concept|Hospital Course|14101,14110|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Finding|Hospital Course|14114,14123|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Event|Event|Hospital Course|14124,14135|false|false|false|||hematemesis
Finding|Sign or Symptom|Hospital Course|14124,14135|false|false|false|C0018926|Hematemesis|hematemesis
Finding|Idea or Concept|Hospital Course|14140,14145|false|false|false|C1552828|Table Frame - above|above
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14153,14163|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|Hospital Course|14153,14163|false|false|false|||Depression
Finding|Functional Concept|Hospital Course|14153,14163|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|Hospital Course|14153,14163|false|false|false|C0460137;C1579931|Depression - motion|Depression
Event|Event|Hospital Course|14169,14177|false|false|false|||appeared
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14178,14187|false|false|false|C0344315|Depressed mood|depressed
Event|Event|Hospital Course|14178,14187|false|false|false|||depressed
Finding|Finding|Hospital Course|14193,14204|false|false|false|C0233471|Flat affect|flat affect
Event|Event|Hospital Course|14198,14204|false|false|false|||affect
Finding|Mental Process|Hospital Course|14198,14204|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Hospital Course|14198,14204|false|false|false|C2237113|assessment of affect|affect
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14218,14227|false|false|false|C0178417|Anhedonia|anhedonia
Event|Event|Hospital Course|14218,14227|false|false|false|||anhedonia
Event|Event|Hospital Course|14239,14248|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|14239,14248|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|14255,14265|false|false|false|||underlying
Finding|Finding|Hospital Course|14255,14265|false|false|false|C4722602|Underlying|underlying
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14267,14277|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|14267,14277|false|false|false|||depression
Finding|Functional Concept|Hospital Course|14267,14277|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|14267,14277|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Finding|Hospital Course|14278,14284|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|14278,14284|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|14285,14294|false|false|false|||affecting
Event|Event|Hospital Course|14295,14305|false|false|false|||motivation
Finding|Mental Process|Hospital Course|14295,14305|false|true|false|C0026605|Motivation|motivation
Attribute|Clinical Attribute|Hospital Course|14314,14323|false|false|false|C0945731||diagnosis
Event|Event|Hospital Course|14314,14323|false|false|false|||diagnosis
Finding|Classification|Hospital Course|14314,14323|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|14314,14323|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14314,14323|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|Hospital Course|14329,14338|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|14329,14338|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|14329,14338|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|14329,14338|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|14329,14338|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Neoplastic Process|Hospital Course|14348,14358|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|14348,14358|false|false|false|||malignancy
Event|Event|Hospital Course|14364,14370|true|false|false|||denied
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14378,14386|true|false|false|C0438696|Suicidal|suicidal
Event|Event|Hospital Course|14378,14386|true|false|false|||suicidal
Event|Event|Hospital Course|14388,14396|true|false|false|||ideation
Finding|Mental Process|Hospital Course|14388,14396|true|false|false|C0392348|ideation|ideation
Event|Event|Hospital Course|14412,14420|true|false|false|||declined
Finding|Idea or Concept|Hospital Course|14421,14425|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|14421,14425|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|14421,14425|true|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|14426,14436|true|false|false|C0074393|sertraline|sertraline
Drug|Pharmacologic Substance|Hospital Course|14426,14436|true|false|false|C0074393|sertraline|sertraline
Event|Event|Hospital Course|14426,14436|true|false|false|||sertraline
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14461,14466|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|14461,14466|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|14461,14466|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|14461,14466|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|14461,14466|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|14461,14466|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|14461,14466|false|false|false|||liver
Finding|Finding|Hospital Course|14461,14466|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|14461,14466|false|false|false|C0872387|Procedures on liver|liver
Procedure|Diagnostic Procedure|Hospital Course|14461,14473|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Procedure|Health Care Activity|Hospital Course|14461,14473|false|false|false|C0193388;C1548877|Biopsy of liver (procedure);Consent Type - Liver Biopsy|liver biopsy
Event|Event|Hospital Course|14467,14473|false|false|false|||biopsy
Finding|Finding|Hospital Course|14467,14473|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|14467,14473|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|14467,14473|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|14467,14473|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|14475,14484|false|false|false|||believing
Event|Event|Hospital Course|14497,14505|false|false|false|||supposed
Event|Event|Hospital Course|14512,14516|false|false|false|||held
Event|Event|Hospital Course|14542,14553|false|false|false|||explanation
Finding|Intellectual Product|Hospital Course|14542,14553|false|false|false|C0681841|Explanation|explanation
Event|Event|Hospital Course|14580,14584|false|false|false|||seen
Finding|Functional Concept|Hospital Course|14588,14594|false|false|false|C0728831|Social|social
Event|Event|Hospital Course|14595,14599|false|false|false|||work
Event|Occupational Activity|Hospital Course|14595,14599|false|false|false|C0043227|Work|work
Event|Event|Hospital Course|14611,14620|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|14611,14620|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|14639,14645|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|14639,14645|false|false|false|||anemia
Attribute|Clinical Attribute|Hospital Course|14647,14657|false|false|false|C1542366|hematocrit attribute|Hematocrit
Event|Event|Hospital Course|14647,14657|false|false|false|||Hematocrit
Finding|Finding|Hospital Course|14647,14657|false|false|false|C0518014|Hematocrit level|Hematocrit
Procedure|Laboratory Procedure|Hospital Course|14647,14657|false|false|false|C0018935|Hematocrit Measurement|Hematocrit
Event|Event|Hospital Course|14667,14673|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|14667,14673|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|14679,14689|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|14679,14689|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|14679,14694|false|false|false|C0332290|Consistent with|consistent with
Drug|Biomedical or Dental Material|Hospital Course|14702,14710|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|14702,14710|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|14702,14710|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|14735,14744|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|14735,14744|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|14763,14769|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|14763,14769|false|false|false|||anemia
Disorder|Disease or Syndrome|Hospital Course|14763,14788|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic disease
Finding|Intellectual Product|Hospital Course|14773,14780|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|14773,14780|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|14773,14788|false|false|false|C0008679|Chronic disease|chronic disease
Disorder|Disease or Syndrome|Hospital Course|14781,14788|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|14781,14788|false|false|false|||disease
Drug|Pharmacologic Substance|Hospital Course|14797,14802|false|false|false|C1874451|Basis|basis
Event|Event|Hospital Course|14797,14802|false|false|false|||basis
Finding|Functional Concept|Hospital Course|14797,14802|false|false|false|C1527178|Basis - conceptual entity|basis
Event|Event|Hospital Course|14819,14823|false|false|false|||labs
Lab|Laboratory or Test Result|Hospital Course|14819,14823|false|false|false|C0587081|Laboratory test finding|labs
Drug|Food|Hospital Course|14825,14830|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|Hospital Course|14825,14836|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|Hospital Course|14825,14836|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|Hospital Course|14831,14836|false|false|false|||signs
Finding|Finding|Hospital Course|14831,14836|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|14831,14836|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|14846,14852|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|14846,14852|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|14864,14873|true|false|false|||exception
Finding|Conceptual Entity|Hospital Course|14864,14873|true|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Idea or Concept|Hospital Course|14864,14873|true|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Event|Event|Hospital Course|14888,14899|true|false|false|||tachycardia
Finding|Finding|Hospital Course|14888,14899|true|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Hospital Course|14909,14914|true|false|false|||signs
Finding|Finding|Hospital Course|14909,14914|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|14909,14914|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|14926,14934|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|14926,14934|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Functional Concept|Hospital Course|14946,14954|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Finding|Idea or Concept|Hospital Course|14946,14954|false|false|false|C0205409;C1548221|Bed Status - Isolated;Isolated|isolated
Disorder|Disease or Syndrome|Hospital Course|14955,14960|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|14955,14960|false|false|false|||blood
Finding|Body Substance|Hospital Course|14955,14960|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Hospital Course|14970,14976|false|false|false|||emesis
Finding|Body Substance|Hospital Course|14970,14976|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|14970,14976|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|14970,14976|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Idea or Concept|Hospital Course|14980,14985|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|Hospital Course|14993,15005|false|false|false|C0005779|Blood Coagulation Disorders|Coagulopathy
Event|Event|Hospital Course|14993,15005|false|false|false|||Coagulopathy
Attribute|Clinical Attribute|Hospital Course|15007,15010|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|Hospital Course|15007,15010|false|false|false|||INR
Procedure|Laboratory Procedure|Hospital Course|15007,15010|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15007,15010|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|Hospital Course|15029,15033|false|false|false|||felt
Event|Event|Hospital Course|15037,15044|false|false|false|||reflect
Finding|Mental Process|Hospital Course|15037,15044|false|false|false|C0558058|Reflecting|reflect
Event|Activity|Hospital Course|15046,15055|false|false|false|C1883254|Synthesis|synthetic
Disorder|Disease or Syndrome|Hospital Course|15056,15067|false|true|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|15056,15067|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|15056,15067|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|15056,15067|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|15056,15067|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Mental Process|Hospital Course|15075,15082|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Location or Region|Hospital Course|15086,15093|false|false|false|C0205054|Hepatic|hepatic
Event|Event|Hospital Course|15094,15106|false|false|false|||infiltration
Finding|Functional Concept|Hospital Course|15094,15106|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|Hospital Course|15094,15106|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15094,15106|false|false|false|C0702249|Infiltration (procedure)|infiltration
Disorder|Neoplastic Process|Hospital Course|15111,15121|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|15111,15121|false|false|false|||malignancy
Finding|Finding|Hospital Course|15126,15130|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|Hospital Course|15134,15138|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Anatomy|Body Space or Junction|Hospital Course|15139,15143|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|15139,15143|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|15139,15143|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|15139,15143|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Finding|Hospital Course|15139,15150|false|false|false|C2137071|Oral intake|oral intake
Event|Event|Hospital Course|15144,15150|false|false|false|||intake
Finding|Functional Concept|Hospital Course|15144,15150|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|15144,15150|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|Hospital Course|15166,15171|true|false|false|||signs
Finding|Finding|Hospital Course|15166,15171|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|15166,15171|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|15183,15191|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|15183,15191|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|15202,15211|false|false|false|||exception
Finding|Conceptual Entity|Hospital Course|15202,15211|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Idea or Concept|Hospital Course|15202,15211|false|false|false|C1554961;C1705847|Exception - Property or Attribute;exception - ResponseLevel|exception
Finding|Finding|Hospital Course|15215,15224|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Event|Event|Hospital Course|15225,15236|false|false|false|||hematemesis
Finding|Sign or Symptom|Hospital Course|15225,15236|false|false|false|C0018926|Hematemesis|hematemesis
Finding|Idea or Concept|Hospital Course|15241,15246|false|false|false|C1552828|Table Frame - above|above
Finding|Idea or Concept|Hospital Course|15249,15261|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Body Substance|Hospital Course|15271,15278|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|15271,15278|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|15271,15278|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Health Care Activity|Hospital Course|15271,15288|false|false|false|C0030685|Patient Discharge|Patient discharge
Event|Event|Hospital Course|15279,15288|false|false|false|||discharge
Finding|Body Substance|Hospital Course|15279,15288|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|15279,15288|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|15279,15288|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|15279,15288|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15279,15293|false|false|false|C0184713|Discharge to home|discharge home
Event|Event|Hospital Course|15289,15293|false|false|false|||home
Finding|Idea or Concept|Hospital Course|15289,15293|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|15289,15293|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|15289,15293|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|15299,15303|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|15299,15303|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|15299,15303|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|Hospital Course|15299,15311|false|false|false|C3275086|Home Hospice|home hospice
Event|Event|Hospital Course|15304,15311|false|false|false|||hospice
Procedure|Health Care Activity|Hospital Course|15304,15311|false|false|false|C0085555|Hospice Care|hospice
Attribute|Clinical Attribute|Hospital Course|15314,15325|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|15314,15325|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|15314,15325|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|15314,15325|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|15314,15338|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|15329,15338|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|15329,15338|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|15357,15367|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|15357,15367|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|15357,15372|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|15368,15372|false|false|false|||list
Finding|Intellectual Product|Hospital Course|15368,15372|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|15380,15390|false|false|false|||inaccurate
Event|Event|Hospital Course|15395,15403|false|false|false|||requires
Event|Event|Hospital Course|15412,15425|false|false|false|||investigation
Finding|Intellectual Product|Hospital Course|15412,15425|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Hospital Course|15412,15425|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Hospital Course|15430,15439|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|15430,15439|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|15440,15447|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|15464,15467|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|15468,15471|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|15468,15471|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Hospital Course|15476,15485|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|Hospital Course|15476,15485|false|false|false|C0085208|bupropion|BuPROPion
Drug|Organic Chemical|Hospital Course|15506,15516|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|15506,15516|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|Hospital Course|15534,15544|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|15534,15544|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|15565,15574|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|Hospital Course|15565,15574|false|false|false|C0040805|trazodone|traZODONE
Finding|Gene or Genome|Hospital Course|15588,15591|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|15592,15597|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|15592,15597|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|15592,15597|false|false|false|||sleep
Finding|Organism Function|Hospital Course|15592,15597|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|15602,15613|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|Hospital Course|15602,15613|false|false|false|C0061851|ondansetron|Ondansetron
Finding|Gene or Genome|Hospital Course|15626,15629|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|15630,15636|false|false|false|C4255480||nausea
Event|Event|Hospital Course|15630,15636|false|false|false|||nausea
Finding|Sign or Symptom|Hospital Course|15630,15636|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|Hospital Course|15641,15650|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|15641,15650|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|Hospital Course|15669,15672|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|15673,15685|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|15673,15685|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|15690,15699|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|15690,15699|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|15690,15699|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|15690,15699|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|15701,15710|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|15701,15710|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|15701,15718|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|15711,15718|false|false|false|||Release
Finding|Functional Concept|Hospital Course|15711,15718|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|15711,15718|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15711,15718|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|15733,15736|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|15737,15741|false|false|false|C2598155||pain
Event|Event|Hospital Course|15737,15741|false|false|false|||pain
Finding|Functional Concept|Hospital Course|15737,15741|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|15737,15741|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|15750,15754|false|false|false|||hold
Event|Event|Hospital Course|15759,15767|false|false|false|||sedation
Finding|Finding|Hospital Course|15759,15767|false|false|false|C0235195;C5400562|Sedated state;Sedation|sedation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15759,15767|false|false|false|C0344106|Sedation procedure|sedation
Drug|Organic Chemical|Hospital Course|15779,15789|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|15779,15789|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|15779,15789|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|15779,15796|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|15779,15796|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|15790,15796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|15790,15796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|15790,15796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|15790,15796|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|15790,15796|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|15790,15796|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|15816,15825|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|15816,15825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|15816,15825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|15816,15825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|15816,15825|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|15816,15837|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|15826,15837|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|15826,15837|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|15826,15837|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|15826,15837|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|15842,15851|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|Hospital Course|15842,15851|false|false|false|C0085208|bupropion|BuPROPion
Drug|Organic Chemical|Hospital Course|15872,15883|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|Hospital Course|15872,15883|false|false|false|C0061851|ondansetron|Ondansetron
Finding|Gene or Genome|Hospital Course|15896,15899|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|15900,15906|false|false|false|C4255480||nausea
Event|Event|Hospital Course|15900,15906|false|false|false|||nausea
Finding|Sign or Symptom|Hospital Course|15900,15906|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|Hospital Course|15911,15919|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|Hospital Course|15911,15919|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|Hospital Course|15911,15919|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|Hospital Course|15911,15919|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|Hospital Course|15921,15927|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|Hospital Course|15921,15927|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|Hospital Course|15942,15945|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|15946,15950|false|false|false|C2598155||pain
Event|Event|Hospital Course|15946,15950|false|false|false|||pain
Finding|Functional Concept|Hospital Course|15946,15950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|15946,15950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|15956,15964|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|15956,15964|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|15956,15964|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|15956,15964|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|15973,15979|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|15983,15991|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|15986,15991|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|15986,15991|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|16024,16030|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|16031,16038|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|16031,16038|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|16045,16050|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|16045,16050|false|false|false|C3489575|sennosides, USP|Senna
Drug|Biomedical or Dental Material|Hospital Course|16053,16056|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|16053,16056|false|false|false|||TAB
Disorder|Mental or Behavioral Dysfunction|Hospital Course|16060,16063|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|16060,16063|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|16060,16063|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|16060,16063|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|16060,16063|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|16064,16067|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|16068,16080|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|16068,16080|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|16086,16096|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|Hospital Course|16086,16096|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Biomedical or Dental Material|Hospital Course|16112,16118|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|16112,16118|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|16119,16127|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|16122,16127|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|16122,16127|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|16137,16140|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|16137,16140|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|16151,16157|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|16158,16165|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|16158,16165|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|16172,16182|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|16172,16182|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|16203,16213|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|16203,16213|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|16203,16213|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|16222,16229|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|16222,16229|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|16222,16229|false|false|false|C0006935|capsule (pharmacologic)|capsule
Event|Event|Hospital Course|16230,16237|false|false|false|||delayed
Anatomy|Body Location or Region|Hospital Course|16246,16251|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|16246,16251|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|16268,16275|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|16268,16275|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|16268,16275|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|16276,16283|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|16276,16283|false|false|false|C0807726|refill|Refills
Finding|Idea or Concept|Hospital Course|16290,16298|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Disorder|Disease or Syndrome|Hospital Course|16299,16302|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|Hospital Course|16299,16302|false|false|false|||Bed
Finding|Intellectual Product|Hospital Course|16299,16302|false|false|false|C2346952|Bachelor of Education|Bed
Finding|Idea or Concept|Hospital Course|16313,16321|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Disorder|Disease or Syndrome|Hospital Course|16322,16325|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|Hospital Course|16322,16325|false|false|false|||Bed
Finding|Intellectual Product|Hospital Course|16322,16325|false|false|false|C2346952|Bachelor of Education|Bed
Drug|Organic Chemical|Hospital Course|16330,16341|false|false|false|C0723712|Therapeutic brand of coal tar|Therapeutic
Drug|Pharmacologic Substance|Hospital Course|16330,16341|false|false|false|C0723712|Therapeutic brand of coal tar|Therapeutic
Event|Event|Hospital Course|16330,16341|false|false|false|||Therapeutic
Finding|Functional Concept|Hospital Course|16330,16341|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|Therapeutic
Finding|Intellectual Product|Hospital Course|16330,16341|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|Therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|16330,16341|false|false|false|C0087111|Therapeutic procedure|Therapeutic
Procedure|Health Care Activity|Hospital Course|16367,16374|false|false|false|C0085555|Hospice Care|Hospice
Event|Activity|Hospital Course|16375,16380|false|false|false|C1705178|Order (action)|Order
Event|Event|Hospital Course|16375,16380|false|false|false|||Order
Finding|Classification|Hospital Course|16375,16380|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|Order
Finding|Idea or Concept|Hospital Course|16375,16380|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|Order
Finding|Intellectual Product|Hospital Course|16375,16380|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|Order
Phenomenon|Natural Phenomenon or Process|Hospital Course|16375,16380|false|false|false|C1373200|Order [PK]|Order
Event|Event|Hospital Course|16388,16394|false|false|false|||Screen
Event|Event|Hospital Course|16399,16404|false|false|false|||Admit
Event|Event|Hospital Course|16408,16415|false|false|false|||Hospice
Procedure|Health Care Activity|Hospital Course|16408,16415|false|false|false|C0085555|Hospice Care|Hospice
Drug|Organic Chemical|Hospital Course|16420,16429|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|16420,16429|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|Hospital Course|16448,16451|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|16452,16464|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|16452,16464|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|16469,16477|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|16469,16477|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|16469,16477|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|16469,16484|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|16469,16484|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|16478,16484|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|16478,16484|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|16478,16484|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|16478,16484|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|16478,16484|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|16478,16484|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|16495,16498|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|16495,16498|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|16495,16498|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|16495,16498|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|16495,16498|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|16504,16514|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|16504,16514|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|16536,16545|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|Hospital Course|16536,16545|false|false|false|C0040805|trazodone|traZODONE
Finding|Gene or Genome|Hospital Course|16559,16562|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|16563,16568|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|16563,16568|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|16563,16568|false|false|false|||sleep
Finding|Organism Function|Hospital Course|16563,16568|false|false|false|C0037313|Sleep|sleep
Drug|Biomedical or Dental Material|Hospital Course|16574,16586|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|16574,16586|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|16574,16586|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|16574,16593|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|16574,16593|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|16587,16593|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|16587,16593|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|16587,16593|false|false|false|||Glycol
Finding|Gene or Genome|Hospital Course|16608,16611|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|16612,16624|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|16612,16624|false|false|false|C0009806|Constipation|constipation
Event|Event|Hospital Course|16629,16638|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|16629,16638|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|16629,16638|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|16629,16638|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|16629,16638|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|16629,16650|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|16629,16650|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|16639,16650|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|16639,16650|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|16639,16650|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|16652,16656|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|16652,16656|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|16652,16656|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|16652,16656|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|16662,16669|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|16662,16669|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|16672,16680|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|16672,16680|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|16688,16697|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|16688,16697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|16688,16697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|16688,16697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|16688,16697|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|16688,16707|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|16698,16707|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|16698,16707|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|16698,16707|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|16698,16707|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|16698,16707|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|16718,16728|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|Hospital Course|16718,16749|false|false|false|C4324497|Adenocarcinoma of colon metastatic|Metastatic colon adenocarcinoma
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|16729,16734|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Hospital Course|16729,16734|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Hospital Course|16729,16734|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Hospital Course|16729,16734|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Hospital Course|16729,16749|false|false|false|C0338106|Adenocarcinoma of colon|colon adenocarcinoma
Disorder|Neoplastic Process|Hospital Course|16735,16749|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|16735,16749|false|false|false|||adenocarcinoma
Finding|Mental Process|Discharge Condition|16774,16780|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|16774,16787|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|16774,16787|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|16781,16787|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|16781,16787|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|16789,16797|false|false|false|C0009676|Confusion|Confused
Event|Event|Discharge Condition|16789,16797|false|false|false|||Confused
Finding|Finding|Discharge Condition|16789,16797|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|16789,16797|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Event|Discharge Condition|16811,16816|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|16811,16833|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|16811,16833|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|16820,16833|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|16820,16833|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|16820,16833|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|16835,16840|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|16835,16840|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|16835,16840|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|16835,16840|false|false|false|||Alert
Finding|Finding|Discharge Condition|16835,16840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|16835,16840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|16835,16840|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|16845,16856|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|16845,16856|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|16858,16866|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|16858,16866|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|16858,16866|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|16867,16873|false|false|false|C5889824||Status
Event|Event|Discharge Condition|16867,16873|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|16867,16873|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|16875,16883|false|false|false|||Bedbound
Finding|Finding|Discharge Condition|16875,16883|false|false|false|C0425251|Bed-ridden|Bedbound
Finding|Gene or Genome|Discharge Instructions|16912,16916|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|16935,16943|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|16935,16943|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|16935,16943|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|Discharge Instructions|16951,16955|false|false|false|||part
Finding|Idea or Concept|Discharge Instructions|16951,16955|false|false|false|C1552020|Role Class - part|part
Event|Activity|Discharge Instructions|16964,16968|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|16964,16968|false|false|false|||care
Finding|Finding|Discharge Instructions|16964,16968|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|16964,16968|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|16981,16990|false|false|false|||admission
Procedure|Health Care Activity|Discharge Instructions|16981,16990|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Discharge Instructions|17023,17031|false|false|false|||admitted
Event|Event|Discharge Instructions|17036,17045|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|17036,17055|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|17036,17055|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|17049,17055|false|false|false|C0225386|Breath|breath
Finding|Finding|Discharge Instructions|17057,17063|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|17057,17063|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Discharge Instructions|17076,17086|true|false|false|||underlying
Finding|Finding|Discharge Instructions|17076,17086|true|false|false|C4722602|Underlying|underlying
Disorder|Neoplastic Process|Discharge Instructions|17088,17094|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Discharge Instructions|17088,17094|true|false|false|||cancer
Event|Event|Discharge Instructions|17113,17121|true|false|false|||evidence
Finding|Idea or Concept|Discharge Instructions|17113,17121|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|17113,17124|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Discharge Instructions|17125,17134|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|17125,17134|true|false|false|||pneumonia
Disorder|Disease or Syndrome|Discharge Instructions|17138,17143|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|17138,17143|true|false|false|||blood
Finding|Body Substance|Discharge Instructions|17138,17143|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|Discharge Instructions|17138,17148|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|Discharge Instructions|17144,17148|true|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|17144,17148|true|false|false|C0009074|clotrimazole|clot
Event|Event|Discharge Instructions|17144,17148|true|false|false|||clot
Finding|Pathologic Function|Discharge Instructions|17144,17148|true|false|false|C0302148|Blood Clot|clot
Disorder|Disease or Syndrome|Discharge Instructions|17157,17162|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|17157,17162|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|17157,17162|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17157,17170|false|false|false|C0005847|Blood Vessel|blood vessels
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17163,17170|false|false|false|C0005847|Blood Vessel|vessels
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17179,17184|false|false|false|C0024109|Lung|lungs
Event|Event|Discharge Instructions|17191,17200|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|17191,17210|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|17191,17210|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|17204,17210|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|17212,17220|false|false|false|||resolved
Event|Event|Discharge Instructions|17235,17240|false|false|false|||found
Event|Event|Discharge Instructions|17249,17257|false|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|17249,17257|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Functional Concept|Discharge Instructions|17266,17270|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17266,17276|false|false|false|C0230426|Structure of left thigh|left thigh
Anatomy|Body Location or Region|Discharge Instructions|17271,17276|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Anatomy|Body Location or Region|Discharge Instructions|17282,17291|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|17282,17296|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Discharge Instructions|17292,17296|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|17292,17296|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|17292,17296|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|17292,17296|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|17311,17318|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Discharge Instructions|17311,17318|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Procedure|Diagnostic Procedure|Discharge Instructions|17311,17326|true|false|false|C1881134|imaging studies|imaging studies
Event|Event|Discharge Instructions|17319,17326|true|false|false|||studies
Procedure|Research Activity|Discharge Instructions|17319,17326|true|false|false|C0947630|Scientific Study|studies
Event|Event|Discharge Instructions|17340,17353|true|false|false|||investigation
Finding|Intellectual Product|Discharge Instructions|17340,17353|true|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Discharge Instructions|17340,17353|true|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Attribute|Clinical Attribute|Discharge Instructions|17363,17371|false|false|false|C2926606||findings
Event|Event|Discharge Instructions|17363,17371|false|false|false|||findings
Finding|Functional Concept|Discharge Instructions|17363,17371|false|false|false|C2607943|findings aspects|findings
Event|Event|Discharge Instructions|17387,17393|false|false|false|||biopsy
Finding|Finding|Discharge Instructions|17387,17393|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Discharge Instructions|17387,17393|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Discharge Instructions|17387,17393|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Discharge Instructions|17387,17393|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17403,17408|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|17403,17408|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|17403,17408|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|17403,17408|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|17403,17408|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|17403,17408|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Discharge Instructions|17403,17408|false|false|false|||liver
Finding|Finding|Discharge Instructions|17403,17408|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|17403,17408|false|false|false|C0872387|Procedures on liver|liver
Event|Event|Discharge Instructions|17414,17422|false|false|false|||revealed
Disorder|Neoplastic Process|Discharge Instructions|17432,17438|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Discharge Instructions|17432,17438|false|false|false|||cancer
Event|Event|Discharge Instructions|17439,17444|false|false|false|||known
Event|Event|Discharge Instructions|17448,17454|false|false|false|||affect
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17460,17465|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|17460,17465|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|17460,17465|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|17460,17465|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|17460,17465|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|17460,17465|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Discharge Instructions|17460,17465|false|false|false|||liver
Finding|Finding|Discharge Instructions|17460,17465|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|17460,17465|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17471,17476|false|false|false|C0024109|Lung|lungs
Event|Event|Discharge Instructions|17477,17487|false|false|false|||originated
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17496,17501|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Discharge Instructions|17496,17501|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Discharge Instructions|17496,17501|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Discharge Instructions|17496,17501|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Gene or Genome|Discharge Instructions|17503,17508|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17503,17514|false|false|false|C0021851|Large Intestine|large bowel
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|17509,17514|false|false|false|C0021853|Intestines|bowel
Event|Event|Discharge Instructions|17527,17538|false|false|false|||transferred
Disorder|Neoplastic Process|Discharge Instructions|17546,17554|false|false|false|C0027651|Neoplasms|oncology
Event|Event|Discharge Instructions|17546,17554|false|false|false|||oncology
Procedure|Health Care Activity|Discharge Instructions|17546,17554|false|false|false|C1555459|oncology services|oncology
Procedure|Health Care Activity|Discharge Instructions|17546,17562|false|false|false|C1555459|oncology services|oncology service
Event|Occupational Activity|Discharge Instructions|17555,17562|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Discharge Instructions|17555,17562|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Discharge Instructions|17583,17595|false|false|false|||chemotherapy
Finding|Functional Concept|Discharge Instructions|17583,17595|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17583,17595|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Discharge Instructions|17610,17614|false|false|false|||harm
Event|Event|Discharge Instructions|17628,17632|false|false|false|||good
Finding|Idea or Concept|Discharge Instructions|17628,17632|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|Discharge Instructions|17649,17659|false|false|false|||discussion
Finding|Social Behavior|Discharge Instructions|17649,17659|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17649,17659|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Idea or Concept|Discharge Instructions|17678,17684|false|false|false|C0018684|Health|health
Procedure|Health Care Activity|Discharge Instructions|17678,17689|false|false|false|C0086388|Health Care|health care
Event|Activity|Discharge Instructions|17685,17689|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|17685,17689|false|false|false|||care
Finding|Finding|Discharge Instructions|17685,17689|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|17685,17689|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|17690,17695|false|false|false|C3897813|Advance Directive - Proxy|proxy
Event|Event|Discharge Instructions|17704,17711|false|false|false|||decided
Event|Event|Discharge Instructions|17730,17734|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|17730,17734|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|17730,17734|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|17730,17734|false|false|false|C1553498|home health encounter|home
Finding|Classification|Discharge Instructions|17751,17757|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|17751,17757|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|17751,17757|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|17751,17757|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Mental Process|Discharge Instructions|17762,17767|false|false|false|C0024028|Love|loved
Event|Event|Discharge Instructions|17789,17792|false|false|false|||set
Procedure|Health Care Activity|Discharge Instructions|17796,17803|false|false|false|C0085555|Hospice Care|hospice
Event|Occupational Activity|Discharge Instructions|17796,17812|false|false|false|C5423046|Purchased Services, Clinical and Biomedical, Home Healthcare, Hospice|hospice services
Event|Event|Discharge Instructions|17804,17812|false|false|false|||services
Event|Occupational Activity|Discharge Instructions|17804,17812|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Discharge Instructions|17804,17812|false|false|false|C1704289|Clinical Service|services
Event|Event|Discharge Instructions|17838,17842|true|false|false|||help
Event|Event|Discharge Instructions|17853,17859|true|false|false|||issues
Event|Event|Discharge Instructions|17865,17870|true|false|false|||arise
Finding|Finding|Discharge Instructions|17885,17892|false|false|false|C4534363|At home|at home
Event|Event|Discharge Instructions|17888,17892|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|17888,17892|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|17888,17892|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|17888,17892|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|Discharge Instructions|17898,17906|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|17907,17919|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|17907,17919|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|17907,17919|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

