 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|40,49|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|40,54|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|74,83|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|74,88|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|130,133|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|141,148|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|141,148|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|150,158|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Finding|Body Substance|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|Allergies|209,218|true|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|209,218|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|222,227|false|false|false|C0013227|Pharmaceutical Preparations|Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|222,227|false|false|false|C3687832|Drugs - dental services|Drugs
Finding|Functional Concept|Allergies|230,239|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|265,274|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|Chief Complaint|265,285|false|false|false|C0000731|Abdomen distended|Abdominal distention
Finding|Finding|Chief Complaint|275,285|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Chief Complaint|275,285|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|Chief Complaint|286,290|false|false|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|286,290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|286,290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Chief Complaint|286,300|false|false|false|C3499958|Pain and Fever|pain and fever
Drug|Pharmacologic Substance|Chief Complaint|286,300|false|false|false|C3499958|Pain and Fever|pain and fever
Finding|Finding|Chief Complaint|295,300|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Chief Complaint|295,300|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Classification|Chief Complaint|303,308|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|309,317|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|309,317|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|321,339|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|330,339|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|330,339|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|330,339|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|330,339|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|341,353|false|false|false|C0034115|Paracentesis|Paracentesis
Drug|Indicator, Reagent, or Diagnostic Aid|Chief Complaint|359,369|false|false|false|C0358514|Diagnostic agents|diagnostic
Finding|Functional Concept|Chief Complaint|359,369|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|Chief Complaint|359,369|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|Chief Complaint|359,369|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Drug|Organic Chemical|Chief Complaint|380,391|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Chief Complaint|380,391|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Finding|Functional Concept|Chief Complaint|380,391|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Chief Complaint|380,391|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|380,391|false|false|false|C0087111|Therapeutic procedure|therapeutic
Disorder|Disease or Syndrome|History of Present Illness|452,471|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|History of Present Illness|462,471|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Disorder|Disease or Syndrome|History of Present Illness|485,492|false|false|false|C0003962|Ascites|ascites
Finding|Pathologic Function|History of Present Illness|485,492|false|false|false|C5441966|Peritoneal Effusion|ascites
Finding|Sign or Symptom|History of Present Illness|509,515|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|History of Present Illness|520,532|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|History of Present Illness|520,532|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Disorder|Disease or Syndrome|History of Present Illness|567,576|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Finding|Idea or Concept|History of Present Illness|610,619|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|History of Present Illness|620,629|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|620,640|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|History of Present Illness|630,640|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|630,640|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|History of Present Illness|642,646|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Pathologic Function|History of Present Illness|652,668|false|false|false|C0476474|Persistent fever|persistent fever
Finding|Finding|History of Present Illness|663,668|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|663,668|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|682,688|true|false|false|C0085593|Chills|chills
Finding|Intellectual Product|History of Present Illness|697,708|false|false|false|C4084908|Have Sweats|have sweats
Finding|Body Substance|History of Present Illness|702,708|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|702,708|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Procedure|Health Care Activity|History of Present Illness|728,737|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Individual Behavior|History of Present Illness|769,778|false|false|false|C1321605|Compliance behavior|compliant
Finding|Finding|History of Present Illness|788,791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|788,791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Food|History of Present Illness|799,803|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|History of Present Illness|799,803|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|799,803|false|false|false|C0012159|Diet therapy|diet
Drug|Substance|History of Present Illness|809,814|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|809,814|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|809,826|false|false|false|C0204700|Fluid restriction|fluid restriction
Finding|Functional Concept|History of Present Illness|815,826|false|false|false|C0443288|Restricted|restriction
Finding|Finding|History of Present Illness|843,852|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|History of Present Illness|843,852|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Drug|Substance|History of Present Illness|853,858|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|853,858|true|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Biologically Active Substance|History of Present Illness|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|History of Present Illness|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|History of Present Illness|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|History of Present Illness|862,868|true|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|History of Present Illness|862,868|true|false|false|C0337443|Sodium measurement|sodium
Finding|Functional Concept|History of Present Illness|870,876|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|History of Present Illness|870,876|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Individual Behavior|History of Present Illness|890,898|false|false|false|C0680686|sobriety|sobriety
Drug|Organic Chemical|History of Present Illness|904,911|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|History of Present Illness|904,911|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|History of Present Illness|904,911|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Sign or Symptom|History of Present Illness|939,946|false|false|false|C0015967|Fever|febrile
Procedure|Diagnostic Procedure|History of Present Illness|961,970|false|false|false|C0030247|Palpation|palpation
Finding|Idea or Concept|History of Present Illness|1020,1027|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1028,1033|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1028,1039|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1028,1039|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|History of Present Illness|1034,1039|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1034,1039|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Gene or Genome|History of Present Illness|1080,1084|false|false|false|C1823816|C1orf210 gene|temp
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1080,1084|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|temp
Attribute|Clinical Attribute|History of Present Illness|1112,1117|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|History of Present Illness|1112,1117|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|History of Present Illness|1112,1117|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|History of Present Illness|1112,1117|false|false|false|C0034107|Pulse taking|pulse
Drug|Organic Chemical|History of Present Illness|1146,1152|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|History of Present Illness|1146,1152|false|false|false|C0699194|Ativan|Ativan
Drug|Organic Chemical|History of Present Illness|1167,1175|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|History of Present Illness|1167,1175|false|false|false|C0026549|morphine|morphine
Attribute|Clinical Attribute|History of Present Illness|1191,1195|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1191,1195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1191,1195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|1197,1204|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|History of Present Illness|1197,1204|false|false|false|C0699142|Tylenol|tylenol
Finding|Finding|History of Present Illness|1220,1225|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1220,1225|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|History of Present Illness|1227,1238|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|History of Present Illness|1227,1238|false|false|false|C0061851|ondansetron|ondansetron
Attribute|Clinical Attribute|History of Present Illness|1253,1259|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|1253,1259|false|false|false|C0027497|Nausea|nausea
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1292,1299|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|History of Present Illness|1292,1299|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|1317,1327|false|false|false|C0358514|Diagnostic agents|diagnostic
Finding|Functional Concept|History of Present Illness|1317,1327|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|History of Present Illness|1317,1327|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|History of Present Illness|1317,1327|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1329,1341|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Antibiotic|History of Present Illness|1401,1412|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|History of Present Illness|1401,1412|false|false|false|C0007561|ceftriaxone|ceftriaxone
Finding|Finding|History of Present Illness|1426,1434|false|false|false|C0332149|Possible|possible
Attribute|Clinical Attribute|History of Present Illness|1435,1438|false|true|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1435,1438|false|true|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|1435,1438|false|true|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|History of Present Illness|1435,1438|false|true|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|1435,1438|false|true|false|C1306620|Systolic blood pressure measurement|SBP
Drug|Pharmacologic Substance|History of Present Illness|1461,1469|false|false|false|C0013227|Pharmaceutical Preparations|Medicine
Event|Occupational Activity|History of Present Illness|1482,1492|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|1482,1492|false|false|false|C0376636|Disease Management|management
Anatomy|Anatomical Structure|History of Present Illness|1556,1561|false|false|false|C3714591|Floor (anatomic)|floor
Anatomy|Anatomical Structure|History of Present Illness|1576,1581|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|History of Present Illness|1586,1590|false|false|false|C2713234||mood
Finding|Conceptual Entity|History of Present Illness|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|History of Present Illness|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|History of Present Illness|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Disorder|Disease or Syndrome|History of Present Illness|1612,1617|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Finding|History of Present Illness|1618,1625|false|false|false|C0424109|Weepiness|tearful
Disorder|Disease or Syndrome|History of Present Illness|1634,1639|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Mental Process|History of Present Illness|1640,1648|false|false|false|C2987187|Pleasant|pleasant
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1690,1698|true|false|false|C0009676|Confusion|confused
Finding|Finding|History of Present Illness|1690,1698|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Finding|Intellectual Product|History of Present Illness|1690,1698|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Drug|Organic Chemical|History of Present Illness|1741,1746|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1741,1746|true|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|1741,1746|true|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|History of Present Illness|1748,1755|true|false|false|C0013428|Dysuria|dysuria
Finding|Finding|History of Present Illness|1758,1766|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1758,1766|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|History of Present Illness|1771,1775|false|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|History of Present Illness|1771,1775|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|1771,1775|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Finding|History of Present Illness|1794,1803|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Finding|Idea or Concept|History of Present Illness|1836,1842|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|1836,1842|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|1836,1845|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|1836,1853|false|false|false|C0488564;C0488565||Review of Systems
Procedure|Health Care Activity|History of Present Illness|1836,1853|false|false|false|C0489633|Review of systems (procedure)|Review of Systems
Finding|Functional Concept|History of Present Illness|1846,1853|false|false|false|C0449913|System|Systems
Disorder|Disease or Syndrome|History of Present Illness|1865,1868|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Finding|Finding|History of Present Illness|1865,1868|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|1865,1868|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Sign or Symptom|History of Present Illness|1882,1888|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|1897,1905|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|History of Present Illness|1907,1912|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|1907,1912|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|1907,1912|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|1907,1912|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Mental Process|History of Present Illness|1913,1923|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|1913,1923|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|1925,1935|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Finding|Pathologic Function|History of Present Illness|1940,1950|false|false|false|C0700148|Congestion|congestion
Anatomy|Body Location or Region|History of Present Illness|1959,1964|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1959,1964|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1959,1969|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1959,1969|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1965,1969|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1965,1969|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1965,1969|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|1984,1996|false|false|false|C0030252|Palpitations|palpitations
Drug|Organic Chemical|History of Present Illness|2006,2011|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|2006,2011|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|2006,2011|false|false|false|C0010200|Coughing|cough
Attribute|Clinical Attribute|History of Present Illness|2013,2032|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|2013,2032|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|2026,2032|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|History of Present Illness|2037,2044|true|false|false|C0043144|Wheezing|wheezes
Attribute|Clinical Attribute|History of Present Illness|2053,2059|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|2053,2059|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|2062,2070|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|History of Present Illness|2072,2080|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2072,2080|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2082,2094|false|false|false|C0009806|Constipation|constipation
Finding|Functional Concept|History of Present Illness|2106,2112|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2106,2112|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|History of Present Illness|2106,2115|true|false|false|C0392747|Changing|change in
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2116,2121|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2126,2133|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|2126,2133|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2126,2133|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Finding|History of Present Illness|2134,2140|false|false|false|C0018464;C2242848|Behaviorial Habits;habits (history)|habits
Finding|Individual Behavior|History of Present Illness|2134,2140|false|false|false|C0018464;C2242848|Behaviorial Habits;habits (history)|habits
Finding|Sign or Symptom|History of Present Illness|2145,2152|true|false|false|C0013428|Dysuria|dysuria
Finding|Sign or Symptom|History of Present Illness|2161,2172|true|false|false|C0003862|Arthralgia|arthralgias
Finding|Sign or Symptom|History of Present Illness|2176,2184|true|false|false|C0231528|Myalgia|myalgias
Finding|Sign or Symptom|History of Present Illness|2194,2200|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Anatomy|Body System|History of Present Illness|2204,2208|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|History of Present Illness|2204,2208|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|History of Present Illness|2204,2208|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|History of Present Illness|2204,2208|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|History of Present Illness|2204,2208|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|History of Present Illness|2204,2218|true|false|false|C0150077;C4048181|Broken skin;Impaired skin integrity|skin breakdown
Disorder|Acquired Abnormality|History of Present Illness|2209,2218|false|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Finding|Organism Function|History of Present Illness|2209,2218|false|false|false|C0699900|Catabolism|breakdown
Finding|Finding|History of Present Illness|2223,2231|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|2223,2231|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|History of Present Illness|2232,2240|true|false|false|C0030554|Paresthesia|tingling
Finding|Sign or Symptom|History of Present Illness|2232,2240|true|false|false|C2242996|Has tingling sensation|tingling
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2245,2256|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Intellectual Product|History of Present Illness|2261,2269|true|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|History of Present Illness|2261,2269|true|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|2273,2283|true|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Finding|Functional Concept|History of Present Illness|2273,2283|true|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|History of Present Illness|2273,2283|true|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|2287,2294|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|History of Present Illness|2287,2294|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|History of Present Illness|2296,2305|false|false|false|C5425799|All other|All other
Finding|Idea or Concept|History of Present Illness|2307,2313|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|2307,2313|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|2307,2316|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|2307,2324|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|2307,2324|false|false|false|C0489633|Review of systems (procedure)|review of systems
Finding|Functional Concept|History of Present Illness|2317,2324|false|false|false|C0449913|System|systems
Finding|Classification|History of Present Illness|2325,2333|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|2325,2333|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|2325,2333|false|false|false|C5237010|Expression Negative|negative
Drug|Organic Chemical|Past Medical History|2364,2371|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Drug|Pharmacologic Substance|Past Medical History|2364,2371|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Finding|Intellectual Product|Past Medical History|2364,2371|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|Alcohol
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2364,2377|false|false|false|C0085762|Alcohol abuse|Alcohol abuse
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2372,2377|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Past Medical History|2372,2377|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Past Medical History|2372,2377|false|false|false|C0562381|Victim of abuse (finding)|abuse
Disorder|Disease or Syndrome|Past Medical History|2382,2401|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|Past Medical History|2392,2401|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Finding|Pathologic Function|Past Medical History|2408,2424|false|false|false|C0476474|Persistent fever|persistent fever
Finding|Finding|Past Medical History|2419,2424|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Past Medical History|2419,2424|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|Past Medical History|2429,2441|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Past Medical History|2429,2441|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Disorder|Disease or Syndrome|Past Medical History|2444,2451|false|false|false|C0003962|Ascites|Ascites
Finding|Pathologic Function|Past Medical History|2444,2451|false|false|false|C5441966|Peritoneal Effusion|Ascites
Finding|Intellectual Product|Past Medical History|2455,2462|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Past Medical History|2455,2462|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|Past Medical History|2455,2472|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|Past Medical History|2463,2472|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Past Medical History|2468,2472|false|false|false|C2598155||pain
Finding|Functional Concept|Past Medical History|2468,2472|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Past Medical History|2468,2472|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Family Medical History|2514,2520|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Neoplastic Process|Family Medical History|2526,2532|false|false|false|C0006826|Malignant Neoplasms|cancer
Attribute|Clinical Attribute|Family Medical History|2534,2537|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|2534,2537|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|2534,2537|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Classification|Family Medical History|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|2549,2563|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|Family Medical History|2549,2566|true|false|false|C0241889|Family Medical History|family history of
Finding|Conceptual Entity|Family Medical History|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2556,2566|true|false|false|C0262926|Medical History|history of
Finding|Finding|Family Medical History|2556,2580|true|false|false|C0455550||history of liver disease
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2567,2572|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|2567,2572|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|2567,2572|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Family Medical History|2567,2572|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|2567,2572|true|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|2567,2580|true|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Family Medical History|2573,2580|true|false|false|C0012634|Disease|disease
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2609,2619|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcoholism
Finding|Finding|General Exam|2639,2647|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|General Exam|2639,2647|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|General Exam|2639,2647|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|General Exam|2639,2652|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|General Exam|2639,2652|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|General Exam|2648,2652|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|2648,2652|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|General Exam|2656,2665|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Classification|General Exam|2669,2672|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|2669,2672|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Disease or Syndrome|General Exam|2674,2677|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2674,2677|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|2674,2677|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Mental or Behavioral Dysfunction|General Exam|2679,2692|false|false|false|C0233472|Labile affect|labile affect
Finding|Mental Process|General Exam|2686,2692|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|2686,2692|false|false|false|C2237113|assessment of affect|affect
Finding|Mental Process|General Exam|2701,2709|false|false|false|C2987187|Pleasant|pleasant
Finding|Finding|General Exam|2714,2721|false|false|false|C0424109|Weepiness|tearful
Anatomy|Body Location or Region|General Exam|2760,2765|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2781,2788|true|false|false|C0221198|Lesion|lesions
Finding|Intellectual Product|General Exam|2790,2794|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|2795,2802|false|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|2795,2810|false|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|General Exam|2803,2810|false|false|false|C0022346|Icterus|icterus
Finding|Gene or Genome|General Exam|2831,2834|true|false|false|C1422304|MAS1L gene|MRG
Procedure|Health Care Activity|General Exam|2837,2841|false|false|false|C1315068|Pulmonary ventilator management|PULM
Finding|Finding|General Exam|2853,2861|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|2870,2873|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|2870,2873|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|2880,2884|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|General Exam|2886,2895|false|false|false|C0700124|Dilated|distended
Finding|Intellectual Product|General Exam|2919,2923|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|2942,2952|false|false|false|C1275670|Collateral branch of vessel|collateral
Anatomy|Body Part, Organ, or Organ Component|General Exam|2953,2958|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|2953,2958|false|false|false|C0398102|Procedure on vein|veins
Finding|Intellectual Product|General Exam|2965,2969|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|2982,2987|false|false|false|C0015385|Limb structure|LIMBS
Finding|Functional Concept|General Exam|2989,2994|false|false|false|C1883002|Sequence Chromatogram|Trace
Attribute|Clinical Attribute|General Exam|2999,3004|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|2999,3004|false|false|false|C0013604|Edema|edema
Finding|Sign or Symptom|General Exam|3009,3016|true|false|false|C0040822|Tremor|tremors
Finding|Sign or Symptom|General Exam|3020,3029|true|false|false|C0232766|Asterixis|asterixis
Anatomy|Body System|General Exam|3032,3036|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Sign or Symptom|General Exam|3041,3047|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Anatomy|Body System|General Exam|3051,3055|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|3051,3055|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|3051,3055|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|3051,3055|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|3051,3055|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|General Exam|3051,3065|true|false|false|C0150077;C4048181|Broken skin;Impaired skin integrity|skin breakdown
Disorder|Acquired Abnormality|General Exam|3056,3065|true|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Finding|Organism Function|General Exam|3056,3065|true|false|false|C0699900|Catabolism|breakdown
Finding|Pathologic Function|General Exam|3077,3087|true|false|false|C0013491|Ecchymosis|ecchymoses
Disorder|Injury or Poisoning|General Exam|3092,3100|false|false|false|C0033119|Puncture wound|puncture
Procedure|Health Care Activity|General Exam|3092,3100|false|false|false|C0034117|Puncture procedure|puncture
Finding|Pathologic Function|General Exam|3132,3146|true|false|false|C1504476|Pronator drift|pronator drift
Finding|Finding|General Exam|3148,3156|true|false|false|C0034929;C0596002|Observation of reflex;Reflex action|reflexes
Finding|Organ or Tissue Function|General Exam|3148,3156|true|false|false|C0034929;C0596002|Observation of reflex;Reflex action|reflexes
Procedure|Diagnostic Procedure|General Exam|3148,3156|true|false|false|C0436145|Examination of reflexes|reflexes
Anatomy|Body Location or Region|General Exam|3182,3187|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|3182,3187|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|3182,3199|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3188,3199|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Lab|Laboratory or Test Result|General Exam|3223,3227|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3230,3235|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|3230,3235|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Anatomy|Cell|General Exam|3241,3244|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3251,3254|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3251,3254|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3251,3254|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3261,3264|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|3261,3264|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|3261,3264|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|3261,3264|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|3271,3274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|3271,3274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|3281,3284|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3281,3284|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3281,3284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3281,3284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3290,3293|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3290,3293|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3290,3293|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3290,3293|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3290,3293|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3301,3305|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3320,3323|false|false|false|C0201617|Primed lymphocyte test|PLT
Disorder|Neoplastic Process|General Exam|3338,3341|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|3338,3341|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Amino Acid, Peptide, or Protein|General Exam|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|General Exam|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|General Exam|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Finding|Gene or Genome|General Exam|3352,3359|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|General Exam|3352,3359|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|General Exam|3352,3359|false|false|false|C0201838|Albumin measurement|ALBUMIN
Disorder|Neoplastic Process|General Exam|3365,3368|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3365,3368|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3365,3368|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3365,3368|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3369,3373|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|3369,3373|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Finding|Gene or Genome|General Exam|3369,3373|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|3369,3373|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|3378,3381|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3378,3381|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|3378,3381|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3382,3386|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|3382,3386|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Finding|Gene or Genome|General Exam|3382,3386|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|3382,3386|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|3393,3396|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|3393,3396|false|false|false|C1663627|ALK protein, human|ALK
Finding|Gene or Genome|General Exam|3393,3396|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|3393,3396|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|General Exam|3393,3401|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|General Exam|3393,3401|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|General Exam|3393,3401|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Finding|Body Substance|General Exam|3422,3435|false|false|false|C5441965|Ascitic Fluid|Ascitic Fluid
Drug|Substance|General Exam|3430,3435|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|General Exam|3430,3435|false|false|false|C1546638|Fluid Specimen Code|Fluid
Anatomy|Cell|General Exam|3443,3446|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3451,3454|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3451,3454|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3451,3454|false|false|false|C0014792|Erythrocytes|RBC
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3459,3464|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|POLYS
Finding|Body Substance|General Exam|3469,3475|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|3488,3491|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|3488,3491|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Finding|Gene or Genome|General Exam|3528,3532|false|false|false|C1420218|SLC6A7 gene|PROT
Drug|Amino Acid, Peptide, or Protein|General Exam|3540,3543|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|3540,3543|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|General Exam|3540,3543|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|3540,3543|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|General Exam|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|General Exam|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Finding|Gene or Genome|General Exam|3548,3555|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|General Exam|3548,3555|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|General Exam|3548,3555|false|false|false|C0201838|Albumin measurement|ALBUMIN
Finding|Body Substance|General Exam|3562,3575|false|false|false|C5441965|Ascitic Fluid|Ascitic Fluid
Drug|Substance|General Exam|3570,3575|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|General Exam|3570,3575|false|false|false|C1546638|Fluid Specimen Code|Fluid
Anatomy|Cell|General Exam|3581,3584|false|false|false|C0023516|Leukocytes|WBC
Finding|Gene or Genome|General Exam|3590,3593|false|false|false|C1428294;C3812663|NACC2 gene;NACC2 wt Allele|RBB
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3599,3604|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|POLYS
Finding|Body Substance|General Exam|3609,3615|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|3629,3632|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|3629,3632|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Disease or Syndrome|General Exam|3654,3659|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|3654,3659|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Anatomy|Cell|General Exam|3665,3668|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|General Exam|3674,3677|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|3674,3677|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Finding|Finding|General Exam|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Idea or Concept|General Exam|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Intellectual Product|General Exam|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Procedure|Diagnostic Procedure|General Exam|3685,3694|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|RADIOLOGY
Anatomy|Body Location or Region|General Exam|3696,3708|false|false|false|C5452879|Lumbo-sacral|Lumbo-sacral
Anatomy|Body Location or Region|General Exam|3702,3708|false|false|false|C0036033;C0036037|Bone structure of sacrum;Sacral Region|sacral
Anatomy|Body Part, Organ, or Organ Component|General Exam|3702,3708|false|false|false|C0036033;C0036037|Bone structure of sacrum;Sacral Region|sacral
Finding|Idea or Concept|General Exam|3724,3732|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|3724,3735|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|General Exam|3736,3749|true|false|false|C0029443|Osteomyelitis|osteomyelitis
Anatomy|Body Part, Organ, or Organ Component|General Exam|3750,3759|false|false|false|C0549207|Bone structure of spine|vertebral
Finding|Functional Concept|General Exam|3761,3772|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|General Exam|3761,3772|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|General Exam|3761,3772|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|General Exam|3761,3772|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|General Exam|3761,3781|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|General Exam|3773,3781|false|false|false|C0016658|Fracture|fracture
Anatomy|Body Location or Region|Hospital Course|3810,3819|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|Hospital Course|3810,3830|false|false|false|C0000731|Abdomen distended|Abdominal distention
Finding|Finding|Hospital Course|3820,3830|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Hospital Course|3820,3830|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|Hospital Course|3831,3835|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3831,3835|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3831,3835|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Hospital Course|3872,3879|false|false|false|C2699424|Concern|concern
Finding|Functional Concept|Hospital Course|3884,3895|false|false|false|C0205359|Spontaneous|spontaneous
Disorder|Disease or Syndrome|Hospital Course|3897,3918|false|false|false|C0275550;C0341503|Acute bacterial peritonitis;Bacterial peritonitis|bacterial peritonitis
Finding|Pathologic Function|Hospital Course|3907,3918|false|false|false|C0031154|Peritonitis|peritonitis
Drug|Antibiotic|Hospital Course|3924,3935|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|3924,3935|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|3947,3957|false|false|false|C0358514|Diagnostic agents|diagnostic
Finding|Functional Concept|Hospital Course|3947,3957|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|Hospital Course|3947,3957|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|Hospital Course|3947,3957|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3959,3971|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Body Substance|Hospital Course|3998,4011|false|false|false|C5441965|Ascitic Fluid|Ascitic fluid
Drug|Substance|Hospital Course|4006,4011|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|4006,4011|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|Hospital Course|4012,4020|false|false|false|C1524024|analysis aspect|analysis
Procedure|Laboratory Procedure|Hospital Course|4012,4020|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Procedure|Research Activity|Hospital Course|4012,4020|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Finding|Functional Concept|Hospital Course|4038,4049|false|false|false|C0205359|Spontaneous|Spontaneous
Disorder|Disease or Syndrome|Hospital Course|4038,4071|false|false|false|C0275551;C2062979|Primary bacterial peritonitis;acute spontaneous bacterial peritonitis|Spontaneous bacterial peritonitis
Disorder|Disease or Syndrome|Hospital Course|4050,4071|false|false|false|C0275550;C0341503|Acute bacterial peritonitis;Bacterial peritonitis|bacterial peritonitis
Finding|Pathologic Function|Hospital Course|4060,4071|false|false|false|C0031154|Peritonitis|peritonitis
Drug|Substance|Hospital Course|4102,4107|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|4102,4107|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Cell|Hospital Course|4108,4112|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|4108,4112|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|Hospital Course|4108,4118|false|false|false|C0007584|Cell Count|cell count
Anatomy|Cell|Hospital Course|4134,4137|false|false|false|C0023516|Leukocytes|WBC
Drug|Antibiotic|Hospital Course|4139,4150|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Mental Process|Hospital Course|4178,4185|false|false|false|C0542559|contextual factors|setting
Finding|Gene or Genome|Hospital Course|4204,4209|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|Hospital Course|4210,4216|false|false|false|C1705102|Volume (publication)|volume
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4218,4230|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Substance|Hospital Course|4265,4271|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|Hospital Course|4265,4271|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4265,4271|false|false|false|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Hospital Course|4292,4301|false|false|false|C0945766||procedure
Event|Occupational Activity|Hospital Course|4292,4301|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|4292,4301|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4292,4301|false|false|false|C0184661|Interventional procedure|procedure
Anatomy|Body Location or Region|Hospital Course|4307,4314|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|4307,4314|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|4307,4314|false|false|false|C0941288|Abdomen problem|abdomen
Finding|Finding|Hospital Course|4324,4333|false|false|false|C0700124|Dilated|distended
Finding|Sign or Symptom|Hospital Course|4344,4351|false|false|false|C0030193|Pain|painful
Drug|Substance|Hospital Course|4354,4359|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|Hospital Course|4354,4359|false|false|false|C1546638|Fluid Specimen Code|Fluid
Finding|Functional Concept|Hospital Course|4360,4368|false|false|false|C1524024|analysis aspect|analysis
Procedure|Laboratory Procedure|Hospital Course|4360,4368|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Procedure|Research Activity|Hospital Course|4360,4368|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Attribute|Clinical Attribute|Hospital Course|4390,4393|true|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4390,4393|true|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|4390,4393|true|false|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|Hospital Course|4390,4393|true|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|4390,4393|true|false|false|C1306620|Systolic blood pressure measurement|SBP
Disorder|Disease or Syndrome|Hospital Course|4400,4419|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|4410,4419|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Finding|Body Substance|Hospital Course|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4431,4436|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|4431,4436|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|4431,4436|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|4431,4436|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|4431,4436|false|false|false|C0872387|Procedures on liver|liver
Event|Activity|Hospital Course|4437,4446|false|false|false|C1883254|Synthesis|synthetic
Finding|Finding|Hospital Course|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Idea or Concept|Hospital Course|4517,4521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4517,4521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4517,4521|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|Hospital Course|4522,4529|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4522,4529|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Organic Chemical|Hospital Course|4534,4543|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|Hospital Course|4534,4543|false|false|false|C0022957|lactulose|lactulose
Finding|Body Substance|Hospital Course|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Procedure|Laboratory Procedure|Hospital Course|4564,4580|false|false|false|C0200354|Urine Specimen Collection|urine collection
Finding|Conceptual Entity|Hospital Course|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Biologically Active Substance|Hospital Course|4585,4591|false|false|false|C0009968|copper|copper
Drug|Element, Ion, or Isotope|Hospital Course|4585,4591|false|false|false|C0009968|copper|copper
Drug|Pharmacologic Substance|Hospital Course|4585,4591|false|false|false|C0009968|copper|copper
Procedure|Laboratory Procedure|Hospital Course|4585,4591|false|false|false|C0373587|Copper measurement|copper
Disorder|Disease or Syndrome|Hospital Course|4613,4620|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Hospital Course|4626,4638|false|false|false|C0023518|Leukocytosis|Leukocytosis
Finding|Finding|Hospital Course|4626,4638|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Finding|Intellectual Product|Hospital Course|4643,4647|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Hospital Course|4643,4653|false|false|false|C0239574|Low grade fever|mild fever
Finding|Finding|Hospital Course|4648,4653|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|4648,4653|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Idea or Concept|Hospital Course|4689,4701|false|false|false|C0449450|Presentation|presentation
Finding|Finding|Hospital Course|4726,4731|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|4726,4731|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|4735,4743|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|4735,4743|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|Hospital Course|4751,4760|true|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|4751,4760|true|false|false|C3714514|Infection|infection
Finding|Body Substance|Hospital Course|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|Hospital Course|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|Hospital Course|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|Hospital Course|4763,4776|false|false|false|C0430404|Urine culture|Urine culture
Drug|Biomedical or Dental Material|Hospital Course|4769,4776|false|false|false|C1706355|Culture Dose Form|culture
Finding|Functional Concept|Hospital Course|4769,4776|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|4769,4776|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|4769,4776|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Idea or Concept|Hospital Course|4800,4810|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|4800,4815|false|false|false|C0332290|Consistent with|consistent with
Finding|Idea or Concept|Hospital Course|4816,4829|false|false|false|C2349974|Contamination|contamination
Phenomenon|Human-caused Phenomenon or Process|Hospital Course|4816,4829|false|false|false|C0259846|adulteration|contamination
Event|Activity|Hospital Course|4837,4844|false|false|false|C1706079||arrival
Finding|Functional Concept|Hospital Course|4837,4844|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|Hospital Course|4853,4858|false|false|false|C3714591|Floor (anatomic)|floor
Procedure|Health Care Activity|Hospital Course|4863,4874|false|false|false|C0886414|Body temperature measurement|temperature
Finding|Intellectual Product|Hospital Course|4879,4885|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Cell|Hospital Course|4917,4920|false|false|false|C0023516|Leukocytes|WBC
Procedure|Health Care Activity|Hospital Course|4949,4964|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Finding|Hospital Course|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4992,5001|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|5010,5021|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|Tachycardia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5027,5032|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|5027,5032|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|5027,5032|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Hospital Course|5027,5037|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Hospital Course|5027,5037|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Hospital Course|5027,5037|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Hospital Course|5033,5037|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|5033,5037|false|false|false|C1549480|Amount type - Rate|rate
Procedure|Health Care Activity|Hospital Course|5083,5098|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Idea or Concept|Hospital Course|5108,5112|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Cell Function|Hospital Course|5113,5124|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Organ or Tissue Function|Hospital Course|5113,5124|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Finding|Hospital Course|5136,5146|true|false|false|C5441521|Complaint (finding)|complaints
Finding|Sign or Symptom|Hospital Course|5151,5154|false|false|false|C0013404|Dyspnea|SOB
Finding|Finding|Hospital Course|5156,5163|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5156,5163|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Anatomy|Body Location or Region|Hospital Course|5165,5170|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|5165,5170|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|5165,5175|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|5165,5175|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|5171,5175|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5171,5175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5171,5175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|5177,5189|false|false|false|C0030252|Palpitations|palpitations
Finding|Idea or Concept|Hospital Course|5195,5206|false|false|false|C0750501|most likely|most likely
Finding|Finding|Hospital Course|5200,5206|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|5200,5206|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Conceptual Entity|Hospital Course|5208,5216|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|Hospital Course|5208,5216|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Attribute|Clinical Attribute|Hospital Course|5228,5232|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5228,5232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5228,5232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5234,5241|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|5234,5241|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|Hospital Course|5251,5254|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|5251,5254|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Functional Concept|Hospital Course|5255,5268|false|false|false|C2960476|Intravascular Route of Administration|intravascular
Finding|Intellectual Product|Hospital Course|5270,5276|false|false|false|C1705102|Volume (publication)|volume
Finding|Body Substance|Hospital Course|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5316,5325|false|false|false|C0030685|Patient Discharge|discharge
Finding|Sign or Symptom|Hospital Course|5332,5341|false|false|false|C0004604|Back Pain|Back pain
Attribute|Clinical Attribute|Hospital Course|5337,5341|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5337,5341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5337,5341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5343,5360|false|false|false|C0223603|Lumbosacral spine|Lumbosacral spine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5355,5360|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Hospital Course|5355,5360|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Hospital Course|5355,5360|false|false|false|C0150920|Spine Problem|spine
Drug|Biomedical or Dental Material|Hospital Course|5361,5365|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Drug|Substance|Hospital Course|5361,5365|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Finding|Intellectual Product|Hospital Course|5361,5365|false|false|false|C4019020||film
Disorder|Anatomical Abnormality|Hospital Course|5378,5400|true|false|false|C4021790|Abnormality of the skeletal system|skeletal abnormalities
Disorder|Congenital Abnormality|Hospital Course|5387,5400|true|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|Hospital Course|5387,5400|true|false|false|C0000769|teratologic|abnormalities
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5403,5412|false|false|false|C0549207|Bone structure of spine|vertebral
Finding|Pathologic Function|Hospital Course|5403,5424|false|false|false|C0262431|Compression fracture of vertebral column|vertebral compression
Finding|Pathologic Function|Hospital Course|5403,5433|false|false|false|C0262431|Compression fracture of vertebral column|vertebral compression fracture
Finding|Functional Concept|Hospital Course|5413,5424|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|5413,5424|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|5413,5424|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5413,5424|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|Hospital Course|5413,5433|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|Hospital Course|5425,5433|false|false|false|C0016658|Fracture|fracture
Disorder|Disease or Syndrome|Hospital Course|5438,5451|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Attribute|Clinical Attribute|Hospital Course|5459,5463|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5459,5463|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5459,5463|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|5469,5476|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Hospital Course|5469,5476|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Finding|Hospital Course|5481,5485|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|Hospital Course|5512,5527|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Organic Chemical|Hospital Course|5534,5543|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|5534,5543|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|Hospital Course|5534,5543|false|false|false|C0524222|Oxycodone measurement|oxycodone
Finding|Gene or Genome|Hospital Course|5552,5555|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5556,5560|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5556,5560|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5556,5560|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|Hospital Course|5595,5607|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|5595,5607|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|Hospital Course|5595,5616|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|Hospital Course|5595,5616|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|Hospital Course|5603,5607|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|5603,5607|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|5603,5607|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Hospital Course|5608,5616|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|5608,5616|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Occupational Activity|Hospital Course|5628,5638|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|5628,5638|false|false|false|C0376636|Disease Management|management
Finding|Intellectual Product|Hospital Course|5646,5653|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|5646,5653|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|Hospital Course|5655,5659|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5655,5659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5655,5659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Food|Hospital Course|5665,5669|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Finding|Functional Concept|Hospital Course|5665,5669|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|Hospital Course|5665,5669|false|false|false|C0012159|Diet therapy|Diet
Finding|Finding|Hospital Course|5671,5674|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Hospital Course|5671,5674|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Finding|Hospital Course|5671,5681|false|false|false|C0860871|Sodium decreased|Low sodium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5671,5681|false|false|false|C0012169|Low sodium diet|Low sodium
Drug|Biologically Active Substance|Hospital Course|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|Hospital Course|5675,5681|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|5675,5681|false|false|false|C0337443|Sodium measurement|sodium
Finding|Idea or Concept|Hospital Course|5686,5689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5686,5689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Substance|Hospital Course|5692,5697|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|5692,5697|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5692,5709|false|false|false|C0204700|Fluid restriction|fluid restriction
Finding|Functional Concept|Hospital Course|5698,5709|false|false|false|C0443288|Restricted|restriction
Finding|Idea or Concept|Hospital Course|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Occupational Activity|Hospital Course|5726,5730|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|5726,5730|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Attribute|Clinical Attribute|Hospital Course|5740,5751|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5740,5751|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|5740,5751|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5740,5764|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|5755,5764|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|5768,5781|false|false|false|C0002600|amitriptyline|AMITRIPTYLINE
Drug|Pharmacologic Substance|Hospital Course|5768,5781|false|false|false|C0002600|amitriptyline|AMITRIPTYLINE
Drug|Organic Chemical|Hospital Course|5800,5809|false|false|false|C0030049|oxycodone|OXYCODONE
Drug|Pharmacologic Substance|Hospital Course|5800,5809|false|false|false|C0030049|oxycodone|OXYCODONE
Procedure|Laboratory Procedure|Hospital Course|5800,5809|false|false|false|C0524222|Oxycodone measurement|OXYCODONE
Finding|Gene or Genome|Hospital Course|5824,5827|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5828,5832|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5828,5832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5828,5832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|Hospital Course|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|Hospital Course|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Procedure|Laboratory Procedure|Hospital Course|5837,5845|false|false|false|C0373727|Thiamine measurement|Thiamine
Drug|Organic Chemical|Hospital Course|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Drug|Pharmacologic Substance|Hospital Course|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Drug|Vitamin|Hospital Course|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Procedure|Laboratory Procedure|Hospital Course|5865,5875|false|false|false|C0523631|Folic acid measurement|Folic acid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5893,5896|false|false|false|C5417720|MVI Regimen|MVI
Finding|Body Substance|Hospital Course|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5910,5919|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5910,5931|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|5920,5931|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5920,5931|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|5920,5931|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|Hospital Course|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|Hospital Course|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Procedure|Laboratory Procedure|Hospital Course|5936,5944|false|false|false|C0373727|Thiamine measurement|Thiamine
Drug|Organic Chemical|Hospital Course|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Pharmacologic Substance|Hospital Course|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Vitamin|Hospital Course|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Disorder|Neoplastic Process|Hospital Course|5945,5948|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Biomedical or Dental Material|Hospital Course|5956,5962|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5976,5982|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Drug|Pharmacologic Substance|Hospital Course|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Drug|Vitamin|Hospital Course|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Procedure|Laboratory Procedure|Hospital Course|6005,6015|false|false|false|C0523631|Folic acid measurement|Folic Acid
Drug|Biomedical or Dental Material|Hospital Course|6021,6027|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6041,6047|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6072,6085|false|false|false|C0002600|amitriptyline|Amitriptyline
Drug|Pharmacologic Substance|Hospital Course|6072,6085|false|false|false|C0002600|amitriptyline|Amitriptyline
Drug|Biomedical or Dental Material|Hospital Course|6092,6098|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6112,6118|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|6145,6168|false|false|false|C0978787|Multivitamin tablet|Multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|6162,6168|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6182,6188|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6213,6222|true|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|Hospital Course|6213,6222|true|false|false|C0022957|lactulose|Lactulose
Drug|Biomedical or Dental Material|Hospital Course|6237,6242|true|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|Syrup
Drug|Food|Hospital Course|6237,6242|true|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|Syrup
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6243,6246|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Organic Chemical|Hospital Course|6287,6296|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|6287,6296|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|Hospital Course|6287,6296|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Biomedical or Dental Material|Hospital Course|6302,6308|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6322,6328|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|Hospital Course|6369,6373|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6369,6373|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6369,6373|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|Hospital Course|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6380,6389|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6380,6401|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6380,6401|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6390,6401|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|6390,6401|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|6403,6407|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6403,6407|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6403,6407|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6410,6419|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6410,6429|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6420,6429|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|6420,6429|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6420,6429|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6420,6429|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|6440,6447|false|false|false|C0003962|Ascites|Ascites
Finding|Pathologic Function|Hospital Course|6440,6447|false|false|false|C5441966|Peritoneal Effusion|Ascites
Anatomy|Body Location or Region|Hospital Course|6448,6454|false|false|false|C0205054|Hepatic|Portal
Disorder|Disease or Syndrome|Hospital Course|6448,6467|false|false|false|C0020541|Portal Hypertension|Portal hypertension
Disorder|Disease or Syndrome|Hospital Course|6455,6467|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Hospital Course|6468,6487|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|6478,6487|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Disorder|Neoplastic Process|Hospital Course|6490,6499|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|6490,6499|false|false|false|C1522484|metastatic qualifier|Secondary
Finding|Intellectual Product|Hospital Course|6501,6508|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|6501,6508|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|Hospital Course|6501,6518|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|Hospital Course|6509,6518|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Hospital Course|6514,6518|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6514,6518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6514,6518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Condition|6543,6548|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|6543,6548|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|6543,6548|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Finding|Discharge Condition|6553,6561|false|false|false|C1961028|Oriented to place|Oriented
Finding|Intellectual Product|Discharge Condition|6575,6587|false|false|false|C3827452|Without Help|without help
Finding|Intellectual Product|Discharge Condition|6583,6587|true|false|false|C1552861|Help document|help
Finding|Intellectual Product|Discharge Condition|6607,6613|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|Discharge Condition|6615,6623|false|false|false|C0277797|Apyrexial|afebrile
Finding|Finding|Discharge Instructions|6709,6719|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Functional Concept|Discharge Instructions|6723,6733|false|false|false|C0442808|Increasing (qualifier value)|increasing
Anatomy|Body Location or Region|Discharge Instructions|6734,6743|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|Discharge Instructions|6734,6754|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|Discharge Instructions|6734,6763|false|false|false|C2749840|Abdominal distention and pain|abdominal distention and pain
Finding|Finding|Discharge Instructions|6744,6754|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Discharge Instructions|6744,6754|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|Discharge Instructions|6759,6763|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|6759,6763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6759,6763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|Discharge Instructions|6796,6800|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Discharge Instructions|6796,6806|false|false|false|C0239574|Low grade fever|mild fever
Finding|Finding|Discharge Instructions|6801,6806|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|6801,6806|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Finding|Discharge Instructions|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|Discharge Instructions|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|Discharge Instructions|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|Discharge Instructions|6808,6823|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6813,6818|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|6813,6818|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|6813,6818|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|6813,6823|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|6813,6823|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|6813,6823|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|6819,6823|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|6819,6823|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Discharge Instructions|6840,6857|false|false|false|C1821144|White blood count|white blood count
Disorder|Disease or Syndrome|Discharge Instructions|6846,6851|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|6846,6851|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|6846,6857|false|false|false|C0005771|Blood Cell Count|blood count
Finding|Finding|Discharge Instructions|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|6881,6890|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|6881,6890|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Discharge Instructions|6892,6902|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Finding|Idea or Concept|Discharge Instructions|6923,6931|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Health Care Activity|Discharge Instructions|6965,6980|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Body Substance|Discharge Instructions|6986,6999|false|false|false|C5441965|Ascitic Fluid|ascitic fluid
Drug|Substance|Discharge Instructions|6994,6999|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|6994,6999|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|Discharge Instructions|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|Discharge Instructions|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|Discharge Instructions|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Disorder|Disease or Syndrome|Discharge Instructions|7070,7079|true|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|7070,7079|true|false|false|C3714514|Infection|infection
Finding|Body Substance|Discharge Instructions|7088,7101|false|false|false|C5441965|Ascitic Fluid|ascitic fluid
Drug|Substance|Discharge Instructions|7096,7101|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|7096,7101|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Substance|Discharge Instructions|7118,7123|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|7118,7123|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Discharge Instructions|7147,7154|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Discharge Instructions|7147,7154|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Discharge Instructions|7147,7154|false|false|false|C0941288|Abdomen problem|abdomen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7159,7171|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Body Substance|Discharge Instructions|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Discharge Instructions|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Discharge Instructions|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Conceptual Entity|Discharge Instructions|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Discharge Instructions|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Discharge Instructions|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Discharge Instructions|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Biologically Active Substance|Discharge Instructions|7219,7225|false|false|false|C0009968|copper|copper
Drug|Element, Ion, or Isotope|Discharge Instructions|7219,7225|false|false|false|C0009968|copper|copper
Drug|Pharmacologic Substance|Discharge Instructions|7219,7225|false|false|false|C0009968|copper|copper
Procedure|Laboratory Procedure|Discharge Instructions|7219,7225|false|false|false|C0373587|Copper measurement|copper
Finding|Functional Concept|Discharge Instructions|7257,7263|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7273,7278|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|7273,7278|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|7273,7278|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|7273,7278|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|7273,7278|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|7273,7286|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Discharge Instructions|7279,7286|false|false|false|C0012634|Disease|disease
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7293,7298|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|7293,7298|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|7293,7298|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|7293,7298|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|7293,7298|false|false|false|C0872387|Procedures on liver|liver
Finding|Intellectual Product|Discharge Instructions|7362,7367|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|Discharge Instructions|7362,7367|false|false|false|C0022885|Laboratory Procedures|tests
Finding|Sign or Symptom|Discharge Instructions|7378,7387|false|false|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Discharge Instructions|7383,7387|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7383,7387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7383,7387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Health Care Activity|Discharge Instructions|7410,7425|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Pharmacologic Substance|Discharge Instructions|7443,7449|false|false|false|C0885876|X-rays, Homeopathic Preparations|x-rays
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|7443,7449|false|false|false|C0043309|Roentgen Rays|x-rays
Procedure|Diagnostic Procedure|Discharge Instructions|7443,7449|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|x-rays
Finding|Idea or Concept|Discharge Instructions|7466,7474|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|7466,7477|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Injury or Poisoning|Discharge Instructions|7478,7486|true|false|false|C0016658|Fracture|fracture
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7490,7494|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|Discharge Instructions|7490,7494|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|Discharge Instructions|7490,7494|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Disease or Syndrome|Discharge Instructions|7496,7505|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|7496,7505|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|Discharge Instructions|7529,7533|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|7529,7533|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|7529,7533|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|7534,7538|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7534,7538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7534,7538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|Discharge Instructions|7539,7546|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7539,7546|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Intellectual Product|Discharge Instructions|7572,7584|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|7572,7584|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|Discharge Instructions|7572,7593|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|Discharge Instructions|7572,7593|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|Discharge Instructions|7580,7584|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|7580,7584|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|7580,7584|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Discharge Instructions|7585,7593|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Discharge Instructions|7585,7593|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Functional Concept|Discharge Instructions|7600,7607|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|Discharge Instructions|7626,7630|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|7626,7630|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|7626,7630|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|7631,7642|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7631,7642|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|7631,7642|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Discharge Instructions|7673,7682|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|Discharge Instructions|7673,7682|false|false|false|C0022957|lactulose|lactulose
Finding|Sign or Symptom|Discharge Instructions|7687,7699|false|false|false|C0009806|Constipation|constipation
Attribute|Clinical Attribute|Discharge Instructions|7712,7716|false|true|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7712,7716|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7712,7716|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|7718,7729|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7718,7729|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|7718,7729|false|false|false|C4284232|Medications|medications
Finding|Intellectual Product|Discharge Instructions|7757,7763|false|false|false|C0376667|Herbals (publications)|herbal
Drug|Pharmacologic Substance|Discharge Instructions|7767,7772|false|false|false|C3543842|TONICS|tonic
Drug|Pharmacologic Substance|Discharge Instructions|7773,7781|false|false|false|C0920324|Homeopathic Remedies|remedies
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7793,7798|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|7793,7798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|7793,7798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|7793,7798|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|7793,7798|false|false|false|C0872387|Procedures on liver|liver
Finding|Finding|Discharge Instructions|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Discharge Instructions|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Discharge Instructions|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Discharge Instructions|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7838,7847|false|false|false|C0087111|Therapeutic procedure|therapies
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|7872,7879|false|false|false|C1705970|Electrical Current|current
Attribute|Clinical Attribute|Discharge Instructions|7880,7891|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7880,7891|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|7880,7891|false|false|false|C4284232|Medications|medications
Finding|Finding|Discharge Instructions|7903,7912|false|false|false|C0332218|Difficult (qualifier value)|difficult
Attribute|Clinical Attribute|Discharge Instructions|7932,7942|false|false|false|C2598148||laboratory
Finding|Functional Concept|Discharge Instructions|7932,7942|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Finding|Intellectual Product|Discharge Instructions|7932,7942|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Lab|Laboratory or Test Result|Discharge Instructions|7932,7942|false|false|false|C4283904|Laboratory observation|laboratory
Lab|Laboratory or Test Result|Discharge Instructions|7932,7950|false|false|false|C1254595|Laboratory Results|laboratory results
Procedure|Health Care Activity|Discharge Instructions|7954,7962|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7963,7975|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|7963,7975|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

