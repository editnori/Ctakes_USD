 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|Allergies|184,193|true|false|false|C1717415||Allergies
Event|Event|Allergies|184,193|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|184,193|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|196,218|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|204,208|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|204,208|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|204,218|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|209,218|true|false|false|||Reactions
Event|Event|Allergies|221,230|false|false|false|||Attending
Finding|Functional Concept|Allergies|221,230|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|256,265|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Chief Complaint|256,270|false|false|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Chief Complaint|266,270|false|false|false|C2598155||pain
Event|Event|Chief Complaint|266,270|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|266,270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|266,270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Chief Complaint|272,282|false|false|false|||distention
Finding|Finding|Chief Complaint|272,282|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Chief Complaint|272,282|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|Chief Complaint|284,290|false|false|false|C4255480||nausea
Event|Event|Chief Complaint|284,290|false|false|false|||nausea
Finding|Sign or Symptom|Chief Complaint|284,290|false|false|false|C0027497|Nausea|nausea
Finding|Classification|Chief Complaint|293,298|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|299,307|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|299,307|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|311,329|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|320,329|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|320,329|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|320,329|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|320,329|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|320,329|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|Chief Complaint|331,345|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|Interventional
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|331,345|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|Interventional
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|331,355|false|false|false|C0344093|Interventional Radiology Procedure|Interventional radiology
Event|Event|Chief Complaint|346,355|false|false|false|||radiology
Finding|Finding|Chief Complaint|346,355|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Finding|Idea or Concept|Chief Complaint|346,355|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Finding|Intellectual Product|Chief Complaint|346,355|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Procedure|Diagnostic Procedure|Chief Complaint|346,355|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|radiology
Event|Event|Chief Complaint|356,365|false|false|false|||placement
Procedure|Health Care Activity|Chief Complaint|356,365|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|356,365|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Anatomy|Body Location or Region|Chief Complaint|369,378|false|false|false|C0000726|Abdomen|abdominal
Disorder|Disease or Syndrome|Chief Complaint|369,386|false|false|false|C0243001|Abdominal Abscess|abdominal abscess
Disorder|Disease or Syndrome|Chief Complaint|379,386|false|false|false|C0000833|Abscess|abscess
Event|Event|Chief Complaint|379,386|false|false|false|||abscess
Finding|Intellectual Product|Chief Complaint|379,386|false|false|false|C1546533||abscess
Drug|Substance|Chief Complaint|387,392|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Chief Complaint|387,392|false|false|false|||drain
Finding|Intellectual Product|Chief Complaint|387,392|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|439,445|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|History of Present Illness|439,445|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Disorder|Neoplastic Process|History of Present Illness|446,469|false|false|false|C1827293|Carcinoma of urinary bladder, invasive|invasive bladder cancer
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|455,462|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|455,462|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|455,462|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|455,469|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|History of Present Illness|463,469|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|463,469|false|false|false|||cancer
Event|Event|History of Present Illness|471,480|false|false|false|||returning
Anatomy|Body Location or Region|History of Present Illness|504,513|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|504,518|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|514,518|false|false|false|C2598155||pain
Event|Event|History of Present Illness|514,518|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|514,518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|514,518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|520,526|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|520,526|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|520,526|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|532,542|false|false|false|||distension
Finding|Finding|History of Present Illness|532,542|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|History of Present Illness|532,542|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Event|Event|History of Present Illness|558,568|false|false|false|||obstipated
Procedure|Diagnostic Procedure|History of Present Illness|600,607|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|History of Present Illness|603,607|false|false|false|||scan
Procedure|Diagnostic Procedure|History of Present Illness|603,607|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|History of Present Illness|609,616|false|false|false|||notable
Finding|Finding|History of Present Illness|621,628|false|false|false|C0700124|Dilated|dilated
Finding|Finding|History of Present Illness|621,634|false|false|false|C4697734|Dilated loops|dilated loops
Event|Event|History of Present Illness|629,634|false|false|false|||loops
Drug|Inorganic Chemical|History of Present Illness|636,639|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|History of Present Illness|636,639|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|History of Present Illness|636,639|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|History of Present Illness|636,639|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|History of Present Illness|636,639|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|History of Present Illness|636,639|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Substance|History of Present Illness|640,646|true|false|false|C0302908|Liquid substance|fluids
Event|Event|History of Present Illness|640,646|true|false|false|||fluids
Finding|Body Substance|History of Present Illness|640,646|true|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|640,646|true|false|false|C0016286|Fluid Therapy|fluids
Event|Event|History of Present Illness|652,660|true|false|false|||tapering
Anatomy|Body Location or Region|History of Present Illness|661,672|true|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|661,672|true|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|667,672|true|false|false|C0021853|Intestines|bowel
Disorder|Cell or Molecular Dysfunction|History of Present Illness|693,703|true|false|false|C0599156|Transition Mutation|transition
Event|Activity|History of Present Illness|693,703|true|false|false|C2700061|Transition (action)|transition
Event|Event|History of Present Illness|693,703|true|false|false|||transition
Finding|Functional Concept|History of Present Illness|693,709|true|false|false|C4684447|Transition Point|transition point
Disorder|Disease or Syndrome|History of Present Illness|740,752|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|History of Present Illness|740,752|false|false|false|||leukocytosis
Finding|Finding|History of Present Illness|740,752|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Anatomy|Body Location or Region|History of Present Illness|768,779|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|768,779|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Disorder|Disease or Syndrome|History of Present Illness|768,791|false|false|false|C0235329|Small bowel obstruction|small bowel obstruction
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|774,779|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|History of Present Illness|774,791|false|false|false|C0021843|Intestinal Obstruction|bowel obstruction
Event|Event|History of Present Illness|780,791|false|false|false|||obstruction
Finding|Finding|History of Present Illness|780,791|false|false|false|C0028778|Obstruction|obstruction
Disorder|Disease or Syndrome|History of Present Illness|798,803|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|History of Present Illness|798,803|false|false|false|||ileus
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|808,816|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Disorder|Disease or Syndrome|History of Present Illness|825,837|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|History of Present Illness|825,837|false|false|false|||leukocytosis
Finding|Finding|History of Present Illness|825,837|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|History of Present Illness|846,857|false|false|false|||re-admitted
Anatomy|Body Space or Junction|History of Present Illness|862,865|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|History of Present Illness|862,865|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|History of Present Illness|862,865|false|false|false|||IVF
Finding|Gene or Genome|History of Present Illness|862,865|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|862,865|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|868,873|false|false|false|C0021853|Intestines|bowel
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|874,878|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|874,878|false|false|false|C1742913|REST protein, human|rest
Event|Event|History of Present Illness|874,878|false|false|false|||rest
Finding|Daily or Recreational Activity|History of Present Illness|874,878|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|874,878|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|874,878|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|History of Present Illness|884,897|false|false|false|||decompression
Finding|Functional Concept|History of Present Illness|884,897|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|History of Present Illness|884,897|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|884,897|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Disorder|Disease or Syndrome|Past Medical History|924,936|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|924,936|false|false|false|||Hypertension
Procedure|Diagnostic Procedure|Past Medical History|938,950|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|Past Medical History|938,966|false|false|false|C0162522|Cholecystectomy, Laparoscopic|laparoscopic cholecystectomy
Event|Event|Past Medical History|951,966|false|false|false|||cholecystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|951,966|false|false|false|C0008320|Cholecystectomy procedure|cholecystectomy
Finding|Functional Concept|Past Medical History|968,972|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Past Medical History|968,977|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|968,977|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|Past Medical History|973,977|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|973,977|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Past Medical History|973,977|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Past Medical History|973,977|false|false|false|C0562271|Examination of knee joint|knee
Event|Event|Past Medical History|979,990|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|979,990|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|979,990|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|979,990|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Gene or Genome|Past Medical History|1008,1011|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Past Medical History|1013,1024|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1013,1024|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|Past Medical History|1037,1040|false|false|false|C1114365||age
Drug|Biologically Active Substance|Past Medical History|1037,1040|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Past Medical History|1037,1040|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Past Medical History|1037,1040|false|false|false|||age
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1051,1058|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|1051,1058|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|1051,1058|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|1051,1058|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|Past Medical History|1059,1069|false|false|false|||deliveries
Event|Event|Past Medical History|1101,1113|false|false|false|||laparoscopic
Procedure|Diagnostic Procedure|Past Medical History|1101,1113|false|false|false|C0031150|Laparoscopy|laparoscopic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1124,1130|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1124,1141|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|Past Medical History|1131,1136|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1131,1141|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|Past Medical History|1143,1153|false|false|false|||dissection
Finding|Pathologic Function|Past Medical History|1143,1153|false|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1143,1153|false|false|false|C0012737|Tissue Dissection|dissection
Event|Event|Past Medical History|1173,1185|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|1173,1185|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1173,1185|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1190,1212|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|Past Medical History|1200,1212|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1200,1212|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|Past Medical History|1218,1223|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|Past Medical History|1218,1230|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1224,1230|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|Past Medical History|1224,1230|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|Past Medical History|1224,1230|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|Past Medical History|1224,1230|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|Past Medical History|1224,1230|false|false|false|||uterus
Procedure|Diagnostic Procedure|Past Medical History|1224,1230|false|false|false|C0869889|examination of uterus|uterus
Finding|Gene or Genome|Past Medical History|1261,1266|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Neoplastic Process|Past Medical History|1267,1274|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|Past Medical History|1267,1274|false|false|false|||fibroid
Procedure|Diagnostic Procedure|Past Medical History|1279,1291|false|false|false|C0031150|Laparoscopy|Laparoscopic
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1279,1310|false|false|false|C5879917|Laparoscopic radical cystectomy|Laparoscopic radical cystectomy
Drug|Chemical Viewed Structurally|Past Medical History|1292,1299|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1292,1310|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|Past Medical History|1300,1310|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1300,1310|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|Past Medical History|1315,1323|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Past Medical History|1324,1335|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1324,1335|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1342,1349|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|1342,1349|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|1342,1349|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|1342,1349|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1342,1364|false|false|false|C0195196|Reconstruction of vagina|vaginal reconstruction
Event|Event|Past Medical History|1350,1364|false|false|false|||reconstruction
Procedure|Machine Activity|Past Medical History|1350,1364|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1350,1364|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Event|Event|Family Medical History|1405,1413|false|false|false|||Negative
Finding|Classification|Family Medical History|1405,1413|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Family Medical History|1405,1413|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Family Medical History|1405,1413|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|Family Medical History|1405,1417|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1418,1425|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Family Medical History|1418,1425|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Family Medical History|1418,1425|true|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1418,1425|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Family Medical History|1418,1428|true|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Disorder|Disease or Syndrome|General Exam|1454,1457|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1454,1457|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1454,1457|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1454,1457|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1454,1457|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1454,1457|false|false|false|||NAD
Finding|Finding|General Exam|1454,1457|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|1459,1463|false|false|false|||AVSS
Anatomy|Body Location or Region|General Exam|1464,1471|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|1464,1471|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|1464,1471|false|false|false|C0941288|Abdomen problem|Abdomen
Finding|Finding|General Exam|1464,1476|false|false|false|C0426663|Abdomen soft|Abdomen soft
Disorder|Disease or Syndrome|General Exam|1472,1476|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|1472,1476|false|false|false|||soft
Anatomy|Body Location or Region|General Exam|1505,1513|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|General Exam|1505,1513|false|false|false|C0332803|Surgical wound|incision
Event|Event|General Exam|1505,1513|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|General Exam|1505,1513|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|General Exam|1514,1522|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|General Exam|1514,1522|false|false|false|C0332803|Surgical wound|Incision
Event|Event|General Exam|1514,1522|false|false|false|||Incision
Procedure|Therapeutic or Preventive Procedure|General Exam|1514,1522|false|false|false|C0184898|Surgical incisions|Incision
Anatomy|Anatomical Structure|General Exam|1532,1537|false|false|false|C1955856|Surgical Stoma|Stoma
Finding|Finding|General Exam|1541,1545|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|General Exam|1556,1561|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|General Exam|1556,1561|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|General Exam|1556,1561|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Finding|General Exam|1556,1567|false|false|false|C0278030|Color of urine|Urine color
Drug|Biomedical or Dental Material|General Exam|1562,1567|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|1562,1567|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Event|Event|General Exam|1562,1567|false|false|false|||color
Event|Event|General Exam|1571,1577|false|false|false|||yellow
Anatomy|Body Location or Region|General Exam|1588,1593|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|1588,1593|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|1588,1605|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|1594,1605|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|1610,1614|false|false|false|||warm
Finding|Finding|General Exam|1610,1614|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|1610,1614|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|1621,1625|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1626,1634|false|false|false|||perfused
Event|Event|General Exam|1650,1658|true|false|false|||reported
Anatomy|Body Location or Region|General Exam|1659,1663|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|1659,1663|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|General Exam|1659,1668|true|false|false|C0236040|Pain in calf|calf pain
Attribute|Clinical Attribute|General Exam|1664,1668|true|false|false|C2598155||pain
Event|Event|General Exam|1664,1668|true|false|false|||pain
Finding|Functional Concept|General Exam|1664,1668|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|1664,1668|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|General Exam|1672,1676|true|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|General Exam|1672,1686|true|false|false|C0278328|Deep palpation|deep palpation
Event|Event|General Exam|1677,1686|true|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|1677,1686|true|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|1698,1703|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|1698,1703|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|1705,1716|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Finding|General Exam|1722,1738|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|General Exam|1725,1732|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|1725,1738|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|1733,1738|false|false|false|C1717255||edema
Event|Event|General Exam|1733,1738|false|false|false|||edema
Finding|Pathologic Function|General Exam|1733,1738|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|General Exam|1746,1754|true|false|false|C0041834|Erythema|erythema
Event|Event|General Exam|1746,1754|true|false|false|||erythema
Event|Event|General Exam|1756,1762|true|false|false|||callor
Attribute|Clinical Attribute|General Exam|1764,1768|true|false|false|C2598155||pain
Event|Event|General Exam|1764,1768|true|false|false|||pain
Finding|Functional Concept|General Exam|1764,1768|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|1764,1768|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Substance|General Exam|1780,1785|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|General Exam|1780,1785|false|false|false|||drain
Finding|Intellectual Product|General Exam|1780,1785|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|General Exam|1795,1802|false|false|false|||removed
Drug|Biomedical or Dental Material|General Exam|1805,1813|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|General Exam|1805,1813|false|false|false|||dressing
Finding|Daily or Recreational Activity|General Exam|1805,1813|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|General Exam|1805,1813|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|General Exam|1805,1813|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|General Exam|1805,1813|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Disorder|Disease or Syndrome|General Exam|1853,1858|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1853,1858|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1853,1858|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1859,1862|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1867,1870|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1867,1870|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1867,1870|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1877,1880|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1877,1880|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1877,1880|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1877,1880|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1886,1889|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1886,1889|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1897,1900|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|1897,1900|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|1897,1900|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1897,1900|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1897,1900|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1904,1907|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1904,1907|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|1904,1907|false|false|false|||MCH
Finding|Gene or Genome|General Exam|1904,1907|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1904,1907|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1904,1907|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|1913,1917|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|1913,1917|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|1945,1948|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|1965,1970|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1965,1970|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1965,1970|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1971,1974|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1981,1984|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1981,1984|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1981,1984|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1991,1994|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1991,1994|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1991,1994|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1991,1994|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2000,2003|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2000,2003|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2011,2014|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2011,2014|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2011,2014|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2011,2014|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2011,2014|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2018,2021|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2018,2021|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2018,2021|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2018,2021|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2018,2021|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2018,2021|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2027,2031|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2027,2031|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2059,2062|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2079,2084|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2079,2084|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2079,2084|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2085,2088|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2095,2098|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2095,2098|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2095,2098|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2105,2108|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2105,2108|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2105,2108|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2105,2108|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2114,2117|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2114,2117|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2125,2128|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2125,2128|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2125,2128|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2125,2128|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2125,2128|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2132,2135|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2132,2135|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2132,2135|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2132,2135|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2132,2135|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2132,2135|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2141,2145|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2141,2145|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2173,2176|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2193,2198|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2193,2198|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2193,2198|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2199,2202|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2210,2213|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2210,2213|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2210,2213|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2220,2223|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2220,2223|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2220,2223|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2220,2223|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2230,2233|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2230,2233|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2240,2243|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2240,2243|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2240,2243|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2240,2243|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2240,2243|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2247,2250|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2247,2250|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2247,2250|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2247,2250|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2247,2250|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2247,2250|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2256,2260|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2256,2260|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2287,2290|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2307,2312|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2307,2312|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2307,2312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|2331,2337|false|false|false|||Lymphs
Finding|Body Substance|General Exam|2331,2337|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|2341,2346|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|2341,2346|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|2341,2346|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|2351,2354|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|2351,2354|false|false|false|||Eos
Finding|Gene or Genome|General Exam|2351,2354|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|2479,2484|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2479,2484|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2479,2484|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2489,2492|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|2489,2492|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|2489,2492|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2514,2519|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2514,2519|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2514,2519|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2514,2527|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2514,2527|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2514,2527|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2520,2527|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2520,2527|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2520,2527|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2520,2527|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2520,2527|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2520,2527|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2574,2578|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2574,2578|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2574,2578|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2602,2607|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2602,2607|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2602,2607|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2602,2615|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2602,2615|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2602,2615|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2608,2615|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2608,2615|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2608,2615|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2608,2615|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2608,2615|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2608,2615|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2662,2666|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2662,2666|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2662,2666|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2691,2696|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2691,2696|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2691,2696|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2691,2704|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2691,2704|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2691,2704|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2697,2704|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2697,2704|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2697,2704|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2697,2704|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2697,2704|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2697,2704|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2751,2755|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2751,2755|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2751,2755|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2780,2785|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2780,2785|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2780,2785|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2780,2793|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2780,2793|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2780,2793|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2786,2793|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2786,2793|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2786,2793|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2786,2793|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2786,2793|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2786,2793|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2841,2845|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2841,2845|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2841,2845|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2872,2877|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2872,2877|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2872,2877|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2878,2881|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2878,2881|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2878,2881|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|2878,2881|false|false|false|||ALT
Finding|Gene or Genome|General Exam|2878,2881|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2878,2881|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2878,2881|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2878,2881|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|2885,2888|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2885,2888|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2885,2888|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2885,2888|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2885,2888|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|2885,2888|false|false|false|||AST
Finding|Gene or Genome|General Exam|2885,2888|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2892,2899|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|2892,2899|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|2916,2921|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2916,2921|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2916,2921|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2916,2929|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|2922,2929|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2922,2929|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2922,2929|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2922,2929|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2922,2929|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2922,2929|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2922,2929|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2922,2929|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|2963,2968|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2963,2968|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2963,2968|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2963,2976|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|2969,2976|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2969,2976|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2969,2976|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2969,2976|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2969,2976|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2969,2976|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2969,2976|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2969,2976|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3012,3017|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3012,3017|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3012,3017|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3012,3025|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|3018,3025|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|3018,3025|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|3018,3025|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|3018,3025|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|3018,3025|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|3018,3025|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|3018,3025|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|3031,3038|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3031,3038|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3031,3038|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3031,3038|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3031,3038|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3031,3038|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3031,3038|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3031,3038|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|General Exam|3061,3065|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|3061,3065|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|3061,3065|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|General Exam|3061,3065|false|false|false|||Iron
Procedure|Laboratory Procedure|General Exam|3061,3065|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|General Exam|3082,3087|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3082,3087|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3082,3087|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3082,3095|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3088,3095|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3088,3095|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3088,3095|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3088,3095|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3088,3095|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3088,3095|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3088,3095|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3088,3095|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3130,3135|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3130,3135|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3130,3135|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3162,3165|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|3162,3165|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|3162,3165|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|3162,3165|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|3162,3165|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|General Exam|3182,3187|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3182,3187|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3182,3187|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3212,3217|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3212,3217|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3212,3217|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3242,3247|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3242,3247|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3242,3247|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3242,3255|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|3248,3255|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|3248,3255|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|General Exam|3248,3255|false|false|false|||Lactate
Procedure|Laboratory Procedure|General Exam|3248,3255|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|General Exam|3273,3280|false|false|false|C0003962|Ascites|ASCITES
Event|Event|General Exam|3273,3280|false|false|false|||ASCITES
Finding|Pathologic Function|General Exam|3273,3280|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Drug|Amino Acid, Peptide, or Protein|General Exam|3291,3298|false|false|false|C0002712|amylase|Amylase
Drug|Enzyme|General Exam|3291,3298|false|false|false|C0002712|amylase|Amylase
Drug|Pharmacologic Substance|General Exam|3291,3298|false|false|false|C0002712|amylase|Amylase
Event|Event|General Exam|3291,3298|false|false|false|||Amylase
Procedure|Laboratory Procedure|General Exam|3291,3298|false|false|false|C0201883|Amylase measurement|Amylase
Drug|Amino Acid, Peptide, or Protein|General Exam|3314,3320|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|3314,3320|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|3314,3320|false|false|false|C0023764|lipase|Lipase
Event|Event|General Exam|3314,3320|false|false|false|||Lipase
Procedure|Laboratory Procedure|General Exam|3314,3320|false|false|false|C0373670|Lipase measurement|Lipase
Anatomy|Anatomical Structure|General Exam|3341,3345|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|BODY
Anatomy|Body Part, Organ, or Organ Component|General Exam|3341,3345|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|BODY
Finding|Intellectual Product|General Exam|3341,3345|false|false|false|C1551342|Document Body|BODY
Finding|Body Substance|General Exam|3341,3351|false|false|false|C0005889|Body Fluids|BODY FLUID
Drug|Substance|General Exam|3346,3351|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|3346,3351|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|3346,3351|false|false|false|C1546638|Fluid Specimen Code|FLUID
Disorder|Disease or Syndrome|General Exam|3375,3380|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3375,3380|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3375,3388|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|3381,3388|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3381,3388|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3381,3388|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3381,3388|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3381,3388|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|General Exam|3420,3425|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|General Exam|3420,3432|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|General Exam|3426,3432|false|false|false|C4255046||REPORT
Event|Event|General Exam|3426,3432|false|false|false|||REPORT
Finding|Intellectual Product|General Exam|3426,3432|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|General Exam|3426,3432|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|General Exam|3441,3446|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|3441,3446|false|false|false|||Blood
Finding|Body Substance|General Exam|3441,3446|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|3441,3454|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|3447,3454|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|3447,3454|false|false|false|||Culture
Finding|Functional Concept|General Exam|3447,3454|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|3447,3454|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|3447,3454|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|General Exam|3456,3463|false|false|false|||Routine
Finding|Idea or Concept|General Exam|3456,3463|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|General Exam|3456,3463|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|General Exam|3456,3463|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|General Exam|3465,3470|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Idea or Concept|General Exam|3506,3511|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Event|Event|General Exam|3512,3525|false|false|false|||SENSITIVITIES
Finding|Finding|General Exam|3512,3525|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Event|Event|General Exam|3559,3572|false|false|false|||SENSITIVITIES
Finding|Finding|General Exam|3559,3572|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|General Exam|3574,3577|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|General Exam|3574,3577|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|General Exam|3574,3577|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|General Exam|3574,3577|false|false|false|||MIC
Procedure|Laboratory Procedure|General Exam|3574,3577|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|General Exam|3574,3577|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|General Exam|3592,3595|false|false|false|||MCG
Event|Event|General Exam|3721,3727|false|false|false|||KOSERI
Drug|Antibiotic|General Exam|3762,3770|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Organic Chemical|General Exam|3762,3770|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Antibiotic|General Exam|3793,3804|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Organic Chemical|General Exam|3793,3804|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Antibiotic|General Exam|3824,3835|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|General Exam|3824,3835|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|General Exam|3855,3868|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Pharmacologic Substance|General Exam|3855,3868|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Antibiotic|General Exam|3886,3896|false|false|false|C3854019|gentamicin|GENTAMICIN
Drug|Organic Chemical|General Exam|3886,3896|false|false|false|C3854019|gentamicin|GENTAMICIN
Event|Event|General Exam|3886,3896|false|false|false|||GENTAMICIN
Procedure|Laboratory Procedure|General Exam|3886,3896|false|false|false|C0202391|Gentamicin measurement|GENTAMICIN
Drug|Antibiotic|General Exam|3917,3926|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Clinical Drug|General Exam|3917,3926|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Organic Chemical|General Exam|3917,3926|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Antibiotic|General Exam|3948,3960|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Organic Chemical|General Exam|3948,3960|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Antibiotic|General Exam|3961,3965|false|false|false|C0075870|tazobactam|TAZO
Drug|Organic Chemical|General Exam|3961,3965|false|false|false|C0075870|tazobactam|TAZO
Drug|Antibiotic|General Exam|3979,3989|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Drug|Organic Chemical|General Exam|3979,3989|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Event|Event|General Exam|3979,3989|false|false|false|||TOBRAMYCIN
Procedure|Laboratory Procedure|General Exam|3979,3989|false|false|false|C0202490|Tobramycin measurement|TOBRAMYCIN
Drug|Antibiotic|General Exam|4010,4022|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Organic Chemical|General Exam|4010,4022|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Pharmacologic Substance|General Exam|4023,4028|false|false|false|C0749139|sulfa|SULFA
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4060,4070|false|false|false|C0061856|Gram's stain|Gram Stain
Drug|Organic Chemical|General Exam|4060,4070|false|false|false|C0061856|Gram's stain|Gram Stain
Procedure|Laboratory Procedure|General Exam|4060,4070|false|false|false|C0200966|Bacterial stain, routine|Gram Stain
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4065,4070|false|false|false|C0038128|Stains|Stain
Event|Event|General Exam|4065,4070|false|false|false|||Stain
Procedure|Laboratory Procedure|General Exam|4065,4070|false|false|false|C0487602|Staining method|Stain
Finding|Idea or Concept|General Exam|4072,4077|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Classification|General Exam|4095,4103|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4095,4103|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4095,4103|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|General Exam|4104,4107|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|General Exam|4104,4107|true|false|false|C0035086|Renal Osteodystrophy|ROD
Event|Event|General Exam|4104,4107|false|false|false|||ROD
Finding|Gene or Genome|General Exam|4104,4107|true|false|false|C1424852|KNTC1 gene|ROD
Event|Event|General Exam|4119,4127|false|false|false|||Reported
Event|Event|General Exam|4135,4139|false|false|false|||read
Disorder|Disease or Syndrome|General Exam|4187,4194|false|false|false|C0000833|Abscess|ABSCESS
Event|Event|General Exam|4187,4194|false|false|false|||ABSCESS
Finding|Intellectual Product|General Exam|4187,4194|false|false|false|C1546533||ABSCESS
Anatomy|Body Part, Organ, or Organ Component|General Exam|4203,4209|false|false|false|C0030797|Pelvis|PELVIC
Disorder|Injury or Poisoning|General Exam|4210,4220|false|false|false|C1720922|Respiratory Aspiration|ASPIRATION
Event|Event|General Exam|4210,4220|false|false|false|||ASPIRATION
Finding|Finding|General Exam|4210,4220|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|ASPIRATION
Finding|Organ or Tissue Function|General Exam|4210,4220|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|ASPIRATION
Finding|Pathologic Function|General Exam|4210,4220|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|ASPIRATION
Procedure|Therapeutic or Preventive Procedure|General Exam|4210,4220|false|false|false|C0349707||ASPIRATION
Finding|Idea or Concept|General Exam|4254,4259|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|General Exam|4254,4266|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|General Exam|4260,4266|false|false|false|C4255046||REPORT
Event|Event|General Exam|4260,4266|false|false|false|||REPORT
Finding|Intellectual Product|General Exam|4260,4266|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|General Exam|4260,4266|false|false|false|C0700287|Reporting|REPORT
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4275,4285|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|4275,4285|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|4275,4285|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4280,4285|false|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|4280,4285|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|4280,4285|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|4287,4292|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4325,4330|false|false|false|||FIELD
Finding|Conceptual Entity|General Exam|4325,4330|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|4325,4330|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|General Exam|4335,4352|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|General Exam|4354,4364|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|General Exam|4354,4364|false|false|false|||LEUKOCYTES
Finding|Body Substance|General Exam|4354,4364|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|4354,4364|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Event|Event|General Exam|4393,4398|false|false|false|||FIELD
Finding|Conceptual Entity|General Exam|4393,4398|true|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|4393,4398|true|false|false|C1553496|field - patient encounter|FIELD
Finding|Classification|General Exam|4408,4416|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4408,4416|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4408,4416|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|General Exam|4417,4420|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|General Exam|4417,4420|true|false|false|C0035086|Renal Osteodystrophy|ROD
Event|Event|General Exam|4417,4420|false|false|false|||ROD
Finding|Gene or Genome|General Exam|4417,4420|true|false|false|C1424852|KNTC1 gene|ROD
Disorder|Injury or Poisoning|General Exam|4430,4435|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|General Exam|4430,4435|false|false|false|||WOUND
Finding|Body Substance|General Exam|4430,4435|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|General Exam|4430,4435|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|General Exam|4430,4435|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Laboratory Procedure|General Exam|4430,4443|false|false|false|C0855657|Wound Culture|WOUND CULTURE
Drug|Biomedical or Dental Material|General Exam|4436,4443|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4436,4443|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4436,4443|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4436,4443|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4436,4443|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4445,4450|false|false|false|||Final
Finding|Idea or Concept|General Exam|4445,4450|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4462,4468|true|false|false|||GROWTH
Finding|Finding|General Exam|4462,4468|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4462,4468|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4462,4468|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4462,4468|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4462,4468|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|General Exam|4475,4492|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|4485,4492|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4485,4492|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4485,4492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4485,4492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4485,4492|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|General Exam|4494,4499|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Disease or Syndrome|General Exam|4512,4532|false|false|false|C1456246|Bacteroides fragilis infection in conditions classified elsewhere and of unspecified site|BACTEROIDES FRAGILIS
Event|Event|General Exam|4524,4532|false|false|false|||FRAGILIS
Event|Event|General Exam|4533,4538|false|false|false|||GROUP
Finding|Body Substance|General Exam|4533,4538|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Conceptual Entity|General Exam|4533,4538|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Functional Concept|General Exam|4533,4538|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Idea or Concept|General Exam|4533,4538|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Event|Event|General Exam|4550,4556|false|false|false|||GROWTH
Finding|Finding|General Exam|4550,4556|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4550,4556|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4550,4556|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4550,4556|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4550,4556|false|false|false|C2911660|Growth action|GROWTH
Event|Event|General Exam|4568,4572|false|false|false|||BETA
Finding|Intellectual Product|General Exam|4568,4572|false|false|false|C0439096|Greek letter beta|BETA
Drug|Amino Acid, Peptide, or Protein|General Exam|4568,4582|false|false|false|C0597979|beta-Lactamase|BETA LACTAMASE
Drug|Enzyme|General Exam|4568,4582|false|false|false|C0597979|beta-Lactamase|BETA LACTAMASE
Drug|Amino Acid, Peptide, or Protein|General Exam|4573,4582|false|false|false|C2945614|lactamase|LACTAMASE
Drug|Enzyme|General Exam|4573,4582|false|false|false|C2945614|lactamase|LACTAMASE
Disorder|Cell or Molecular Dysfunction|General Exam|4583,4591|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Event|Event|General Exam|4583,4591|false|false|false|||POSITIVE
Finding|Classification|General Exam|4583,4591|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|General Exam|4583,4591|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Body Substance|General Exam|4608,4613|false|false|false|C0015733|Feces|STOOL
Finding|Finding|General Exam|4608,4629|false|false|false|C0426740|Consistency of stool|STOOL     CONSISTENCY
Event|Event|General Exam|4652,4658|true|false|false|||Source
Finding|Finding|General Exam|4652,4658|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Functional Concept|General Exam|4652,4658|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Intellectual Product|General Exam|4652,4658|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Event|Event|General Exam|4660,4665|false|false|false|||Stool
Finding|Body Substance|General Exam|4660,4665|false|false|false|C0015733|Feces|Stool
Finding|Idea or Concept|General Exam|4699,4704|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|General Exam|4699,4711|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|General Exam|4705,4711|false|false|false|C4255046||REPORT
Event|Event|General Exam|4705,4711|false|false|false|||REPORT
Finding|Intellectual Product|General Exam|4705,4711|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|General Exam|4705,4711|false|false|false|C0700287|Reporting|REPORT
Drug|Biologically Active Substance|General Exam|4733,4736|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4733,4736|false|false|false|C0012854|DNA|DNA
Finding|Genetic Function|General Exam|4733,4750|false|false|false|C0683230|dna amplification|DNA amplification
Disorder|Cell or Molecular Dysfunction|General Exam|4737,4750|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|General Exam|4737,4750|false|false|false|||amplification
Phenomenon|Phenomenon or Process|General Exam|4737,4750|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|General Exam|4737,4750|false|false|false|C1517480|Gene Amplification Technique|amplification
Event|Event|General Exam|4751,4756|false|false|false|||assay
Procedure|Laboratory Procedure|General Exam|4751,4756|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Finding|Idea or Concept|General Exam|4758,4763|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4776,4784|false|false|false|||Negative
Finding|Classification|General Exam|4776,4784|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|General Exam|4776,4784|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|General Exam|4776,4784|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|General Exam|4776,4788|false|false|false|C0205160|Negative|Negative for
Finding|Intellectual Product|General Exam|4789,4798|true|false|false|C0445332|Toxigenic|toxigenic
Drug|Biologically Active Substance|General Exam|4830,4833|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4830,4833|false|false|false|C0012854|DNA|DNA
Event|Event|General Exam|4830,4833|false|false|false|||DNA
Disorder|Cell or Molecular Dysfunction|General Exam|4840,4853|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|General Exam|4840,4853|false|false|false|||amplification
Phenomenon|Phenomenon or Process|General Exam|4840,4853|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|General Exam|4840,4853|false|false|false|C1517480|Gene Amplification Technique|amplification
Event|Event|General Exam|4854,4859|false|false|false|||assay
Procedure|Laboratory Procedure|General Exam|4854,4859|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Finding|Conceptual Entity|General Exam|4874,4883|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Idea or Concept|General Exam|4874,4883|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|General Exam|4874,4883|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|General Exam|4884,4889|false|false|false|C3542016|Concept model range (foundation metadata concept)|Range
Event|Event|General Exam|4890,4898|false|false|false|||Negative
Finding|Classification|General Exam|4890,4898|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|General Exam|4890,4898|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|General Exam|4890,4898|false|false|false|C5237010|Expression Negative|Negative
Event|Event|Hospital Course|4940,4948|false|false|false|||admitted
Event|Occupational Activity|Hospital Course|4960,4967|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|4960,4967|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|4973,4983|false|false|false|||management
Event|Occupational Activity|Hospital Course|4973,4983|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|4973,4983|false|false|false|C0376636|Disease Management|management
Disorder|Disease or Syndrome|Hospital Course|4987,4992|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|Hospital Course|4987,4992|false|false|false|||ileus
Event|Event|Hospital Course|5000,5009|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5000,5009|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Location or Region|Hospital Course|5013,5024|false|false|false|C3282907|Nasogastric|nasogastric
Finding|Functional Concept|Hospital Course|5013,5024|false|false|false|C0694637|Nasogastric Route of Administration|nasogastric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5013,5029|false|false|false|C0812428|Nasogastric tube procedures|nasogastric tube
Event|Event|Hospital Course|5025,5029|false|false|false|||tube
Finding|Functional Concept|Hospital Course|5025,5029|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Hospital Course|5025,5029|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|Hospital Course|5035,5041|false|false|false|||placed
Event|Event|Hospital Course|5046,5059|false|false|false|||decompression
Finding|Functional Concept|Hospital Course|5046,5059|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|Hospital Course|5046,5059|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5046,5059|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Event|Event|Hospital Course|5070,5074|false|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5070,5074|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Event|Event|Hospital Course|5079,5085|false|false|false|||placed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5090,5093|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Biologically Active Substance|Hospital Course|5090,5093|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|5090,5093|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Event|Event|Hospital Course|5090,5093|false|false|false|||TPN
Finding|Gene or Genome|Hospital Course|5090,5093|false|false|false|C1420583;C3813711|TAPBP gene;TAPBP wt Allele|TPN
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5090,5093|false|false|false|C0030548|Parenteral Nutrition, Total|TPN
Event|Event|Hospital Course|5095,5102|false|false|false|||started
Disorder|Disease or Syndrome|Hospital Course|5105,5110|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|Hospital Course|5105,5110|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|Hospital Course|5105,5119|true|false|false|C0200949|Blood culture|Blood cultures
Event|Event|Hospital Course|5111,5119|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|5111,5119|false|false|false|C0010453|Culture (Anthropological)|cultures
Finding|Classification|Hospital Course|5130,5138|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5130,5138|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5130,5138|false|false|false|C5237010|Expression Negative|negative
Anatomy|Cell|Hospital Course|5139,5143|false|false|false|C0206427|Rod Photoreceptors|rods
Drug|Antibiotic|Hospital Course|5148,5159|true|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|5148,5159|true|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|5148,5159|false|false|false|||ceftriaxone
Event|Event|Hospital Course|5165,5172|false|false|false|||started
Event|Event|Hospital Course|5186,5193|false|false|false|||started
Event|Event|Hospital Course|5197,5201|false|false|false|||pass
Event|Event|Hospital Course|5208,5214|false|false|false|||amount
Finding|Intellectual Product|Hospital Course|5208,5214|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|Hospital Course|5219,5225|false|false|false|||flatus
Finding|Sign or Symptom|Hospital Course|5219,5225|false|false|false|C0016204|Flatulence|flatus
Procedure|Diagnostic Procedure|Hospital Course|5232,5239|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|5235,5239|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|5235,5239|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|5240,5252|false|false|false|||demonstrated
Disorder|Disease or Syndrome|Hospital Course|5263,5268|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|Hospital Course|5263,5268|false|false|false|||ileus
Event|Event|Hospital Course|5274,5281|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|5274,5281|false|false|false|C2699424|Concern|concern
Finding|Finding|Hospital Course|5287,5295|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|5296,5301|false|false|false|||urine
Finding|Body Substance|Hospital Course|5296,5301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|5296,5301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|5296,5301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Pathologic Function|Hospital Course|5296,5306|false|true|false|C0042024|Urinary Incontinence|urine leak
Event|Event|Hospital Course|5302,5306|false|false|false|||leak
Finding|Functional Concept|Hospital Course|5302,5306|false|true|false|C0332234|Leaking|leak
Event|Event|Hospital Course|5311,5320|false|false|false|||increased
Finding|Functional Concept|Hospital Course|5321,5325|false|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|Hospital Course|5321,5331|false|false|false|C0013687|effusion|free fluid
Drug|Substance|Hospital Course|5326,5331|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Hospital Course|5326,5331|false|false|false|||fluid
Finding|Intellectual Product|Hospital Course|5326,5331|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Hospital Course|5345,5348|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|Hospital Course|5349,5354|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|Hospital Course|5349,5354|false|false|false|||drain
Finding|Intellectual Product|Hospital Course|5349,5354|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|Hospital Course|5359,5365|false|false|false|||placed
Procedure|Diagnostic Procedure|Hospital Course|5369,5383|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|interventional
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5369,5383|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|interventional
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5369,5393|false|false|false|C0344093|Interventional Radiology Procedure|interventional radiology
Event|Event|Hospital Course|5384,5393|false|false|false|||radiology
Finding|Finding|Hospital Course|5384,5393|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Finding|Idea or Concept|Hospital Course|5384,5393|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Finding|Intellectual Product|Hospital Course|5384,5393|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|radiology
Procedure|Diagnostic Procedure|Hospital Course|5384,5393|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|radiology
Event|Event|Hospital Course|5408,5414|false|false|false|||passed
Finding|Functional Concept|Hospital Course|5415,5420|false|false|false|C1418448;C1423795;C1883710;C3810601|Clamping Activity;PDZK1 gene;PDZK1 wt Allele;SPEF1 gene|clamp
Finding|Gene or Genome|Hospital Course|5415,5420|false|false|false|C1418448;C1423795;C1883710;C3810601|Clamping Activity;PDZK1 gene;PDZK1 wt Allele;SPEF1 gene|clamp
Event|Event|Hospital Course|5421,5426|false|false|false|||trial
Procedure|Research Activity|Hospital Course|5421,5426|false|false|false|C0008976|Clinical Trials|trial
Event|Event|Hospital Course|5431,5434|false|false|false|||NGT
Event|Event|Hospital Course|5439,5446|false|false|false|||removed
Event|Event|Hospital Course|5452,5461|false|false|false|||continued
Event|Event|Hospital Course|5465,5469|false|false|false|||pass
Finding|Finding|Hospital Course|5465,5469|false|false|false|C2828386|Pass (indicator)|pass
Event|Event|Hospital Course|5471,5477|false|false|false|||flatus
Finding|Sign or Symptom|Hospital Course|5471,5477|false|false|false|C0016204|Flatulence|flatus
Event|Event|Hospital Course|5487,5494|false|false|false|||started
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5503,5508|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Hospital Course|5503,5518|false|false|false|C0011135|Defecation|bowel movements
Event|Event|Hospital Course|5509,5518|false|false|false|||movements
Finding|Organism Function|Hospital Course|5509,5518|false|false|false|C0026649|Movement|movements
Event|Event|Hospital Course|5537,5545|false|false|false|||advanced
Finding|Idea or Concept|Hospital Course|5551,5556|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|Hospital Course|5551,5563|false|false|false|C4264429|Clear liquid|clear liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5551,5568|false|false|false|C2184084|Clear liquid diet|clear liquid diet
Drug|Biomedical or Dental Material|Hospital Course|5557,5563|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|Hospital Course|5557,5563|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Event|Event|Hospital Course|5557,5563|false|false|false|||liquid
Finding|Finding|Hospital Course|5557,5563|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5557,5563|false|false|false|C0301571|Liquid diet|liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5557,5568|false|false|false|C0301571|Liquid diet|liquid diet
Drug|Food|Hospital Course|5564,5568|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|5564,5568|false|false|false|||diet
Finding|Functional Concept|Hospital Course|5564,5568|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5564,5568|false|false|false|C0012159|Diet therapy|diet
Finding|Functional Concept|Hospital Course|5571,5577|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Disorder|Disease or Syndrome|Hospital Course|5578,5583|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|5578,5583|false|false|false|||blood
Finding|Body Substance|Hospital Course|5578,5583|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Hospital Course|5578,5592|false|true|false|C0200949|Blood culture|blood cultures
Event|Event|Hospital Course|5584,5592|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|5584,5592|false|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|Hospital Course|5599,5607|false|false|false|||negative
Finding|Classification|Hospital Course|5599,5607|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5599,5607|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5599,5607|false|false|false|C5237010|Expression Negative|negative
Disorder|Cell or Molecular Dysfunction|Hospital Course|5612,5620|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|5612,5620|false|false|false|||positive
Finding|Classification|Hospital Course|5612,5620|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|5612,5620|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Lab|Laboratory or Test Result|Hospital Course|5612,5634|false|false|false|C0740299|Organism isolated in blood by culture|positive blood culture
Disorder|Disease or Syndrome|Hospital Course|5621,5626|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|5621,5626|false|false|false|||blood
Finding|Body Substance|Hospital Course|5621,5626|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Hospital Course|5621,5634|false|false|false|C0200949|Blood culture|blood culture
Drug|Biomedical or Dental Material|Hospital Course|5627,5634|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|5627,5634|false|false|false|||culture
Finding|Functional Concept|Hospital Course|5627,5634|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|5627,5634|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|5627,5634|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|Hospital Course|5640,5649|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5640,5649|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|5656,5667|false|false|false|||citrobacter
Drug|Food|Hospital Course|5670,5674|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Event|Event|Hospital Course|5670,5674|false|false|false|||Diet
Finding|Functional Concept|Hospital Course|5670,5674|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|Hospital Course|5670,5674|false|false|false|C0012159|Diet therapy|Diet
Event|Event|Hospital Course|5689,5697|false|false|false|||advanced
Event|Event|Hospital Course|5702,5708|false|false|false|||ensure
Event|Event|Hospital Course|5709,5714|false|false|false|||added
Attribute|Clinical Attribute|Hospital Course|5720,5731|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5720,5731|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|5720,5731|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|5720,5731|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|5747,5756|false|false|false|||converted
Event|Event|Hospital Course|5776,5788|false|false|false|||re-evaluated
Finding|Finding|Hospital Course|5792,5800|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|5792,5800|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|5792,5800|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Hospital Course|5792,5808|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5792,5808|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Hospital Course|5801,5808|false|false|false|||therapy
Finding|Finding|Hospital Course|5801,5808|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|5801,5808|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5801,5808|false|false|false|C0087111|Therapeutic procedure|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5813,5827|false|false|false|C0034991|Rehabilitation therapy|rehabilitative
Finding|Intellectual Product|Hospital Course|5813,5836|false|false|false|C4523774|Rehabilitative Services|rehabilitative services
Event|Event|Hospital Course|5828,5836|false|false|false|||services
Event|Occupational Activity|Hospital Course|5828,5836|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|5828,5836|false|false|false|C1704289|Clinical Service|services
Event|Event|Hospital Course|5847,5857|false|false|false|||ambulating
Event|Event|Hospital Course|5870,5880|false|false|false|||assistance
Finding|Social Behavior|Hospital Course|5870,5880|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|Hospital Course|5885,5893|false|false|false|||prepared
Event|Event|Hospital Course|5899,5908|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5899,5908|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5899,5908|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5899,5908|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5899,5908|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|5920,5928|false|false|false|||facility
Finding|Intellectual Product|Hospital Course|5920,5928|false|false|false|C4695111|ADMIN.FACILITY|facility
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5936,5939|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Biologically Active Substance|Hospital Course|5936,5939|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|5936,5939|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Event|Event|Hospital Course|5936,5939|false|false|false|||TPN
Finding|Gene or Genome|Hospital Course|5936,5939|false|false|false|C1420583;C3813711|TAPBP gene;TAPBP wt Allele|TPN
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5936,5939|false|false|false|C0030548|Parenteral Nutrition, Total|TPN
Event|Event|Hospital Course|5945,5954|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|5964,5967|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5964,5967|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5975,5984|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5975,5984|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5975,5984|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5975,5984|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5975,5984|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|5989,5993|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|5989,5993|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|5989,5993|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|5997,6006|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5997,6006|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5997,6006|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5997,6006|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5997,6006|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6017,6027|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|6028,6040|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|6036,6040|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|6036,6040|false|false|false|||diet
Finding|Functional Concept|Hospital Course|6036,6040|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|6036,6040|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|6042,6049|false|false|false|||passing
Attribute|Clinical Attribute|Hospital Course|6042,6056|false|false|false|C4050437||passing flatus
Finding|Sign or Symptom|Hospital Course|6042,6056|false|false|false|C0016204|Flatulence|passing flatus
Event|Event|Hospital Course|6050,6056|false|false|false|||flatus
Finding|Sign or Symptom|Hospital Course|6050,6056|false|false|false|C0016204|Flatulence|flatus
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6079,6084|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Hospital Course|6079,6094|false|false|false|C0011135|Defecation|bowel movements
Event|Event|Hospital Course|6085,6094|false|false|false|||movements
Finding|Organism Function|Hospital Course|6085,6094|false|false|false|C0026649|Movement|movements
Attribute|Clinical Attribute|Hospital Course|6099,6110|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6099,6110|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6099,6110|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6099,6110|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|6099,6123|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|6114,6123|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|6114,6123|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|6142,6152|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|6142,6152|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|6142,6157|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|6153,6157|false|false|false|||list
Finding|Intellectual Product|Hospital Course|6153,6157|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|6161,6169|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|6174,6182|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|6174,6182|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|6174,6182|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|6174,6182|false|false|false|||complete
Finding|Functional Concept|Hospital Course|6174,6182|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6174,6182|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|6187,6199|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6187,6199|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6217,6230|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|6217,6230|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|6217,6230|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|6217,6230|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6217,6237|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|6217,6237|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|6217,6237|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|6231,6237|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6231,6237|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6231,6237|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6231,6237|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6231,6237|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6231,6237|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|6259,6267|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Hospital Course|6259,6267|false|false|false|C0126174|losartan|Losartan
Event|Event|Hospital Course|6259,6267|false|false|false|||Losartan
Drug|Organic Chemical|Hospital Course|6259,6277|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Hospital Course|6259,6277|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Hospital Course|6268,6277|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|6268,6277|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|6268,6277|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|6268,6277|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|6268,6277|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|6268,6277|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|6268,6277|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|6268,6277|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Hospital Course|6297,6310|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6297,6310|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|6297,6310|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6297,6310|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|6329,6337|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|6329,6337|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|6329,6337|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|6329,6344|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|6329,6344|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|6338,6344|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6338,6344|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6338,6344|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6338,6344|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6338,6344|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6338,6344|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6355,6358|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6355,6358|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6355,6358|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6355,6358|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6355,6358|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6363,6373|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|6363,6373|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|6363,6373|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|6363,6380|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|6363,6380|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|6374,6380|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6374,6380|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6374,6380|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6374,6380|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6374,6380|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6374,6380|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|6400,6414|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Pharmacologic Substance|Hospital Course|6400,6414|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Organic Chemical|Hospital Course|6424,6432|false|false|false|C0591750|Macrobid|MacroBID
Drug|Pharmacologic Substance|Hospital Course|6424,6432|false|false|false|C0591750|Macrobid|MacroBID
Drug|Organic Chemical|Hospital Course|6454,6463|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|Hospital Course|6454,6463|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|Hospital Course|6454,6463|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|Hospital Course|6454,6463|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|Hospital Course|6465,6474|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|6465,6474|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|6465,6482|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|6475,6482|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6475,6482|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6475,6482|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6475,6482|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|6496,6499|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|6500,6504|false|false|false|C2598155||Pain
Event|Event|Hospital Course|6500,6504|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|6500,6504|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|6500,6504|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|6507,6515|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|6507,6515|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|6521,6530|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6521,6530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6521,6530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6521,6530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6521,6530|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6521,6542|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6531,6542|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6531,6542|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6531,6542|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6531,6542|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6548,6561|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|Hospital Course|6548,6561|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Antibiotic|Hospital Course|6548,6565|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Drug|Organic Chemical|Hospital Course|6548,6565|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Disorder|Neoplastic Process|Hospital Course|6562,6565|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|6562,6565|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|6562,6565|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|6562,6565|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|6562,6565|false|false|false|||HCl
Drug|Pharmacologic Substance|Hospital Course|6581,6589|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|6581,6589|false|false|false|||Duration
Drug|Organic Chemical|Hospital Course|6619,6632|false|false|false|C0025872|metronidazole|MetroNIDAZOLE
Drug|Pharmacologic Substance|Hospital Course|6619,6632|false|false|false|C0025872|metronidazole|MetroNIDAZOLE
Drug|Pharmacologic Substance|Hospital Course|6647,6655|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|6647,6655|false|false|false|||Duration
Drug|Organic Chemical|Hospital Course|6685,6690|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|6685,6690|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6701,6704|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6701,6704|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6701,6704|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6701,6704|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6701,6704|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6711,6724|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6711,6724|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|6711,6724|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6711,6724|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|6745,6757|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6745,6757|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|6777,6785|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|6777,6785|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|6777,6785|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|6777,6792|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|6777,6792|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|6786,6792|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6786,6792|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6786,6792|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6786,6792|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6786,6792|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6786,6792|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6803,6806|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6803,6806|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6803,6806|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6803,6806|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6803,6806|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6813,6823|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|6813,6823|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|6813,6823|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|6813,6830|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|6813,6830|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|6824,6830|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6824,6830|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6824,6830|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6824,6830|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6824,6830|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6824,6830|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|6847,6852|false|false|false|||Start
Finding|Idea or Concept|Hospital Course|6871,6875|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|Hospital Course|6876,6883|false|false|false|||Routine
Finding|Idea or Concept|Hospital Course|6876,6883|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|6876,6883|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|6876,6883|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|6884,6898|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6884,6898|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|6899,6903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|6899,6903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|6899,6903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6910,6923|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|6910,6923|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|6910,6923|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|6910,6923|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6910,6930|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|6910,6930|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|6910,6930|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|6924,6930|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6924,6930|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6924,6930|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6924,6930|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6924,6930|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6924,6930|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|6954,6963|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|Hospital Course|6954,6963|false|false|false|C0024002|lorazepam|LORazepam
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6975,6978|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6975,6978|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6975,6978|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6975,6978|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6975,6978|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|6979,6982|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6983,6990|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|6983,6990|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|6983,6990|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|Hospital Course|6998,7006|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Hospital Course|6998,7006|false|false|false|C0126174|losartan|Losartan
Event|Event|Hospital Course|6998,7006|false|false|false|||Losartan
Drug|Organic Chemical|Hospital Course|6998,7016|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Hospital Course|6998,7016|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Hospital Course|7007,7016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|7007,7016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|7007,7016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|7007,7016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|7007,7016|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|7007,7016|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|7007,7016|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|7007,7016|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Hospital Course|7039,7053|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Pharmacologic Substance|Hospital Course|7039,7053|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Organic Chemical|Hospital Course|7063,7071|false|false|false|C0591750|Macrobid|MacroBID
Drug|Pharmacologic Substance|Hospital Course|7063,7071|false|false|false|C0591750|Macrobid|MacroBID
Drug|Organic Chemical|Hospital Course|7096,7105|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|Hospital Course|7096,7105|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|Hospital Course|7096,7105|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|Hospital Course|7096,7105|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|Hospital Course|7107,7116|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|7107,7116|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|7107,7124|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|7117,7124|false|false|false|||Release
Finding|Functional Concept|Hospital Course|7117,7124|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7117,7124|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7117,7124|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|7138,7141|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|7142,7146|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|7142,7146|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|7142,7146|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|7150,7158|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|7150,7158|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|7164,7173|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|7164,7173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7164,7173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7164,7173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7164,7173|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|7164,7185|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|7164,7185|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|7174,7185|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|7174,7185|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|7174,7185|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|7187,7195|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7187,7195|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|7187,7200|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|7196,7200|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|7196,7200|false|false|false|||Care
Finding|Finding|Hospital Course|7196,7200|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|7196,7200|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|7203,7211|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|7203,7211|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|7219,7228|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7219,7228|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7219,7228|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|7219,7238|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|7229,7238|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|7229,7238|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|7229,7238|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|7229,7238|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|7229,7238|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7240,7247|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|7240,7247|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7240,7247|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Hospital Course|7240,7254|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|Hospital Course|7248,7254|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|7248,7254|false|false|false|||cancer
Disorder|Disease or Syndrome|Hospital Course|7271,7276|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|Hospital Course|7271,7276|false|false|false|||ileus
Event|Event|Hospital Course|7278,7288|false|false|false|||bacteremia
Finding|Finding|Hospital Course|7278,7288|false|false|false|C0004610|Bacteremia|bacteremia
Anatomy|Body Location or Region|Hospital Course|7315,7324|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7325,7331|false|false|false|C0030797|Pelvis|pelvic
Disorder|Disease or Syndrome|Hospital Course|7325,7339|false|false|false|C0030785|Pelvic abscess|pelvic abscess
Disorder|Disease or Syndrome|Hospital Course|7332,7339|false|false|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|7332,7339|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|7332,7339|false|false|false|C1546533||abscess
Disorder|Disease or Syndrome|Hospital Course|7341,7361|false|false|false|C1456246|Bacteroides fragilis infection in conditions classified elsewhere and of unspecified site|BACTEROIDES FRAGILIS
Event|Event|Hospital Course|7353,7361|false|false|false|||FRAGILIS
Finding|Body Substance|Hospital Course|7363,7368|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Conceptual Entity|Hospital Course|7363,7368|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Functional Concept|Hospital Course|7363,7368|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Finding|Idea or Concept|Hospital Course|7363,7368|false|false|false|C0441833;C1519504;C1561557;C1705428|Group Object;Group Specimen;Groups;Stage Grouping|GROUP
Event|Event|Hospital Course|7370,7379|false|false|false|||requiring
Event|Event|Hospital Course|7384,7392|false|false|false|||drainage
Finding|Body Substance|Hospital Course|7384,7392|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Hospital Course|7384,7392|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7384,7392|false|false|false|C0013103|Drainage procedure|drainage
Finding|Mental Process|Discharge Condition|7417,7423|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|7417,7430|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|7417,7430|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|7424,7430|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|7424,7430|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7432,7437|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|7432,7437|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|7442,7450|false|false|false|||coherent
Finding|Finding|Discharge Condition|7442,7450|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|7452,7457|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|7452,7474|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|7452,7474|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|7461,7474|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|7461,7474|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|7461,7474|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|7476,7481|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|7476,7481|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|7476,7481|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|7476,7481|false|false|false|||Alert
Finding|Finding|Discharge Condition|7476,7481|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|7476,7481|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|7476,7481|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|7486,7497|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|7486,7497|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|7499,7507|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|7499,7507|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|7499,7507|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|7508,7514|false|false|false|C5889824||Status
Event|Event|Discharge Condition|7508,7514|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|7508,7514|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|7516,7526|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|7516,7526|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|7516,7526|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|7516,7526|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|7529,7537|false|false|false|||requires
Event|Event|Discharge Condition|7538,7548|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|7538,7548|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|7552,7555|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|7552,7555|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|7552,7555|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|7552,7555|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|7552,7555|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|7557,7563|false|false|false|||walker
Event|Event|Discharge Instructions|7615,7620|false|false|false|||refer
Attribute|Clinical Attribute|Discharge Instructions|7628,7640|false|false|false|C3263700||instructions
Event|Event|Discharge Instructions|7628,7640|false|false|false|||instructions
Finding|Intellectual Product|Discharge Instructions|7628,7640|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Attribute|Clinical Attribute|Discharge Instructions|7628,7649|false|false|false|C4554379||instructions provided
Finding|Finding|Discharge Instructions|7628,7649|false|false|false|C4554380|Instructions provided|instructions provided
Event|Event|Discharge Instructions|7641,7649|false|false|false|||provided
Event|Event|Discharge Instructions|7665,7671|false|false|false|||Ostomy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7665,7671|false|false|false|C0029473|Ostomy|Ostomy
Event|Event|Discharge Instructions|7678,7688|false|false|false|||specialist
Finding|Classification|Discharge Instructions|7678,7688|false|false|false|C4521398|United States Military enlisted E4 (qualifier value)|specialist
Event|Event|Discharge Instructions|7694,7701|false|false|false|||details
Finding|Functional Concept|Discharge Instructions|7706,7714|false|false|false|C1514873;C1546857;C1556066;C1619636;C3245501;C3245502|Required - Escort Required;Requirement;required - CodingRationale;required - HL7ConformanceInclusion;required - HL7V3Conformance;required - ParticipationSignature|required
Finding|Idea or Concept|Discharge Instructions|7706,7714|false|false|false|C1514873;C1546857;C1556066;C1619636;C3245501;C3245502|Required - Escort Required;Requirement;required - CodingRationale;required - HL7ConformanceInclusion;required - HL7V3Conformance;required - ParticipationSignature|required
Finding|Intellectual Product|Discharge Instructions|7706,7714|false|false|false|C1514873;C1546857;C1556066;C1619636;C3245501;C3245502|Required - Escort Required;Requirement;required - CodingRationale;required - HL7ConformanceInclusion;required - HL7V3Conformance;required - ParticipationSignature|required
Event|Activity|Discharge Instructions|7715,7719|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|7715,7719|false|false|false|||care
Finding|Finding|Discharge Instructions|7715,7719|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|7715,7719|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|7725,7735|false|false|false|||management
Event|Occupational Activity|Discharge Instructions|7725,7735|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Discharge Instructions|7725,7735|false|false|false|C0376636|Disease Management|management
Anatomy|Anatomical Structure|Discharge Instructions|7744,7752|false|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7744,7752|false|false|false|C0856443|Urostomy procedure|Urostomy
Event|Event|Discharge Instructions|7755,7761|false|false|false|||Resume
Finding|Functional Concept|Discharge Instructions|7755,7761|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Idea or Concept|Discharge Instructions|7755,7761|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Intellectual Product|Discharge Instructions|7755,7761|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Conceptual Entity|Discharge Instructions|7767,7780|false|false|false|C4724283|Pre-admission Encounter|pre-admission
Finding|Idea or Concept|Discharge Instructions|7781,7785|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|7781,7785|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|7781,7785|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|7786,7797|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7786,7797|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|7786,7797|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|7786,7797|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|7808,7813|false|false|false|||noted
Finding|Finding|Discharge Instructions|7816,7822|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|Always
Finding|Idea or Concept|Discharge Instructions|7816,7822|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|Always
Event|Event|Discharge Instructions|7823,7827|true|false|false|||call
Finding|Functional Concept|Discharge Instructions|7823,7827|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Discharge Instructions|7823,7827|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Discharge Instructions|7823,7827|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Discharge Instructions|7823,7827|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Event|Event|Discharge Instructions|7831,7837|true|false|false|||inform
Event|Occupational Activity|Discharge Instructions|7831,7837|true|false|false|C1552002|inform|inform
Procedure|Health Care Activity|Discharge Instructions|7831,7837|true|false|false|C0700287|Reporting|inform
Event|Event|Discharge Instructions|7839,7845|true|false|false|||review
Finding|Idea or Concept|Discharge Instructions|7839,7845|true|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|Discharge Instructions|7839,7845|true|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Event|Event|Discharge Instructions|7850,7857|true|false|false|||discuss
Drug|Pharmacologic Substance|Discharge Instructions|7862,7872|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|7862,7872|true|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|7862,7872|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|7873,7880|true|false|false|||changes
Finding|Functional Concept|Discharge Instructions|7873,7880|true|false|true|C0392747|Changing|changes
Event|Event|Discharge Instructions|7906,7912|true|false|false|||course
Finding|Intellectual Product|Discharge Instructions|7923,7935|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|7923,7935|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Discharge Instructions|7931,7935|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|7931,7935|false|false|false|||care
Finding|Finding|Discharge Instructions|7931,7935|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|7931,7935|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|7936,7942|false|false|false|C2348314|Doctor - Title|doctor
Drug|Organic Chemical|Discharge Instructions|7950,7963|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Discharge Instructions|7950,7963|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Discharge Instructions|7950,7963|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Discharge Instructions|7950,7963|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Organic Chemical|Discharge Instructions|7969,7978|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|7969,7978|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Discharge Instructions|7969,7978|false|false|false|||Ibuprofen
Attribute|Clinical Attribute|Discharge Instructions|7983,7987|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7983,7987|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7983,7987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7983,7987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|7983,7995|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7983,7995|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Discharge Instructions|7988,7995|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|7988,7995|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|7988,7995|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Discharge Instructions|7988,7995|false|false|false|||control
Finding|Conceptual Entity|Discharge Instructions|7988,7995|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|7988,7995|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|7988,7995|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|Discharge Instructions|7999,8012|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|Discharge Instructions|7999,8012|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|Discharge Instructions|7999,8030|false|false|false|C3871468|ciprofloxacin and metronidazole|Ciprofloxacin and Metronidazole
Drug|Organic Chemical|Discharge Instructions|8017,8030|false|false|false|C0025872|metronidazole|Metronidazole
Drug|Pharmacologic Substance|Discharge Instructions|8017,8030|false|false|false|C0025872|metronidazole|Metronidazole
Event|Event|Discharge Instructions|8017,8030|false|false|false|||Metronidazole
Finding|Finding|Discharge Instructions|8035,8038|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|8035,8038|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Antibiotic|Discharge Instructions|8039,8049|false|false|false|C0003232|Antibiotics|ANTIBIOTIC
Attribute|Clinical Attribute|Discharge Instructions|8050,8061|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|8050,8061|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|8050,8061|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|8050,8061|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|8066,8071|false|false|false|||treat
Disorder|Disease or Syndrome|Discharge Instructions|8077,8086|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|8077,8086|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|8077,8086|false|false|false|C3714514|Infection|infection
Event|Event|Discharge Instructions|8088,8096|false|false|false|||Continue
Event|Event|Discharge Instructions|8135,8139|false|false|false|||dose
Drug|Organic Chemical|Discharge Instructions|8143,8150|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|8143,8150|false|false|false|C0699142|Tylenol|Tylenol
Drug|Organic Chemical|Discharge Instructions|8152,8165|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|ACETAMINOPHEN
Drug|Pharmacologic Substance|Discharge Instructions|8152,8165|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|ACETAMINOPHEN
Event|Event|Discharge Instructions|8152,8165|false|false|false|||ACETAMINOPHEN
Procedure|Laboratory Procedure|Discharge Instructions|8152,8165|false|false|false|C0373527|Acetaminophen measurement|ACETAMINOPHEN
Event|Event|Discharge Instructions|8172,8177|false|false|false|||grams
Event|Event|Discharge Instructions|8189,8196|false|false|false|||sources
Finding|Finding|Discharge Instructions|8189,8196|false|false|false|C0449416|Source|sources
Event|Event|Discharge Instructions|8202,8205|false|false|false|||DAY
Finding|Idea or Concept|Discharge Instructions|8202,8205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Discharge Instructions|8202,8205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Event|Event|Discharge Instructions|8220,8226|false|false|false|||taking
Drug|Organic Chemical|Discharge Instructions|8227,8236|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|8227,8236|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Discharge Instructions|8227,8236|false|false|false|||Ibuprofen
Finding|Intellectual Product|Discharge Instructions|8238,8249|false|false|false|C0592503|Proprietary Name|Brand names
Event|Event|Discharge Instructions|8244,8249|false|false|false|||names
Finding|Intellectual Product|Discharge Instructions|8244,8249|false|false|false|C0027365|Name|names
Finding|Finding|Discharge Instructions|8275,8281|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|Discharge Instructions|8275,8281|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Event|Event|Discharge Instructions|8285,8290|false|false|false|||taken
Drug|Food|Discharge Instructions|8296,8300|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|Discharge Instructions|8296,8300|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|Discharge Instructions|8296,8300|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|Discharge Instructions|8296,8300|false|false|false|||food
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8317,8324|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Discharge Instructions|8317,8324|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Discharge Instructions|8317,8324|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Discharge Instructions|8317,8324|false|false|false|||stomach
Finding|Finding|Discharge Instructions|8317,8324|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8317,8324|false|false|false|C0872393|Procedure on stomach|stomach
Attribute|Clinical Attribute|Discharge Instructions|8326,8330|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|8326,8330|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|8326,8330|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8326,8330|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|8334,8338|false|false|false|||note
Finding|Pathologic Function|Discharge Instructions|8339,8350|false|false|false|C0025222;C0474585|Melena|black stool
Finding|Sign or Symptom|Discharge Instructions|8339,8350|false|false|false|C0025222;C0474585|Melena|black stool
Event|Event|Discharge Instructions|8345,8350|false|false|false|||stool
Finding|Body Substance|Discharge Instructions|8345,8350|false|false|false|C0015733|Feces|stool
Event|Event|Discharge Instructions|8352,8356|false|false|false|||stop
Drug|Organic Chemical|Discharge Instructions|8361,8370|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|8361,8370|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Discharge Instructions|8361,8370|false|false|false|||Ibuprofen
Event|Event|Discharge Instructions|8388,8393|true|false|false|||drive
Event|Event|Discharge Instructions|8395,8402|true|false|false|||operate
Disorder|Injury or Poisoning|Discharge Instructions|8413,8422|true|false|false|C0337246|Contact with machinery|machinery
Event|Event|Discharge Instructions|8413,8422|true|false|false|||machinery
Event|Event|Discharge Instructions|8427,8434|false|false|false|||consume
Drug|Organic Chemical|Discharge Instructions|8436,8443|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|8436,8443|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Discharge Instructions|8436,8443|false|false|false|||alcohol
Finding|Intellectual Product|Discharge Instructions|8436,8443|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|Discharge Instructions|8450,8456|false|false|false|||taking
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8457,8465|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|8457,8465|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|8466,8470|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|8466,8470|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|8466,8470|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8466,8470|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|8471,8482|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|8471,8482|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|8471,8482|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|8471,8482|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|8493,8498|true|false|false|||drive
Event|Event|Discharge Instructions|8517,8524|true|false|false|||cleared
Event|Event|Discharge Instructions|8528,8534|false|false|false|||resume
Event|Activity|Discharge Instructions|8541,8551|false|false|false|C0441655|Activities|activities
Event|Event|Discharge Instructions|8541,8551|false|false|false|||activities
Finding|Finding|Discharge Instructions|8541,8551|false|false|false|C2239122|activities (history)|activities
Disorder|Disease or Syndrome|Discharge Instructions|8560,8563|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|8560,8563|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|8560,8563|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|8560,8563|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|8560,8563|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8560,8563|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|8560,8563|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|8560,8563|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Discharge Instructions|8560,8563|false|false|false|||PCP
Finding|Gene or Genome|Discharge Instructions|8560,8563|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|8560,8563|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Discharge Instructions|8567,8576|false|false|false|||urologist
Event|Event|Discharge Instructions|8591,8600|false|false|false|||passenger
Drug|Organic Chemical|Discharge Instructions|8603,8609|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|8603,8609|false|false|false|C0282139|Colace|Colace
Event|Event|Discharge Instructions|8624,8634|false|false|false|||prescribed
Event|Event|Discharge Instructions|8638,8643|false|false|false|||avoid
Event|Event|Discharge Instructions|8649,8657|false|false|false|||surgical
Procedure|Health Care Activity|Discharge Instructions|8649,8657|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8649,8657|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|Discharge Instructions|8659,8671|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|8659,8671|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|8676,8688|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|8676,8688|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Discharge Instructions|8689,8696|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Discharge Instructions|8689,8696|false|false|false|||related
Finding|Finding|Discharge Instructions|8689,8696|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Discharge Instructions|8689,8696|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8700,8708|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|8700,8708|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|8709,8713|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|8709,8713|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|8709,8713|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8709,8713|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|8715,8725|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|8715,8725|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|8715,8725|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|8727,8738|false|false|false|||Discontinue
Finding|Sign or Symptom|Discharge Instructions|8742,8753|false|false|false|C2129214|Loose stool|loose stool
Event|Event|Discharge Instructions|8748,8753|false|false|false|||stool
Finding|Body Substance|Discharge Instructions|8748,8753|false|false|false|C0015733|Feces|stool
Event|Event|Discharge Instructions|8757,8765|false|false|false|||diarrhea
Finding|Finding|Discharge Instructions|8757,8765|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|8757,8765|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|Discharge Instructions|8766,8774|false|false|false|||develops
Drug|Organic Chemical|Discharge Instructions|8777,8783|true|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|8777,8783|true|false|false|C0282139|Colace|Colace
Event|Event|Discharge Instructions|8777,8783|true|false|false|||Colace
Finding|Body Substance|Discharge Instructions|8789,8794|true|false|false|C0015733|Feces|stool
Event|Event|Discharge Instructions|8795,8803|true|false|false|||softener
Drug|Pharmacologic Substance|Discharge Instructions|8811,8819|true|false|false|C0282090|Laxatives|laxative
Event|Event|Discharge Instructions|8811,8819|true|false|false|||laxative
Event|Activity|Discharge Instructions|8832,8839|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|8832,8839|true|false|false|||lifting
Finding|Finding|Discharge Instructions|8866,8875|true|false|false|C3845310|10 pounds|10 pounds
Event|Event|Discharge Instructions|8878,8880|true|false|false|||Do
Event|Event|Discharge Instructions|8891,8900|true|false|false|||sedentary
Finding|Finding|Discharge Instructions|8891,8900|true|false|false|C1532253|Sedentary lifestyle|sedentary
Finding|Daily or Recreational Activity|Discharge Instructions|8902,8906|false|false|false|C0080331|Walking (function)|Walk
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|8919,8924|false|false|false|C1570446|TNFSF14 protein, human|Light
Drug|Biologically Active Substance|Discharge Instructions|8919,8924|false|false|false|C1570446|TNFSF14 protein, human|Light
Event|Event|Discharge Instructions|8919,8924|false|false|false|||Light
Finding|Finding|Discharge Instructions|8919,8924|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|Light
Finding|Functional Concept|Discharge Instructions|8919,8924|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|Light
Finding|Gene or Genome|Discharge Instructions|8919,8924|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|Light
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|8919,8924|false|false|false|C0023693|Light|Light
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8919,8924|false|false|false|C0031765|Phototherapy|Light
Finding|Finding|Discharge Instructions|8925,8941|false|false|false|C2136403|activity level doing household chores|household chores
Event|Event|Discharge Instructions|8935,8941|false|false|false|||chores
Event|Event|Discharge Instructions|8943,8950|false|false|false|||cooking
Finding|Daily or Recreational Activity|Discharge Instructions|8943,8950|false|false|false|C0335326|Cooking (activity)|cooking
Attribute|Clinical Attribute|Discharge Instructions|8961,8968|false|false|false|C1830411||laundry
Event|Event|Discharge Instructions|8961,8968|false|false|false|||laundry
Finding|Daily or Recreational Activity|Discharge Instructions|8961,8968|false|false|false|C1830412|Laundry|laundry
Event|Activity|Discharge Instructions|8970,8977|false|false|false|C0441648|Wash (cleansing action)|washing
Finding|Intellectual Product|Discharge Instructions|8970,8984|false|false|false|C4050473|Washing Dishes question|washing dishes
Event|Event|Discharge Instructions|8978,8984|false|false|false|||dishes
Event|Event|Discharge Instructions|9003,9004|false|false|false|||
Event|Event|Discharge Instructions|9023,9032|true|false|false|||straining
Finding|Physiologic Function|Discharge Instructions|9023,9032|true|false|false|C0442694|Straining (finding)|straining
Event|Event|Discharge Instructions|9034,9041|true|false|false|||pulling
Finding|Finding|Discharge Instructions|9034,9041|true|false|false|C0580846;C2584320|Does pull;Pulling|pulling
Finding|Organism Function|Discharge Instructions|9034,9041|true|false|false|C0580846;C2584320|Does pull;Pulling|pulling
Event|Event|Discharge Instructions|9043,9051|true|false|false|||twisting
Finding|Pathologic Function|Discharge Instructions|9043,9051|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Finding|Physiologic Function|Discharge Instructions|9043,9051|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|9060,9066|true|false|false|C0042221|Vacuum (physical force)|vacuum
Procedure|Health Care Activity|Discharge Instructions|9072,9080|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9081,9093|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9081,9093|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9081,9093|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

