CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Paxil|Drug|false|false||Paxil
null|Paxil|Drug|false|false||Paxilnull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Craniotomy|Procedure|false|false||craniotomynull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|Hardware Removal|Procedure|false|false||hardware removalnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||Craniotomynull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Involvement with|Finding|false|false||involvednull|Involved Anatomy|Modifier|false|false||involvednull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Precision - second|Finding|false|false||second
null|metastatic qualifier|Finding|false|false||second
null|Second Suffix|Finding|false|false||secondnull|seconds|Time|false|false||secondnull|Second Unit of Plane Angle|LabModifier|false|false||second
null|second (number)|LabModifier|false|false||secondnull|Craniotomy|Procedure|false|false||craniotomynull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Recurrent Malignant Neoplasm|Disorder|false|false||recurrencenull|Recurrence (disease attribute)|Finding|false|false||recurrencenull|Recurrence|Phenomenon|false|false||recurrencenull|penciclovir|Drug|false|false||PCV
null|penciclovir|Drug|false|false||PCVnull|Porcine circovirus|Disorder|false|false||PCVnull|Procarbazine-Lomustine-Vincristine (PCV) Regimen|Procedure|false|false||PCV
null|lomustine/procarbazine/vincristine|Procedure|false|false||PCV
null|Hematocrit Measurement|Procedure|false|false||PCVnull|area PCV|Anatomy|false|false||PCVnull|After Dinner|Time|false|false||PCVnull|Combid|Drug|false|false||comb
null|Combid|Drug|false|false||combnull|bleomycin/cyclophosphamide/methotrexate/vincristine protocol|Procedure|false|false||comb
null|bleomycin/cyclophosphamide/semustine/vincristine protocol|Procedure|false|false||combnull|Comb (body structure)|Anatomy|false|false||combnull|Comb (physical object)|Device|false|false||combnull|Chemotherapy Regimen|Procedure|false|false||chemo
null|Chemotherapy|Procedure|false|false||chemonull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Pruritus|Finding|false|false||pruritusnull|sensory perception of itch|Modifier|false|false||pruritusnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|husband|Subject|false|false||husbandnull|Personal appearance|Subject|false|false||looknull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|day|Time|false|false||daysnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Metals|Drug|false|false||metalnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|husband|Subject|false|false||husbandnull|Local Remote Control State - Local|Finding|false|false||localnull|Local|Modifier|false|false||localnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Nausea and vomiting|Finding|true|false||nausea vomitingnull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Vomiting|Finding|true|false||vomitingnull|nuchal|Modifier|false|false||nuchalnull|Muscle Rigidity|Finding|false|false||rigiditynull|plastic property - rigidity|Phenomenon|false|false||rigiditynull|Numbness or tingling|Finding|false|false||numbness or tinglingnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Has tingling sensation|Finding|false|false||tingling sensationnull|Paresthesia|Disorder|false|false||tinglingnull|Has tingling sensation|Finding|false|false||tinglingnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Intestines|Anatomy|false|false||bowelnull|Urinary incontinence due to bladder problem|Disorder|false|false||bladder incontinencenull|urinary incontinence by exam|Finding|false|false||bladder incontinence
null|Urinary Incontinence|Finding|false|false||bladder incontinencenull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Incontinence|Disorder|false|false||incontinencenull|new onset|Finding|true|false||new onsetnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Onset of (contextual qualifier)|Modifier|true|false||onsetnull|Age of Onset|LabModifier|true|false||onsetnull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Tremor|Finding|false|false||tremorsnull|Alveolar rhabdomyosarcoma|Disorder|false|false||armsnull|Adherence to Refills and Medications Scale|Finding|false|false||arms
null|KIDINS220 gene|Finding|false|false||armsnull|Upper arm|Anatomy|false|false||armsnull|null|Attribute|false|false||armsnull|Hyperthyroidism|Disorder|false|false||hyperthyroidnull|Disease|Disorder|false|false||diseasenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Left hemiparesis|Finding|false|false||left sided weaknessnull|Left sided|Modifier|false|false||left sided
null|Left|Modifier|false|false||left sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Ambulate|Finding|true|false||ambulatenull|Walkers|Device|true|false||walkernull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||Craniotomynull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Craniotomy|Procedure|false|false||craniotomynull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Disease|Disorder|false|false||diseasenull|Tubal Ligation|Procedure|false|false||tubal ligationnull|Ligation|Procedure|false|false||ligationnull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Acute bronchitis|Disorder|false|false||bronchitis
null|Bronchitis|Disorder|false|false||bronchitisnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Seizures|Finding|false|false||seizuresnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Alveolar rhabdomyosarcoma|Disorder|false|false||armsnull|Adherence to Refills and Medications Scale|Finding|false|false||arms
null|KIDINS220 gene|Finding|false|false||armsnull|Upper arm|Anatomy|false|false||armsnull|null|Attribute|false|false||armsnull|Trembling|Finding|false|false||tremulousnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hyperthyroidism|Disorder|false|false||hyperthyroidnull|Disease|Disorder|false|false||diseasenull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Mental Recall|Finding|false|false||Recallnull|Recall (activity)|Event|false|false||Recallnull|Physical object|Entity|false|false||objectsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|true|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|examination of extraocular movements|Procedure|true|false||Extraocular movementsnull|Extraocular|Finding|true|false||Extraocularnull|Movement|Finding|true|false||movementsnull|Gender Status - Intact|Finding|true|false||intactnull|Intact|Modifier|true|false||intactnull|Nystagmus|Disorder|true|false||nystagmusnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Palate|Anatomy|false|false||Palatalnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|true|false||Tongue midlinenull|Benign neoplasm of tongue|Disorder|true|false||Tonguenull|Procedure on tongue|Procedure|true|false||Tonguenull|Tongue|Anatomy|true|false||Tonguenull|midline cell component|Anatomy|true|false||midlinenull|Midline (qualifier value)|Modifier|true|false||midlinenull|Muscular fasciculation|Finding|true|false||fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Dyskinetic syndrome|Disorder|true|false||abnormal movementsnull|Abnormal movement|Finding|true|false||abnormal movementsnull|Observation Interpretation - Abnormal|Finding|true|false||abnormal
null|Abnormal|Finding|true|false||abnormalnull|Movement|Finding|true|false||movementsnull|Tremor|Finding|true|false||tremorsnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Power (Psychology)|Finding|false|false||powernull|Power|LabModifier|false|false||powernull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pronator drift|Finding|true|false||pronator driftnull|Observation of Sensation|Finding|true|false||Sensation
null|Sensory perception|Finding|true|false||Sensationnull|sensory exam|Procedure|true|false||Sensationnull|Sensation quality|Modifier|true|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Lower extremity>Toes|Anatomy|false|false||Toes
null|Toes|Anatomy|false|false||Toesnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Rapid|Modifier|false|false||rapidnull|Alternating|Finding|false|false||alternatingnull|Movement|Finding|false|false||movementsnull|Heel|Anatomy|false|false||heelnull|Shin|Anatomy|false|false||shinnull|CAT scan of head|Procedure|false|false||CT Headnull|null|Attribute|false|false||CT Headnull|Problems with head|Disorder|false|false||Headnull|Procedure on head|Procedure|false|false||Headnull|Structure of head of caudate nucleus|Anatomy|false|false||Head
null|Head|Anatomy|false|false||Headnull|Head Device|Device|false|false||Headnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Abscess formation|Finding|true|false||abscess formationnull|Abscess|Disorder|true|false||abscessnull|null|Finding|true|false||abscessnull|Formation|Finding|true|false||formationnull|Anabolism|Phenomenon|true|false||formationnull|Formations|Modifier|true|false||formationnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Postoperative Period|Time|false|false||postoperativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||mass
null|Mass of body structure|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Residual|Modifier|false|false||residualnull|Encephalomalacia|Disorder|false|false||encephalomalacianull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Similarity|Modifier|false|false||similarnull|Distribution [PK]|Finding|false|false||distribution
null|Distribution|Finding|false|false||distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Complaint (finding)|Finding|false|false||complaintsnull|Pruritus|Finding|false|false||itchynull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Examination and observation for unspecified reason|Finding|false|false||observation
null|null|Finding|false|false||observation
null|null|Finding|false|false||observation
null|Observation (finding)|Finding|false|false||observationnull|Observation - diagnostic procedure|Procedure|false|false||observation
null|Observation in research|Procedure|false|false||observation
null|Patient observation|Procedure|false|false||observationnull|Preoperative|Time|false|false||pre-operativenull|null|Finding|false|false||planning
null|Planned|Finding|false|false||planningnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Further|Modifier|false|false||furthernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Morning|Time|false|false||morningnull|Fit and well|Finding|false|false||fit
null|Prosthesis fit|Finding|false|false||fit
null|Fit by Myeloma Frailty Index|Finding|false|false||fit
null|Seizures|Finding|false|false||fitnull|Fecal Immunochemical Test|Procedure|false|false||fitnull|Fit (action)|Event|false|false||fitnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Pentasa|Drug|false|false||Pentasa
null|Pentasa|Drug|false|false||Pentasanull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|zolpidem|Drug|false|false||zolpidem
null|zolpidem|Drug|false|false||zolpidemnull|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl er
null|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl ernull|venlafaxine hydrochloride|Drug|false|false||venlafaxine hcl
null|venlafaxine hydrochloride|Drug|false|false||venlafaxine hclnull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|Flinders medical centre-7 marker|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hclnull|Hairy Cell Leukemia|Disorder|false|false||hclnull|promethazine|Drug|true|false||promethazine
null|promethazine|Drug|true|false||promethazinenull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Dosage|LabModifier|true|false||dosesnull|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Every six hours|Time|false|false||Q6Hnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|promethazine|Drug|false|false||promethazine
null|promethazine|Drug|false|false||promethazinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every six hours|Time|false|false||Q6Hnull|Hour|Time|false|false||hoursnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|cephalexin|Drug|false|false||cephalexin
null|cephalexin|Drug|false|false||cephalexinnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Every six hours|Time|false|false||Q6Hnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|day|Time|false|false||daysnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|zolpidem|Drug|false|false||zolpidem
null|zolpidem|Drug|false|false||zolpidemnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|mesalamine|Drug|false|false||mesalamine
null|mesalamine|Drug|false|false||mesalaminenull|Extended Release Oral Capsule|Drug|false|false||Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Extended Release Oral Capsule|Drug|false|false||Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Four times daily|Time|false|false||QIDnull|4 times|Finding|false|false||4 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|propylthiouracil|Drug|false|false||propylthiouracil
null|propylthiouracil|Drug|false|false||propylthiouracilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every eight hours|Time|false|false||Q8Hnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Every eight hours|Time|false|false||Q8Hnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Injury due to exposure to external cause|Disorder|false|false||exposurenull|exposure history|Finding|false|false||exposurenull|Accident due to exposure to weather conditions|Phenomenon|false|false||exposurenull|Exposure to|Modifier|false|false||exposurenull|Craniotomy|Procedure|false|false||craniotomynull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Relationship - Friend|Finding|false|false||friendnull|friend|Subject|false|false||friendnull|Family member|Subject|false|false||family membernull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Member Organization|Subject|false|false||member
null|Role Class - member|Subject|false|false||member
null|member|Subject|false|false||membernull|Surgical wound|Disorder|false|true||incisionnull|Surgical incisions|Procedure|false|true||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Daily|Time|false|false||dailynull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Lifting|Event|true|false||liftingnull|Straining (finding)|Finding|true|false||strainingnull|Excessive (qualifier value)|Modifier|true|false||excessivenull|Decompression Sickness|Disorder|false|false||bendingnull|Bending - Changing basic body position|Finding|false|false||bending
null|Does bend|Finding|false|false||bendingnull|Bent|Modifier|false|false||bendingnull|Hair Specimen Code|Finding|false|false||hair
null|Hair Specimen|Finding|false|false||hairnull|Hair|Anatomy|false|false||hairnull|Suture Joint|Anatomy|false|false||suturesnull|Surgical sutures|Device|false|false||suturesnull|Staple, Surgical|Device|false|false||staplesnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Fiber brand of calcium polycarbophil|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false||fibernull|Tissue fiber|Anatomy|false|false||fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||over the counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Doctor - Title|Finding|true|false||doctornull|Physicians|Subject|true|false||doctornull|Anti-Inflammatory Agents|Drug|true|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|true|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|true|false||medicinesnull|Motrin|Drug|true|false||Motrin
null|Motrin|Drug|true|false||Motrinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Etc.|Finding|false|false||etcnull|Clearance procedure|Procedure|false|false||Clearancenull|Clearance of substance|Attribute|false|false||Clearancenull|Clearance [PK]|Phenomenon|false|false||Clearancenull|Clearance|Modifier|false|false||Clearancenull|Work|Event|false|false||worknull|Postoperative Period|Time|false|false||post-operativenull|Office Visits|Procedure|false|false||office visitnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Visit|Finding|false|false||visitnull|Make - Instruction Imperative|Finding|false|false||Make
null|Manufacturer Name|Finding|false|false||Makenull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Continuous|Finding|false|false||continuenull|Incentive spirometry|Procedure|false|false||incentive spirometernull|Incentive Spirometers (device)|Device|false|false||incentive spirometernull|Incentives|Modifier|false|false||incentivenull|Spirometer Device|Device|false|false||spirometernull|At home|Finding|true|false||at homenull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|Call - dosing instruction fragment|Finding|false|false||CALL
null|Call (Instruction)|Finding|false|false||CALL
null|Decision|Finding|false|false||CALL
null|CHL1 gene|Finding|false|false||CALLnull|null|Attribute|false|false||SURGEONnull|Surgeon|Subject|false|false||SURGEONnull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Experience (Practice)|Finding|true|false||EXPERIENCE
null|Experience|Finding|true|false||EXPERIENCEnull|Following|Time|true|false||FOLLOWING
null|Status post|Time|true|false||FOLLOWINGnull|new onset|Finding|false|false||New onsetnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Tremor|Finding|false|false||tremorsnull|Seizures|Finding|false|false||seizuresnull|Confusion|Disorder|true|false||confusionnull|Clouded consciousness|Finding|true|false||confusionnull|Mental status changes|Finding|true|false||change in mental statusnull|null|Attribute|true|false||change in mental statusnull|Changing|Finding|true|false||change innull|Changed status|LabModifier|true|false||change innull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Changed status|LabModifier|true|false||change
null|Delta (difference)|LabModifier|true|false||changenull|Mental state|Finding|true|false||mental statusnull|null|Attribute|true|false||mental status
null|null|Attribute|true|false||mental statusnull|Psyche structure|Finding|true|false||mentalnull|What subject filter - Status|Finding|true|false||statusnull|null|Attribute|true|false||statusnull|Social status|Modifier|true|false||status
null|Status|Modifier|true|false||statusnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|true|false||tinglingnull|Has tingling sensation|Finding|true|false||tinglingnull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Headache|Finding|true|false||headachenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Traumatic Wound|Disorder|true|false||wound
null|Wounds and Injuries|Disorder|true|false||wound
null|Traumatic injury|Disorder|true|false||woundnull|Route of Administration - Wound|Finding|true|false||wound
null|null|Finding|true|false||wound
null|Specimen Type - Wound|Finding|true|false||woundnull|null|Finding|true|false||sitenull|Anatomic Site|Anatomy|true|false||sitenull|Study Site|Modifier|true|false||site
null|Site|Modifier|true|false||sitenull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than or Equal To|LabModifier|false|false||greater than or equal tonull|Greater Than or Equal To|LabModifier|false|false||greater than or equalnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Equal|Modifier|false|false||equal tonull|Relational Operator - Equal|Finding|false|false||equalnull|Equal|Modifier|false|false||equalnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions