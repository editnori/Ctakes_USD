 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|45,54|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|79,88|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Body Substance|Allergies|180,187|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|180,187|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|180,187|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Allergies|188,196|true|false|false|||recorded
Attribute|Clinical Attribute|Allergies|216,225|true|false|false|C1717415||Allergies
Event|Event|Allergies|216,225|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|216,225|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|229,234|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|Allergies|229,234|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|229,234|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|Allergies|237,246|true|false|false|||Attending
Finding|Functional Concept|Allergies|237,246|true|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|283,294|false|false|false|||overwhelmed
Event|Event|Chief Complaint|301,305|false|false|false|||felt
Disorder|Mental or Behavioral Dysfunction|Chief Complaint|306,314|false|false|false|C0438696|Suicidal|suicidal
Event|Event|Chief Complaint|306,314|false|false|false|||suicidal
Finding|Classification|Chief Complaint|320,325|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|326,334|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|326,334|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|338,356|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|347,356|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|347,356|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|347,356|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|347,356|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|347,356|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|394,397|true|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|394,397|true|false|false|||HPI
Finding|Finding|History of Present Illness|394,397|true|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|394,397|true|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|452,461|false|false|false|C0344315|Depressed mood|depressed
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|452,466|false|false|false|C0344315|Depressed mood|depressed mood
Attribute|Clinical Attribute|History of Present Illness|462,466|false|false|false|C2713234||mood
Event|Event|History of Present Illness|462,466|false|false|false|||mood
Finding|Conceptual Entity|History of Present Illness|462,466|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|History of Present Illness|462,466|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|History of Present Illness|462,466|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|471,478|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|History of Present Illness|471,478|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Sign or Symptom|History of Present Illness|471,487|false|false|false|C0860603|Anxiety symptoms|anxiety symptoms
Event|Event|History of Present Illness|479,487|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|479,487|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|479,487|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|History of Present Illness|489,494|false|false|false|C0030318|Panic|panic
Event|Event|History of Present Illness|504,508|false|false|false|||sent
Event|Event|History of Present Illness|519,533|false|false|false|||recommendation
Finding|Idea or Concept|History of Present Illness|519,533|false|false|false|C0034866|Recommendation|recommendation
Event|Event|History of Present Illness|546,555|false|false|false|||therapist
Event|Event|History of Present Illness|579,589|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|579,589|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|579,589|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|614,624|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|History of Present Illness|614,624|false|false|false|||depression
Finding|Functional Concept|History of Present Illness|614,624|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|History of Present Illness|614,624|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|630,639|false|false|false|C0178417|Anhedonia|anhedonia
Event|Event|History of Present Illness|630,639|false|false|false|||anhedonia
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|630,647|false|false|false|C3178803|Social Anhedonia|anhedonia, social
Finding|Functional Concept|History of Present Illness|641,647|false|false|false|C0728831|Social|social
Finding|Social Behavior|History of Present Illness|641,657|false|false|false|C0037421|Social isolation|social isolation
Event|Event|History of Present Illness|648,657|false|false|false|||isolation
Finding|Finding|History of Present Illness|648,657|false|false|false|C0037421;C0205409;C0260397;C1608299;C1608300|Isolated;Level of Care - Isolation;Need for isolation;Privacy Level - Isolation;Social isolation|isolation
Finding|Functional Concept|History of Present Illness|648,657|false|false|false|C0037421;C0205409;C0260397;C1608299;C1608300|Isolated;Level of Care - Isolation;Need for isolation;Privacy Level - Isolation;Social isolation|isolation
Finding|Idea or Concept|History of Present Illness|648,657|false|false|false|C0037421;C0205409;C0260397;C1608299;C1608300|Isolated;Level of Care - Isolation;Need for isolation;Privacy Level - Isolation;Social isolation|isolation
Finding|Social Behavior|History of Present Illness|648,657|false|false|false|C0037421;C0205409;C0260397;C1608299;C1608300|Isolated;Level of Care - Isolation;Need for isolation;Privacy Level - Isolation;Social isolation|isolation
Procedure|Laboratory Procedure|History of Present Illness|648,657|false|false|false|C0204727;C0220862|Isolation procedure;isolation aspects|isolation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|648,657|false|false|false|C0204727;C0220862|Isolation procedure;isolation aspects|isolation
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|660,670|false|false|false|C2825032|Withdrawal (dysfunction)|withdrawal
Event|Activity|History of Present Illness|660,670|false|false|false|C2349954|Withdraw (activity)|withdrawal
Event|Event|History of Present Illness|660,670|false|false|false|||withdrawal
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|660,670|false|false|false|C3812880|Withdrawal - birth control|withdrawal
Event|Event|History of Present Illness|672,682|false|false|false|||escalating
Event|Event|History of Present Illness|683,691|false|false|false|||feelings
Finding|Intellectual Product|History of Present Illness|683,691|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|History of Present Illness|683,691|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|History of Present Illness|683,700|false|false|false|C0018379|Guilt|feelings of guilt
Event|Event|History of Present Illness|695,700|false|false|false|||guilt
Finding|Mental Process|History of Present Illness|695,700|false|false|false|C0018379|Guilt|guilt
Finding|Intellectual Product|History of Present Illness|702,706|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Sign or Symptom|History of Present Illness|702,712|false|false|false|C0235162|Difficulty sleeping|poor sleep
Drug|Organic Chemical|History of Present Illness|707,712|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|History of Present Illness|707,712|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|History of Present Illness|707,712|false|false|false|||sleep
Finding|Organism Function|History of Present Illness|707,712|false|false|false|C0037313|Sleep|sleep
Disorder|Neoplastic Process|History of Present Illness|713,722|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|History of Present Illness|713,722|false|false|false|||secondary
Finding|Functional Concept|History of Present Illness|713,722|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|727,738|false|false|false|C0154575|Rumination Disorders|ruminations
Event|Event|History of Present Illness|727,738|false|false|false|||ruminations
Phenomenon|Biologic Function|History of Present Illness|727,738|false|false|false|C0232604|Rumination|ruminations
Event|Event|History of Present Illness|742,747|false|false|false|||guilt
Finding|Mental Process|History of Present Illness|742,747|false|false|false|C0018379|Guilt|guilt
Finding|Body Substance|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|773,780|false|false|false|||trouble
Event|Event|History of Present Illness|781,794|false|false|false|||concentrating
Event|Event|History of Present Illness|818,825|false|false|false|||classes
Finding|Intellectual Product|History of Present Illness|818,825|false|false|false|C0456387|Class|classes
Procedure|Health Care Activity|History of Present Illness|818,825|false|false|false|C4019422|Classes - encounter|classes
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|841,851|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|History of Present Illness|841,851|false|false|false|||depression
Finding|Functional Concept|History of Present Illness|841,851|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|History of Present Illness|841,851|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|856,863|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|856,863|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|856,863|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|History of Present Illness|878,884|false|false|false|||eating
Event|Activity|History of Present Illness|901,905|false|false|false|C1947933|care activity|care
Event|Event|History of Present Illness|901,905|false|false|false|||care
Finding|Finding|History of Present Illness|901,905|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|901,905|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|History of Present Illness|941,949|false|false|false|||reported
Event|Event|History of Present Illness|971,977|false|false|false|||caused
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|997,1004|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|997,1004|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|997,1004|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|History of Present Illness|1012,1023|false|false|false|||culmination
Attribute|Clinical Attribute|History of Present Illness|1027,1033|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|History of Present Illness|1027,1033|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|History of Present Illness|1027,1033|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|History of Present Illness|1027,1033|false|false|false|||stress
Finding|Finding|History of Present Illness|1027,1033|false|false|false|C0038435|Stress|stress
Finding|Idea or Concept|History of Present Illness|1039,1051|false|false|false|C1548286;C1571886|Charge type - professional;Entity Name Part Qualifier - professional|professional
Finding|Intellectual Product|History of Present Illness|1039,1051|false|false|false|C1548286;C1571886|Charge type - professional;Entity Name Part Qualifier - professional|professional
Event|Event|History of Present Illness|1052,1064|false|false|false|||relationship
Finding|Idea or Concept|History of Present Illness|1052,1064|false|false|false|C1705630;C1706279|Concept Relationship;Object Relationship|relationship
Event|Event|History of Present Illness|1081,1089|false|false|false|||teachers
Drug|Organic Chemical|History of Present Illness|1098,1105|false|false|false|C2728259|Program|program
Drug|Pharmacologic Substance|History of Present Illness|1098,1105|false|false|false|C2728259|Program|program
Event|Event|History of Present Illness|1098,1105|false|false|false|||program
Finding|Conceptual Entity|History of Present Illness|1098,1105|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Functional Concept|History of Present Illness|1098,1105|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Intellectual Product|History of Present Illness|1098,1105|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Event|Event|History of Present Illness|1112,1119|true|false|false|||reasons
Finding|Idea or Concept|History of Present Illness|1112,1119|true|false|false|C0392360|Indication of (contextual qualifier)|reasons
Finding|Intellectual Product|History of Present Illness|1133,1143|true|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|History of Present Illness|1144,1149|true|false|false|||clear
Finding|Idea or Concept|History of Present Illness|1144,1149|true|true|false|C1550016|Remote control command - Clear|clear
Finding|Body Substance|History of Present Illness|1151,1158|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1151,1158|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1151,1158|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1163,1170|true|false|false|||removed
Event|Event|History of Present Illness|1185,1190|false|false|false|||class
Finding|Classification|History of Present Illness|1185,1190|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Functional Concept|History of Present Illness|1185,1190|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Intellectual Product|History of Present Illness|1185,1190|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Event|Event|History of Present Illness|1209,1219|false|false|false|||instructor
Finding|Body Substance|History of Present Illness|1222,1229|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1222,1229|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1222,1229|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1230,1238|false|false|false|||referred
Finding|Finding|History of Present Illness|1245,1250|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Idea or Concept|History of Present Illness|1245,1250|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Individual Behavior|History of Present Illness|1245,1250|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Event|Event|History of Present Illness|1263,1270|false|false|false|||explain
Event|Event|History of Present Illness|1276,1285|false|false|false|||specifics
Event|Event|History of Present Illness|1303,1312|true|false|false|||available
Finding|Functional Concept|History of Present Illness|1303,1312|true|false|false|C0470187|Availability of|available
Finding|Body Substance|History of Present Illness|1317,1324|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1317,1324|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1317,1324|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1325,1329|true|false|false|||felt
Finding|Functional Concept|History of Present Illness|1370,1376|false|false|false|C1561567|detail - Response Level|detail
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1381,1385|false|false|false|C5552605|FACT Complex|fact
Drug|Biologically Active Substance|History of Present Illness|1381,1385|false|false|false|C5552605|FACT Complex|fact
Finding|Gene or Genome|History of Present Illness|1381,1385|false|false|false|C1420522;C5551287|SSRP1 wt Allele;SUPT16H gene|fact
Event|Event|History of Present Illness|1392,1397|false|false|false|||panic
Finding|Finding|History of Present Illness|1392,1397|false|false|false|C0030318|Panic|panic
Event|Event|History of Present Illness|1398,1404|false|false|false|||attack
Finding|Finding|History of Present Illness|1398,1404|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|History of Present Illness|1398,1404|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Event|Event|History of Present Illness|1416,1420|false|false|false|||talk
Finding|Finding|History of Present Illness|1416,1420|false|false|false|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Finding|Individual Behavior|History of Present Illness|1416,1420|false|false|false|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Finding|Organism Function|History of Present Illness|1416,1420|false|false|false|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Event|Event|History of Present Illness|1455,1462|false|false|false|||removed
Finding|Classification|History of Present Illness|1472,1477|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Functional Concept|History of Present Illness|1472,1477|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Intellectual Product|History of Present Illness|1472,1477|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Event|Event|History of Present Illness|1499,1506|true|false|false|||letters
Finding|Intellectual Product|History of Present Illness|1499,1506|true|false|false|C0282413||letters
Event|Event|History of Present Illness|1508,1514|true|false|false|||called
Event|Event|History of Present Illness|1531,1539|true|false|false|||messages
Finding|Intellectual Product|History of Present Illness|1531,1539|true|false|false|C0470166|Message|messages
Event|Event|History of Present Illness|1545,1552|true|false|false|||emailed
Event|Event|History of Present Illness|1558,1568|true|false|false|||instructor
Event|Event|History of Present Illness|1585,1593|true|false|false|||response
Finding|Finding|History of Present Illness|1585,1593|true|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|History of Present Illness|1585,1593|true|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|History of Present Illness|1585,1593|true|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|History of Present Illness|1608,1616|false|false|false|||response
Finding|Finding|History of Present Illness|1608,1616|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|History of Present Illness|1608,1616|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|History of Present Illness|1608,1616|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|History of Present Illness|1621,1627|false|false|false|||caused
Event|Event|History of Present Illness|1642,1649|false|false|false|||pattern
Event|Event|History of Present Illness|1653,1658|false|false|false|||guilt
Finding|Mental Process|History of Present Illness|1653,1658|false|false|false|C0018379|Guilt|guilt
Event|Event|History of Present Illness|1681,1688|false|false|false|||dealing
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1697,1704|false|false|false|C0424376|Cutting self|cutting
Event|Event|History of Present Illness|1697,1704|false|false|false|||cutting
Finding|Finding|History of Present Illness|1697,1704|false|false|false|C2321228|self-mutilation by cutting (history)|cutting
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1697,1704|false|false|false|C0152060|Transection (procedure)|cutting
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1727,1730|true|false|false|C0228549|Cuneate tubercle structure|cut
Disorder|Injury or Poisoning|History of Present Illness|1727,1730|true|false|false|C0000925|Incised wound|cut
Finding|Finding|History of Present Illness|1727,1730|true|false|false|C1413827;C2136694|CUX1 gene;reported cut of tissue (history)|cut
Finding|Gene or Genome|History of Present Illness|1727,1730|true|false|false|C1413827;C2136694|CUX1 gene;reported cut of tissue (history)|cut
Finding|Functional Concept|History of Present Illness|1731,1735|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1731,1741|true|false|false|C0230366|Structure of left wrist|left wrist
Anatomy|Body Location or Region|History of Present Illness|1736,1741|true|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Anatomy|Body Space or Junction|History of Present Illness|1736,1741|true|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Event|Event|History of Present Illness|1746,1754|true|false|false|||stitches
Event|Event|History of Present Illness|1777,1784|true|false|false|||context
Finding|Idea or Concept|History of Present Illness|1777,1784|true|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|History of Present Illness|1777,1784|true|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|History of Present Illness|1777,1784|true|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Event|Event|History of Present Illness|1793,1798|true|false|false|||guilt
Finding|Mental Process|History of Present Illness|1793,1798|true|false|false|C0018379|Guilt|guilt
Event|Event|History of Present Illness|1804,1812|true|false|false|||sleeping
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1829,1836|true|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|1829,1836|true|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|1829,1836|true|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|History of Present Illness|1846,1851|false|false|false|||began
Finding|Finding|History of Present Illness|1852,1868|false|false|false|C0424000|Feeling suicidal (finding)|feeling suicidal
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1860,1868|false|false|false|C0438696|Suicidal|suicidal
Event|Event|History of Present Illness|1860,1868|false|false|false|||suicidal
Event|Event|History of Present Illness|1873,1882|false|false|false|||developed
Event|Event|Plan|1894,1898|false|false|false|||kill
Event|Event|Plan|1944,1951|false|false|false|||decided
Event|Event|Plan|1980,1984|false|false|false|||deal
Event|Event|Plan|2007,2015|false|false|false|||feelings
Finding|Intellectual Product|Plan|2007,2015|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|Plan|2007,2015|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Disorder|Mental or Behavioral Dysfunction|Plan|2025,2032|false|false|false|C0812393|Cancer patients and suicide and depression|suicide
Event|Event|Plan|2025,2032|false|false|false|||suicide
Finding|Finding|Plan|2025,2032|false|false|false|C0038661|Suicide|suicide
Event|Event|Plan|2043,2047|false|false|false|||told
Event|Event|Plan|2052,2061|false|false|false|||counselor
Finding|Finding|Plan|2052,2061|false|false|true|C1561602|counselor|counselor
Event|Event|Plan|2075,2083|false|false|false|||thoughts
Finding|Idea or Concept|Plan|2075,2083|false|false|false|C0039869;C4319827|Thought|thoughts
Finding|Mental Process|Plan|2075,2083|false|false|false|C0039869;C4319827|Thought|thoughts
Event|Event|Plan|2092,2101|false|false|false|||counselor
Finding|Finding|Plan|2092,2101|false|false|false|C1561602|counselor|counselor
Event|Event|Plan|2102,2113|false|false|false|||recommended
Event|Event|Plan|2122,2126|false|false|false|||come
Event|Event|Plan|2149,2157|false|false|false|||reported
Event|Event|Plan|2170,2174|false|false|false|||felt
Finding|Idea or Concept|Plan|2210,2213|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Plan|2210,2213|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Plan|2224,2233|true|false|false|||impacting
Drug|Organic Chemical|Plan|2234,2239|true|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Plan|2234,2239|true|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Plan|2234,2239|true|false|false|||sleep
Finding|Organism Function|Plan|2234,2239|true|false|false|C0037313|Sleep|sleep
Event|Event|Plan|2243,2252|true|false|false|||resulting
Finding|Functional Concept|Plan|2269,2277|false|false|false|C0221099|Impaired|impaired
Finding|Finding|Plan|2269,2293|false|false|false|C3845552|Impaired decision-making|impaired decision-making
Event|Event|Plan|2278,2286|false|false|false|||decision
Finding|Mental Process|Plan|2278,2286|false|false|false|C0679006|Decision|decision
Finding|Mental Process|Plan|2278,2293|false|false|false|C0011109|Decision Making|decision-making
Event|Event|Plan|2287,2293|false|false|false|||making
Finding|Finding|Plan|2310,2318|false|false|false|C3843660|Too much|too much
Event|Event|Plan|2314,2318|false|false|false|||much
Finding|Finding|Plan|2314,2318|false|false|false|C4281574|Much|much
Finding|Behavior|Plan|2335,2341|false|false|false|C0036864|Sex Behavior|sexual
Finding|Social Behavior|Plan|2335,2355|false|false|false|C2371571|Sexual relationships|sexual relationships
Event|Event|Plan|2342,2355|false|false|false|||relationships
Finding|Idea or Concept|Plan|2357,2360|false|false|false|C1548556|Etc.|etc
Event|Event|Plan|2384,2385|true|false|false|||_
Disorder|Mental or Behavioral Dysfunction|Plan|2387,2396|false|false|false|C0033975|Psychotic Disorders|psychotic
Finding|Finding|Plan|2387,2396|false|false|false|C0459435|Psychotic symptom present|psychotic
Finding|Sign or Symptom|Plan|2387,2405|false|false|false|C0871189|Psychotic symptom|psychotic symptoms
Event|Event|Plan|2397,2405|false|false|false|||symptoms
Finding|Functional Concept|Plan|2397,2405|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Plan|2397,2405|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Mental Process|Plan|2429,2434|false|false|false|C0018379|Guilt|guilt
Event|Event|Plan|2439,2446|false|false|false|||reached
Disorder|Mental or Behavioral Dysfunction|Plan|2454,2463|false|false|false|C0033975|Psychotic Disorders|psychotic
Event|Event|Plan|2454,2463|false|false|false|||psychotic
Finding|Finding|Plan|2454,2463|false|false|false|C0459435|Psychotic symptom present|psychotic
Event|Event|Plan|2485,2491|false|false|false|||denied
Event|Event|Plan|2503,2508|true|false|false|||asked
Event|Event|Plan|2536,2543|true|false|false|||contact
Event|Event|Plan|2556,2561|true|false|false|||feels
Event|Event|Plan|2581,2590|true|false|false|||answering
Event|Event|Plan|2595,2600|true|false|false|||calls
Event|Event|Plan|2604,2614|true|false|false|||responding
Event|Event|Plan|2618,2624|true|false|false|||emails
Finding|Intellectual Product|Plan|2618,2624|true|false|false|C0013849|Email|emails
Event|Event|Plan|2625,2630|true|false|false|||means
Event|Event|Plan|2660,2664|true|false|false|||like
Event|Event|Plan|2674,2680|true|false|false|||denied
Event|Event|Plan|2685,2693|true|false|false|||thoughts
Finding|Idea or Concept|Plan|2685,2693|true|false|false|C0039869;C4319827|Thought|thoughts
Finding|Mental Process|Plan|2685,2693|true|false|false|C0039869;C4319827|Thought|thoughts
Event|Event|Plan|2697,2703|true|false|false|||trying
Event|Event|Plan|2707,2711|true|false|false|||harm
Event|Event|Plan|2716,2726|false|false|false|||instructor
Event|Event|Plan|2739,2747|false|false|false|||reported
Event|Event|Plan|2748,2755|false|false|false|||feeling
Disorder|Mental or Behavioral Dysfunction|Plan|2748,2763|false|false|false|C0003467|Anxiety|feeling anxious
Finding|Finding|Plan|2748,2763|false|false|false|C2239195|Anxious mood|feeling anxious
Disorder|Mental or Behavioral Dysfunction|Plan|2756,2763|false|false|false|C0003467|Anxiety|anxious
Event|Event|Plan|2756,2763|false|false|false|||anxious
Finding|Gene or Genome|Plan|2766,2771|false|false|false|C1424898|RXFP2 gene|great
Event|Event|Plan|2772,2776|false|false|false|||deal
Finding|Gene or Genome|Plan|2788,2792|false|false|false|C1514917|Retinoic Acid Response Element|rare
Finding|Finding|Plan|2793,2798|false|false|false|C0030318|Panic|panic
Disorder|Mental or Behavioral Dysfunction|Plan|2793,2805|false|false|false|C0086769|Panic Attacks|panic attack
Event|Event|Plan|2799,2805|false|false|false|||attack
Finding|Finding|Plan|2799,2805|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Plan|2799,2805|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2838,2843|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|Past Medical History|2838,2843|false|false|false|||PSYCH
Drug|Pharmacologic Substance|Past Medical History|2861,2871|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Past Medical History|2861,2871|true|false|false|||medication
Finding|Intellectual Product|Past Medical History|2861,2871|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Past Medical History|2872,2878|true|false|false|||trials
Event|Event|Past Medical History|2882,2893|true|false|false|||psychiatric
Finding|Finding|Past Medical History|2882,2893|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|Past Medical History|2882,2893|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2882,2893|true|false|false|C3526598|Psychiatric service|psychiatric
Event|Event|Past Medical History|2894,2910|true|false|false|||hospitalizations
Procedure|Health Care Activity|Past Medical History|2894,2910|true|false|false|C0019993|Hospitalization|hospitalizations
Event|Event|Past Medical History|2926,2933|false|false|false|||episode
Event|Event|Past Medical History|2943,2947|false|false|false|||kept
Event|Event|Past Medical History|2953,2964|false|false|false|||psychiatric
Finding|Finding|Past Medical History|2953,2964|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|Past Medical History|2953,2964|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2953,2964|false|false|false|C3526598|Psychiatric service|psychiatric
Event|Event|Past Medical History|2982,2989|false|false|false|||context
Finding|Idea or Concept|Past Medical History|2982,2989|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|Past Medical History|2982,2989|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|Past Medical History|2982,2989|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Anatomy|Body Location or Region|Past Medical History|3000,3005|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Past Medical History|3000,3005|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Past Medical History|3006,3010|false|false|false|C2598155||pain
Event|Event|Past Medical History|3006,3010|false|false|false|||pain
Finding|Functional Concept|Past Medical History|3006,3010|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Past Medical History|3006,3010|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Past Medical History|3017,3023|false|false|false|||turned
Finding|Finding|Past Medical History|3036,3041|false|false|false|C0030318|Panic|panic
Disorder|Mental or Behavioral Dysfunction|Past Medical History|3036,3048|false|true|false|C0086769|Panic Attacks|panic attack
Event|Event|Past Medical History|3042,3048|false|false|false|||attack
Finding|Finding|Past Medical History|3042,3048|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Past Medical History|3042,3048|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Event|Event|Past Medical History|3056,3066|false|false|false|||occasional
Finding|Finding|Past Medical History|3067,3072|false|false|false|C0030318|Panic|panic
Disorder|Mental or Behavioral Dysfunction|Past Medical History|3067,3080|false|false|false|C0086769|Panic Attacks|panic attacks
Event|Event|Past Medical History|3073,3080|false|false|false|||attacks
Finding|Finding|Past Medical History|3073,3080|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attacks
Finding|Social Behavior|Past Medical History|3073,3080|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attacks
Finding|Finding|Diagnosis|3137,3142|false|false|false|C0030318|Panic|panic
Event|Event|Diagnosis|3159,3165|false|false|false|||seeing
Event|Event|Diagnosis|3168,3177|false|false|false|||counselor
Finding|Finding|Diagnosis|3168,3177|false|false|false|C1561602|counselor|counselor
Finding|Gene or Genome|Diagnosis|3219,3222|true|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Idea or Concept|Diagnosis|3231,3235|true|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|Diagnosis|3231,3235|true|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Individual Behavior|Diagnosis|3231,3255|true|false|false|C0085271|Self-Injurious Behavior|self-injurious behaviors
Event|Event|Diagnosis|3246,3255|true|false|false|||behaviors
Finding|Behavior|Diagnosis|3246,3255|true|false|false|C0004927;C0677505|Behavior;Behaviors and observations relating to behavior|behaviors
Finding|Finding|Diagnosis|3246,3255|true|false|false|C0004927;C0677505|Behavior;Behaviors and observations relating to behavior|behaviors
Disorder|Mental or Behavioral Dysfunction|Diagnosis|3274,3282|false|false|false|C0438696|Suicidal|suicidal
Attribute|Clinical Attribute|Diagnosis|3274,3291|false|false|false|C5203396||suicidal ideation
Finding|Finding|Diagnosis|3274,3291|false|false|false|C5942421|Suicidal thoughts|suicidal ideation
Event|Event|Diagnosis|3283,3291|false|false|false|||ideation
Finding|Mental Process|Diagnosis|3283,3291|false|false|false|C0392348|ideation|ideation
Finding|Intellectual Product|Diagnosis|3305,3309|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Diagnosis|3355,3361|true|false|false|||intent
Finding|Idea or Concept|Diagnosis|3355,3361|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|Diagnosis|3355,3361|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Event|Event|Diagnosis|3380,3389|false|false|false|||counselor
Finding|Finding|Diagnosis|3380,3389|false|false|false|C1561602|counselor|counselor
Finding|Finding|Diagnosis|3393,3397|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Diagnosis|3393,3397|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Diagnosis|3393,3397|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Diagnosis|3393,3404|false|false|false|C0683862|high school level|high school
Event|Event|Diagnosis|3408,3412|false|false|false|||help
Event|Event|Diagnosis|3419,3425|false|false|false|||coping
Finding|Finding|Diagnosis|3419,3425|false|false|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Finding|Individual Behavior|Diagnosis|3419,3425|false|false|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Procedure|Therapeutic or Preventive Procedure|Diagnosis|3419,3425|false|false|false|C2700390;C3502819|COPING - Dental Restorative Procedure;COPING - Fixed Prosthodontics|coping
Event|Event|Diagnosis|3432,3439|false|false|false|||feeling
Finding|Mental Process|Diagnosis|3432,3439|false|false|false|C1527305|Feelings|feeling
Event|Event|Diagnosis|3440,3449|false|false|false|||different
Event|Event|Diagnosis|3470,3478|false|false|false|||reported
Event|Event|Diagnosis|3491,3499|false|false|false|||thoughts
Finding|Idea or Concept|Diagnosis|3491,3499|false|false|false|C0039869;C4319827|Thought|thoughts
Finding|Mental Process|Diagnosis|3491,3499|false|false|false|C0039869;C4319827|Thought|thoughts
Event|Event|Diagnosis|3503,3511|false|false|false|||fighting
Finding|Gene or Genome|Diagnosis|3547,3550|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Diagnosis|3568,3575|false|false|false|||started
Event|Event|Diagnosis|3579,3589|false|false|false|||counseling
Finding|Finding|Diagnosis|3579,3589|false|false|false|C0740209;C2148587|Encounter due to counseling;duration of counseling|counseling
Procedure|Health Care Activity|Diagnosis|3579,3589|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Procedure|Therapeutic or Preventive Procedure|Diagnosis|3579,3589|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Event|Event|Diagnosis|3594,3598|false|false|false|||said
Event|Event|Diagnosis|3610,3614|true|false|false|||want
Event|Event|Diagnosis|3618,3621|true|false|false|||get
Event|Event|Diagnosis|3644,3653|false|false|false|||situation
Event|Event|Diagnosis|3659,3663|false|false|false|||said
Event|Event|Diagnosis|3687,3691|false|false|false|||able
Finding|Finding|Diagnosis|3687,3691|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Diagnosis|3695,3699|false|false|false|||come
Attribute|Clinical Attribute|Diagnosis|3719,3725|false|false|false|C5890614||person
Event|Event|Diagnosis|3719,3725|false|false|false|||person
Finding|Intellectual Product|Diagnosis|3719,3725|false|false|false|C1522390|Person Info|person
Event|Event|Diagnosis|3730,3738|false|false|false|||fighting
Event|Event|Diagnosis|3744,3750|true|false|false|||denied
Disorder|Mental or Behavioral Dysfunction|Diagnosis|3759,3766|true|false|false|C0242151|Violent|violent
Event|Event|Diagnosis|3759,3766|true|false|false|||violent
Attribute|Clinical Attribute|Diagnosis|3767,3775|true|false|false|C2707008||behavior
Event|Event|Diagnosis|3767,3775|true|false|false|||behavior
Finding|Behavior|Diagnosis|3767,3775|true|false|false|C0004927|Behavior|behavior
Event|Event|Diagnosis|3778,3781|false|false|false|||PMH
Finding|Finding|Diagnosis|3778,3781|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Event|Event|Diagnosis|3820,3826|false|false|false|||repair
Finding|Functional Concept|Diagnosis|3820,3826|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Diagnosis|3820,3826|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Diagnosis|3820,3826|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Diagnosis|3820,3826|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Diagnosis|3820,3838|false|false|false|C0407887|Repair of meniscus|repair of meniscus
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|3830,3838|false|false|false|C0224498|Meniscus structure of joint|meniscus
Finding|Functional Concept|Diagnosis|3842,3846|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Diagnosis|3842,3851|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|3842,3851|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|Diagnosis|3847,3851|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|3847,3851|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Diagnosis|3847,3851|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Diagnosis|3847,3851|false|false|false|C0562271|Examination of knee joint|knee
Finding|Gene or Genome|Diagnosis|3867,3870|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Disorder|Neoplastic Process|Diagnosis|3871,3880|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Diagnosis|3871,3880|false|false|false|||secondary
Finding|Functional Concept|Diagnosis|3871,3880|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Injury or Poisoning|Diagnosis|3884,3890|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|Diagnosis|3884,3890|false|false|false|||injury
Event|Event|Diagnosis|3897,3904|false|false|false|||running
Event|Event|Diagnosis|3916,3925|true|false|false|||surgeries
Procedure|Therapeutic or Preventive Procedure|Diagnosis|3916,3925|true|false|false|C0543467|Operative Surgical Procedures|surgeries
Finding|Functional Concept|Patient History|3950,3956|false|false|false|C0728831|Social|SOCIAL
Finding|Finding|Patient History|3950,3963|false|false|false|C3841781|Social/family|SOCIAL/FAMILY
Finding|Classification|Patient History|3957,3963|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|FAMILY
Finding|Conceptual Entity|Patient History|3957,3963|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|FAMILY
Finding|Idea or Concept|Patient History|3957,3963|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|FAMILY
Finding|Intellectual Product|Patient History|3957,3963|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|FAMILY
Finding|Idea or Concept|Patient History|3974,3979|false|false|false|C1546495|Relationship - Child|child
Event|Event|Patient History|3980,3984|false|false|false|||born
Finding|Finding|Patient History|3992,4000|false|false|false|C0086170|Divorced state|divorced
Event|Event|Patient History|4001,4008|false|false|false|||parents
Event|Event|Patient History|4019,4028|false|false|false|||separated
Finding|Body Substance|Patient History|4034,4041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Patient History|4034,4041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Patient History|4034,4041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Patient History|4052,4058|false|false|false|||Raised
Finding|Idea or Concept|Patient History|4062,4068|false|false|false|C1546508|Relationship - Mother|mother
Event|Event|Patient History|4092,4104|false|false|false|||relationship
Finding|Idea or Concept|Patient History|4092,4104|false|false|false|C1705630;C1706279|Concept Relationship;Object Relationship|relationship
Event|Event|Patient History|4110,4116|false|false|false|||father
Finding|Conceptual Entity|Patient History|4110,4116|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Patient History|4110,4116|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Conceptual Entity|Patient History|4119,4125|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Patient History|4119,4125|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Patient History|4126,4135|false|false|false|||struggled
Drug|Organic Chemical|Patient History|4148,4155|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Patient History|4148,4155|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Patient History|4148,4155|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Mental or Behavioral Dysfunction|Patient History|4148,4166|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcohol dependence
Disorder|Mental or Behavioral Dysfunction|Patient History|4156,4166|false|false|false|C0439857|Dependence|dependence
Event|Event|Patient History|4156,4166|false|false|false|||dependence
Finding|Individual Behavior|Patient History|4156,4166|false|false|false|C0011546|emotional dependency|dependence
Event|Event|Patient History|4194,4199|false|false|false|||sober
Finding|Body Substance|Patient History|4202,4209|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Patient History|4202,4209|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Patient History|4202,4209|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Patient History|4210,4216|true|false|false|||denied
Event|Event|Patient History|4225,4233|true|false|false|||physical
Finding|Finding|Patient History|4225,4233|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Patient History|4225,4233|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Patient History|4225,4233|true|false|false|C0031809|Physical Examination|physical
Finding|Behavior|Patient History|4237,4243|true|false|false|C0036864|Sex Behavior|sexual
Disorder|Injury or Poisoning|Patient History|4237,4249|true|false|false|C0282350|Sexual abuse|sexual abuse
Disorder|Mental or Behavioral Dysfunction|Patient History|4244,4249|true|false|false|C0013146|Drug abuse|abuse
Event|Event|Patient History|4244,4249|true|false|false|||abuse
Event|Event|Patient History|4244,4249|true|false|false|C1546935|Abuse|abuse
Finding|Finding|Patient History|4244,4249|true|false|false|C0562381|Victim of abuse (finding)|abuse
Event|Event|Patient History|4257,4264|false|false|false|||growing
Event|Event|Patient History|4270,4279|false|false|false|||Described
Event|Event|Patient History|4280,4287|false|false|false|||feeling
Event|Event|Patient History|4289,4298|false|false|false|||different
Event|Event|Patient History|4311,4318|false|false|false|||trouble
Event|Event|Patient History|4319,4326|false|false|false|||fitting
Finding|Sign or Symptom|Patient History|4319,4326|false|false|false|C0036572|Seizures|fitting
Procedure|Health Care Activity|Patient History|4319,4326|false|false|false|C0441548||fitting
Event|Event|Patient History|4355,4362|true|false|false|||details
Finding|Behavior|Patient History|4375,4385|false|false|false|C0004927|Behavior|behavioral
Event|Event|Patient History|4386,4394|false|false|false|||troubles
Finding|Idea or Concept|Patient History|4410,4415|false|false|false|C1546495|Relationship - Child|child
Event|Event|Patient History|4421,4430|false|false|false|||suspended
Finding|Finding|Patient History|4440,4447|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|Patient History|4442,4447|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Patient History|4442,4447|false|false|false|||times
Finding|Finding|Patient History|4451,4455|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Patient History|4451,4455|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Patient History|4451,4455|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Patient History|4451,4462|false|false|false|C0683862|high school level|high school
Event|Event|Patient History|4456,4462|false|false|false|||school
Event|Event|Patient History|4464,4473|false|false|false|||struggled
Event|Event|Patient History|4496,4504|false|false|false|||graduate
Finding|Idea or Concept|Patient History|4496,4504|false|false|false|C1547183|School type - Graduate|graduate
Event|Governmental or Regulatory Activity|Patient History|4544,4548|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|Patient History|4552,4565|false|false|false|||concentration
Finding|Mental Process|Patient History|4552,4565|false|false|false|C0086045|Mental concentration|concentration
Finding|Finding|Patient History|4596,4605|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|Patient History|4606,4610|false|false|false|||time
Finding|Finding|Patient History|4606,4610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Patient History|4606,4610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Patient History|4606,4610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Patient History|4614,4619|false|false|false|C1552828|Table Frame - above|above
Event|Event|Patient History|4630,4635|false|false|false|||lives
Finding|Finding|Patient History|4636,4641|false|false|false|C0439044|Living Alone|alone
Phenomenon|Natural Phenomenon or Process|Patient History|4666,4673|true|false|false|C1705970|Electrical Current|current
Finding|Mental Process|Patient History|4674,4682|true|false|false|C0683275|romantic|romantic
Finding|Social Behavior|Patient History|4674,4696|true|false|false|C2371569|Romantic relationships|romantic relationships
Event|Event|Patient History|4683,4696|true|false|false|||relationships
Event|Event|Patient History|4737,4749|true|false|false|||relationship
Finding|Idea or Concept|Patient History|4737,4749|true|false|false|C1705630;C1706279|Concept Relationship;Object Relationship|relationship
Event|Event|Patient History|4750,4755|true|false|false|||ended
Event|Event|Patient History|4781,4785|true|false|false|||feel
Event|Event|Patient History|4795,4803|true|false|false|||continue
Event|Event|Patient History|4814,4820|true|false|false|||denied
Event|Event|Patient History|4825,4830|true|false|false|||legal
Finding|Conceptual Entity|Patient History|4825,4830|true|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|legal
Finding|Functional Concept|Patient History|4825,4830|true|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|legal
Finding|Intellectual Product|Patient History|4825,4830|true|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|legal
Event|Event|Patient History|4831,4839|true|false|false|||problems
Finding|Idea or Concept|Patient History|4831,4839|true|false|false|C1546466|Problems - What subject filter|problems
Event|Event|Patient History|4844,4850|true|false|false|||denied
Event|Event|Patient History|4858,4864|true|false|false|||access
Finding|Functional Concept|Patient History|4858,4864|true|false|false|C1554204|Role Class - access|access
Event|Event|Patient History|4872,4876|true|false|false|||guns
Event|Event|Family Medical History|4914,4924|false|false|false|||remarkable
Event|Event|Family Medical History|4929,4935|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|4929,4935|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|4929,4935|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Drug|Organic Chemical|Family Medical History|4941,4948|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Family Medical History|4941,4948|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Family Medical History|4941,4948|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Mental or Behavioral Dysfunction|Family Medical History|4941,4957|false|false|false|C0549393|Alcohol Problem|alcohol problems
Event|Event|Family Medical History|4949,4957|false|false|false|||problems
Finding|Idea or Concept|Family Medical History|4949,4957|false|false|false|C1546466|Problems - What subject filter|problems
Event|Event|Family Medical History|4958,4959|false|false|false|||(
Disorder|Neoplastic Process|Family Medical History|4962,4971|false|false|false|C0687702|Cancer Remission|remission
Event|Event|Family Medical History|4962,4971|false|false|false|||remission
Finding|Finding|Family Medical History|4962,4971|false|false|false|C0544452|Disease remission|remission
Event|Event|Family Medical History|4977,4983|false|false|false|||mother
Finding|Idea or Concept|Family Medical History|4977,4983|false|false|false|C1546508|Relationship - Mother|mother
Disorder|Disease or Syndrome|Family Medical History|4993,5007|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Event|Event|Family Medical History|4993,5007|false|false|false|||hypothyroidism
Event|Event|Family Medical History|5019,5025|true|false|false|||family
Finding|Classification|Family Medical History|5019,5025|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|5019,5025|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|5019,5025|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|5019,5025|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Family Medical History|5026,5033|true|false|false|||medical
Finding|Functional Concept|Family Medical History|5026,5033|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Family Medical History|5026,5033|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Family Medical History|5026,5033|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Family Medical History|5026,5033|true|false|false|C0199168|Medical service|medical
Finding|Finding|Family Medical History|5037,5048|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|Family Medical History|5037,5048|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5037,5048|true|false|false|C3526598|Psychiatric service|psychiatric
Disorder|Mental or Behavioral Dysfunction|Family Medical History|5037,5057|true|false|false|C1306597|Psychiatric problem|psychiatric problems
Event|Event|Family Medical History|5049,5057|true|false|false|||problems
Finding|Idea or Concept|Family Medical History|5049,5057|true|true|false|C1546466|Problems - What subject filter|problems
Event|Event|Family Medical History|5058,5063|false|false|false|||known
Finding|Body Substance|Family Medical History|5067,5074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|5067,5074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|5067,5074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|General Exam|5094,5097|false|false|false|C1414405;C3537320|ENO3 gene;MYELINATING SCHWANN CELL ELEMENT|MSE
Finding|Finding|General Exam|5122,5126|false|false|false|C1706180|Male Gender|male
Event|Event|General Exam|5128,5135|false|false|false|||dressed
Finding|Idea or Concept|General Exam|5139,5147|false|false|false|C1547192|Organization unit type - Hospital|hospital
Disorder|Mental or Behavioral Dysfunction|General Exam|5162,5169|false|false|false|C0003467|Anxiety|anxious
Event|Event|General Exam|5162,5169|false|false|false|||anxious
Finding|Finding|General Exam|5177,5182|false|false|false|C0030318|Panic|panic
Disorder|Mental or Behavioral Dysfunction|General Exam|5177,5189|false|false|false|C0086769|Panic Attacks|panic attack
Event|Event|General Exam|5183,5189|false|false|false|||attack
Finding|Finding|General Exam|5183,5189|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|General Exam|5183,5189|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Event|Activity|General Exam|5201,5210|false|false|false|C0021822|Interview|interview
Event|Event|General Exam|5201,5210|false|false|false|||interview
Finding|Intellectual Product|General Exam|5201,5210|false|false|false|C0935630|Published Interview|interview
Event|Event|General Exam|5213,5219|false|false|false|||Speech
Finding|Organism Function|General Exam|5213,5219|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|5213,5219|false|false|false|C0846595|Speech assessment|Speech
Finding|Finding|General Exam|5213,5226|false|false|false|C0395017||Speech normal
Event|Event|General Exam|5220,5226|false|false|false|||normal
Event|Activity|General Exam|5227,5231|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|5227,5231|false|false|false|||rate
Finding|Idea or Concept|General Exam|5227,5231|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|5233,5237|false|false|false|||tone
Event|Event|General Exam|5240,5246|false|false|false|||volume
Finding|Intellectual Product|General Exam|5240,5246|false|false|false|C1705102|Volume (publication)|volume
Attribute|Clinical Attribute|General Exam|5256,5264|false|false|false|C2706915||language
Event|Event|General Exam|5256,5264|false|false|false|||language
Finding|Intellectual Product|General Exam|5256,5264|false|false|false|C0033348|Programming Languages|language
Attribute|Clinical Attribute|General Exam|5267,5271|false|false|false|C2713234||Mood
Finding|Conceptual Entity|General Exam|5267,5271|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|5267,5271|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|5267,5271|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Disorder|Mental or Behavioral Dysfunction|General Exam|5276,5285|false|false|false|C0344315|Depressed mood|depressed
Event|Event|General Exam|5276,5285|false|false|false|||depressed
Finding|Finding|General Exam|5294,5305|false|false|false|C1444778|Constricting sensation quality|constricted
Event|Event|General Exam|5316,5321|false|false|false|||range
Finding|Intellectual Product|General Exam|5316,5321|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Disorder|Mental or Behavioral Dysfunction|General Exam|5325,5332|false|false|false|C0003467|Anxiety|anxious
Event|Event|General Exam|5333,5338|false|false|false|||realm
Finding|Idea or Concept|General Exam|5333,5338|false|false|false|C3244047|Realm|realm
Event|Event|General Exam|5341,5349|false|false|false|||Thoughts
Finding|Idea or Concept|General Exam|5341,5349|false|false|false|C0039869;C4319827|Thought|Thoughts
Finding|Mental Process|General Exam|5341,5349|false|false|false|C0039869;C4319827|Thought|Thoughts
Event|Event|General Exam|5350,5359|false|false|false|||organized
Finding|Functional Concept|General Exam|5350,5359|false|false|false|C1300196|Organized|organized
Event|Event|General Exam|5375,5380|false|false|false|||guilt
Finding|Mental Process|General Exam|5375,5380|false|false|false|C0018379|Guilt|guilt
Disorder|Mental or Behavioral Dysfunction|General Exam|5392,5400|false|false|false|C0438696|Suicidal|suicidal
Event|Event|General Exam|5392,5400|false|false|false|||suicidal
Attribute|Clinical Attribute|General Exam|5392,5409|false|false|false|C5203396||suicidal ideation
Finding|Finding|General Exam|5392,5409|false|false|false|C5942421|Suicidal thoughts|suicidal ideation
Event|Event|General Exam|5401,5409|false|false|false|||ideation
Finding|Mental Process|General Exam|5401,5409|false|false|false|C0392348|ideation|ideation
Disorder|Disease or Syndrome|General Exam|5415,5419|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|General Exam|5415,5419|false|false|false|||plan
Finding|Functional Concept|General Exam|5415,5419|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|General Exam|5415,5419|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|General Exam|5415,5419|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Drug|Organic Chemical|General Exam|5423,5429|false|false|false|C1171947|Commit Lozenge|commit
Drug|Pharmacologic Substance|General Exam|5423,5429|false|false|false|C1171947|Commit Lozenge|commit
Event|Event|General Exam|5423,5429|false|false|false|||commit
Procedure|Machine Activity|General Exam|5423,5429|false|false|false|C2347840|Commit Operation|commit
Disorder|Mental or Behavioral Dysfunction|General Exam|5430,5437|false|false|false|C0812393|Cancer patients and suicide and depression|suicide
Event|Event|General Exam|5430,5437|false|false|false|||suicide
Finding|Finding|General Exam|5430,5437|false|false|false|C0038661|Suicide|suicide
Event|Event|General Exam|5468,5479|false|false|false|||vacillating
Event|Event|General Exam|5480,5486|false|false|false|||intent
Finding|Idea or Concept|General Exam|5480,5486|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|General Exam|5480,5486|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Event|Event|General Exam|5496,5504|true|false|false|||thoughts
Finding|Idea or Concept|General Exam|5496,5504|true|false|false|C0039869;C4319827|Thought|thoughts
Finding|Mental Process|General Exam|5496,5504|true|false|false|C0039869;C4319827|Thought|thoughts
Event|Event|General Exam|5516,5522|true|false|false|||others
Event|Event|General Exam|5525,5532|false|false|false|||Insight
Finding|Mental Process|General Exam|5525,5532|false|false|false|C0233820|Insight|Insight
Event|Event|General Exam|5538,5542|false|false|false|||need
Finding|Functional Concept|General Exam|5538,5542|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Event|Event|General Exam|5547,5551|false|false|false|||help
Finding|Intellectual Product|General Exam|5547,5551|false|false|false|C1552861|Help document|help
Event|Event|General Exam|5555,5559|false|false|false|||good
Finding|Idea or Concept|General Exam|5555,5559|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|5561,5569|false|false|false|||judgment
Finding|Mental Process|General Exam|5561,5569|false|false|false|C0022423|Judgment|judgment
Drug|Biologically Active Substance|General Exam|5612,5619|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|5612,5619|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|5612,5619|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|5612,5619|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|5612,5619|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|5612,5619|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|5623,5627|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|5623,5627|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|5623,5627|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|5623,5627|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|5623,5627|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|5643,5649|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|5643,5649|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|5643,5649|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|5643,5649|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|5643,5649|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|5643,5649|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|5655,5664|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5655,5664|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|5655,5664|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|5655,5664|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|5655,5664|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|5655,5664|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|5655,5664|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5669,5677|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|5669,5677|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|5669,5677|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|5669,5677|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|5688,5691|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|5688,5691|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|5688,5691|false|false|false|||CO2
Finding|Finding|General Exam|5688,5691|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|5688,5691|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|5695,5700|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|5695,5704|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|5695,5704|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|5695,5704|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|5701,5704|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|5701,5704|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|5701,5704|false|false|false|||GAP
Finding|Gene or Genome|General Exam|5701,5704|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Attribute|Clinical Attribute|General Exam|5754,5757|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|5754,5757|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|5754,5757|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|5754,5757|false|false|false|C0040160|thyrotropin|TSH
Event|Event|General Exam|5754,5757|false|false|false|||TSH
Procedure|Laboratory Procedure|General Exam|5754,5757|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|5776,5779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|General Exam|5776,5779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|General Exam|5776,5779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|General Exam|5776,5779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|General Exam|5776,5779|false|false|false|||ASA
Finding|Gene or Genome|General Exam|5776,5779|false|false|false|C1412553|ARSA gene|ASA
Event|Event|General Exam|5780,5783|false|false|false|||NEG
Finding|Finding|General Exam|5780,5783|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|General Exam|5784,5791|false|false|false|C0161679|Toxic effect of ethyl alcohol|ETHANOL
Drug|Organic Chemical|General Exam|5784,5791|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Drug|Pharmacologic Substance|General Exam|5784,5791|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Event|Event|General Exam|5784,5791|false|false|false|||ETHANOL
Procedure|Laboratory Procedure|General Exam|5784,5791|false|false|false|C0202304|Ethanol measurement|ETHANOL
Event|Event|General Exam|5792,5795|false|false|false|||NEG
Finding|Finding|General Exam|5792,5795|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5806,5809|false|false|false|||NEG
Finding|Finding|General Exam|5806,5809|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|5820,5823|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5833,5836|false|false|false|||NEG
Finding|Finding|General Exam|5833,5836|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5847,5850|false|false|false|||NEG
Finding|Finding|General Exam|5847,5850|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|5863,5868|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5863,5868|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5863,5868|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|5876,5882|false|false|false|||RANDOM
Finding|Body Substance|General Exam|5895,5900|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5895,5900|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5895,5900|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|5908,5914|false|false|false|||RANDOM
Finding|Body Substance|General Exam|5927,5932|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5927,5932|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5927,5932|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Activity|General Exam|5937,5941|false|false|false|C1948035|Hold (action)|HOLD
Event|Event|General Exam|5937,5941|false|false|false|||HOLD
Finding|Functional Concept|General Exam|5937,5941|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Intellectual Product|General Exam|5937,5941|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Event|Activity|General Exam|5942,5946|false|false|false|C1948035|Hold (action)|HOLD
Event|Event|General Exam|5942,5946|false|false|false|||HOLD
Finding|Functional Concept|General Exam|5942,5946|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Intellectual Product|General Exam|5942,5946|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Body Substance|General Exam|5959,5964|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5959,5964|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5959,5964|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|5975,5978|false|false|false|||NEG
Finding|Finding|General Exam|5975,5978|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|5988,5991|false|false|false|C5848551|Neg - answer|NEG
Drug|Hazardous or Poisonous Substance|General Exam|5992,5999|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Organic Chemical|General Exam|5992,5999|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Pharmacologic Substance|General Exam|5992,5999|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Event|Event|General Exam|5992,5999|false|false|false|||opiates
Procedure|Laboratory Procedure|General Exam|5992,5999|false|false|false|C0242401|Opiate Measurement|opiates
Event|Event|General Exam|6000,6003|false|false|false|||NEG
Finding|Finding|General Exam|6000,6003|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|General Exam|6005,6012|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|General Exam|6005,6012|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|General Exam|6005,6012|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|General Exam|6005,6012|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|General Exam|6005,6012|false|false|false|C0009170|cocaine|cocaine
Event|Event|General Exam|6005,6012|false|false|false|||cocaine
Procedure|Laboratory Procedure|General Exam|6005,6012|false|false|false|C0202362|Cocaine measurement|cocaine
Event|Event|General Exam|6013,6016|false|false|false|||NEG
Finding|Finding|General Exam|6013,6016|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|6026,6029|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|6038,6041|false|false|false|||NEG
Finding|Finding|General Exam|6038,6041|false|false|false|C5848551|Neg - answer|NEG
Anatomy|Cell|General Exam|6056,6059|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6064,6067|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6064,6067|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6064,6067|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6073,6076|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|6073,6076|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|6073,6076|false|false|false|||HGB
Finding|Gene or Genome|General Exam|6073,6076|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|6073,6076|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|General Exam|6082,6085|false|false|false|||HCT
Procedure|Laboratory Procedure|General Exam|6082,6085|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|6082,6085|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|6091,6094|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|6091,6094|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|6091,6094|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6091,6094|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6091,6094|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6099,6102|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6099,6102|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6099,6102|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6099,6102|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6099,6102|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6099,6102|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6108,6112|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6108,6112|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Antibiotic|General Exam|6156,6161|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|6156,6161|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|6156,6161|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|6166,6169|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|General Exam|6166,6169|false|false|false|||EOS
Finding|Gene or Genome|General Exam|6166,6169|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|General Exam|6199,6202|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|6199,6202|false|false|false|C0201617|Primed lymphocyte test|PLT
Event|Event|General Exam|6225,6230|false|false|false|||URINE
Finding|Body Substance|General Exam|6225,6230|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6225,6230|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6225,6230|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|6225,6237|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|6232,6237|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6232,6237|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Finding|Idea or Concept|General Exam|6252,6257|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|6277,6282|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6277,6282|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6277,6282|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|6277,6289|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|6284,6289|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6284,6289|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6284,6289|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|6290,6293|false|false|false|||NEG
Finding|Finding|General Exam|6290,6293|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|6294,6301|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|6294,6301|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|6294,6301|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|6302,6305|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|6306,6313|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|6306,6313|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|General Exam|6306,6313|false|false|false|||PROTEIN
Finding|Conceptual Entity|General Exam|6306,6313|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|6306,6313|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|General Exam|6314,6317|false|false|false|||NEG
Finding|Finding|General Exam|6314,6317|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|6319,6326|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|6319,6326|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|6319,6326|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|6319,6326|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|6319,6326|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|6319,6326|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|General Exam|6327,6330|false|false|false|||NEG
Finding|Finding|General Exam|6327,6330|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|6331,6337|false|false|false|C0022634|Ketones|KETONE
Event|Event|General Exam|6338,6341|false|false|false|||NEG
Finding|Finding|General Exam|6338,6341|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|6342,6351|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|6342,6351|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|6342,6351|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|6342,6351|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|General Exam|6352,6355|false|false|false|||NEG
Finding|Finding|General Exam|6352,6355|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|6366,6369|false|false|false|||NEG
Finding|Finding|General Exam|6366,6369|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|6383,6386|false|false|false|||NEG
Finding|Finding|General Exam|6383,6386|false|false|false|C5848551|Neg - answer|NEG
Event|Event|Hospital Course|6415,6426|false|false|false|||Psychiatric
Finding|Finding|Hospital Course|6415,6426|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|Psychiatric
Finding|Functional Concept|Hospital Course|6415,6426|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|Psychiatric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6415,6426|false|false|false|C3526598|Psychiatric service|Psychiatric
Event|Event|Hospital Course|6431,6438|true|false|false|||arrived
Anatomy|Anatomical Structure|Hospital Course|6442,6447|true|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|6448,6455|false|false|false|||denying
Anatomy|Body Location or Region|Hospital Course|6464,6467|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|Hospital Course|6464,6467|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|Hospital Course|6479,6485|true|false|false|||intent
Finding|Idea or Concept|Hospital Course|6479,6485|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|Hospital Course|6479,6485|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Disorder|Disease or Syndrome|Hospital Course|6487,6491|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|6487,6491|false|false|false|||plan
Finding|Functional Concept|Hospital Course|6487,6491|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|6487,6491|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|6487,6491|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Hospital Course|6497,6505|false|false|false|||admitted
Disorder|Disease or Syndrome|Hospital Course|6509,6514|false|false|false|C1410088|Still|still
Event|Event|Hospital Course|6515,6522|false|false|false|||feeling
Attribute|Clinical Attribute|Hospital Course|6515,6532|false|false|false|C5671242||feeling depressed
Finding|Finding|Hospital Course|6515,6532|false|false|false|C0497307|Feeling depressed|feeling depressed
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6523,6532|false|false|false|C0344315|Depressed mood|depressed
Event|Event|Hospital Course|6523,6532|false|false|false|||depressed
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6534,6541|false|false|false|C0003467|Anxiety|anxious
Event|Event|Hospital Course|6534,6541|false|false|false|||anxious
Event|Event|Hospital Course|6550,6555|false|false|false|||eager
Finding|Mental Process|Hospital Course|6550,6555|false|false|false|C0558083|Enthusiastic|eager
Event|Event|Hospital Course|6560,6565|false|false|false|||start
Event|Event|Hospital Course|6566,6575|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|6566,6575|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6566,6575|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6566,6575|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6566,6575|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|Hospital Course|6580,6584|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|6580,6584|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|6580,6584|false|false|false|C4284232|Medications|meds
Drug|Organic Chemical|Hospital Course|6600,6606|false|false|false|C0719199|Celexa|celexa
Drug|Pharmacologic Substance|Hospital Course|6600,6606|false|false|false|C0719199|Celexa|celexa
Event|Event|Hospital Course|6600,6606|false|false|false|||celexa
Drug|Organic Chemical|Hospital Course|6618,6626|false|false|false|C0699315|Klonopin|klonopin
Drug|Pharmacologic Substance|Hospital Course|6618,6626|false|false|false|C0699315|Klonopin|klonopin
Event|Event|Hospital Course|6618,6626|false|false|false|||klonopin
Event|Event|Hospital Course|6631,6634|false|false|false|||QHS
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6643,6646|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6643,6646|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6643,6646|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6643,6646|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6652,6659|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|6652,6659|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|6652,6659|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|Hospital Course|6665,6672|false|false|false|||started
Event|Event|Hospital Course|6683,6690|true|false|false|||effects
Event|Event|Hospital Course|6695,6703|true|false|false|||reported
Finding|Idea or Concept|Hospital Course|6704,6715|true|false|false|C0750502|Significant|significant
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6716,6723|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|6716,6723|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|6716,6723|false|false|false|C0860603|Anxiety symptoms|anxiety
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6716,6733|false|false|false|C0150135|Alleviating anxiety|anxiety reduction
Event|Event|Hospital Course|6724,6733|false|false|false|||reduction
Finding|Finding|Hospital Course|6724,6733|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|6724,6733|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6724,6733|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Event|Event|Hospital Course|6739,6749|false|false|false|||resolution
Finding|Conceptual Entity|Hospital Course|6739,6749|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|6739,6749|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6753,6772|false|false|false|C0086132|Depressive Symptoms|depressive symptoms
Event|Event|Hospital Course|6764,6772|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|6764,6772|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|6764,6772|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|6818,6823|false|false|false|||urges
Event|Activity|Hospital Course|6839,6846|false|false|false|C1706079||arrival
Event|Event|Hospital Course|6839,6846|false|false|false|||arrival
Finding|Functional Concept|Hospital Course|6839,6846|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|Hospital Course|6851,6857|false|false|false|||stated
Event|Event|Hospital Course|6878,6889|false|false|false|||overreacted
Finding|Finding|Hospital Course|6915,6922|false|false|false|C3245517|Patient's teacher when immunized|teacher
Event|Event|Hospital Course|6928,6934|false|false|false|||wanted
Event|Event|Hospital Course|6941,6951|false|false|false|||discharged
Event|Event|Hospital Course|6969,6975|false|false|false|||return
Event|Event|Hospital Course|7000,7008|false|false|false|||speaking
Event|Event|Hospital Course|7019,7028|false|false|false|||counselor
Finding|Finding|Hospital Course|7019,7028|false|false|false|C1561602|counselor|counselor
Finding|Intellectual Product|Hospital Course|7050,7058|false|false|false|C3242376|Academic title|Academic
Event|Event|Hospital Course|7114,7122|false|false|false|||repeated
Event|Event|Hospital Course|7123,7127|false|false|false|||acts
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7131,7142|false|false|false|C0021125|Impulsive Behavior|impulsivity
Event|Event|Hospital Course|7131,7142|false|false|false|||impulsivity
Finding|Idea or Concept|Hospital Course|7144,7154|false|false|false|C0750541|apparently|apparently
Event|Event|Hospital Course|7165,7168|false|false|false|||got
Finding|Social Behavior|Hospital Course|7174,7179|false|false|false|C0424324|Fighting|fight
Event|Event|Hospital Course|7194,7201|false|false|false|||student
Event|Event|Hospital Course|7209,7216|false|false|false|||thought
Event|Event|Hospital Course|7221,7228|false|false|false|||talking
Finding|Intellectual Product|Hospital Course|7244,7248|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|7249,7252|false|false|false|||ran
Event|Event|Hospital Course|7285,7290|false|false|false|||asked
Anatomy|Body Location or Region|Hospital Course|7331,7337|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7331,7337|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Hospital Course|7331,7337|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Hospital Course|7331,7337|false|false|false|||throat
Finding|Body Substance|Hospital Course|7331,7337|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Hospital Course|7331,7337|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Hospital Course|7350,7356|false|false|false|||stated
Finding|Finding|Hospital Course|7377,7382|false|false|false|C2984081|Very Much|a lot
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7379,7382|false|false|false|C0162435;C0175218|Olfactory tract;nucleus of the lateral olfactory tract|lot
Finding|Idea or Concept|Hospital Course|7379,7382|false|false|false|C1710198|Stock (in-store merchandise)|lot
Event|Event|Hospital Course|7388,7395|false|false|false|||bridges
Finding|Finding|Hospital Course|7415,7422|false|false|false|C3245517|Patient's teacher when immunized|teacher
Event|Event|Hospital Course|7462,7470|false|false|false|||teachers
Disorder|Disease or Syndrome|Hospital Course|7482,7487|false|false|false|C1410088|Still|still
Event|Event|Hospital Course|7489,7498|false|false|false|||unwilling
Finding|Mental Process|Hospital Course|7489,7498|false|false|false|C0558080|Unwilling|unwilling
Event|Event|Hospital Course|7516,7520|false|false|false|||take
Event|Event|Hospital Course|7560,7570|false|false|false|||reputation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7574,7583|false|false|false|C0021125;C0564567|Impulsive Behavior;Impulsive character (finding)|impulsive
Event|Event|Hospital Course|7574,7583|false|false|false|||impulsive
Event|Event|Hospital Course|7591,7597|false|false|false|||stated
Disorder|Disease or Syndrome|Hospital Course|7602,7605|false|false|false|C0206695;C4082937|Carcinoma, Neuroendocrine;Necrotizing enterocolitis in fetus OR newborn|NEC
Disorder|Neoplastic Process|Hospital Course|7602,7605|false|false|false|C0206695;C4082937|Carcinoma, Neuroendocrine;Necrotizing enterocolitis in fetus OR newborn|NEC
Event|Event|Hospital Course|7602,7605|false|false|false|||NEC
Finding|Intellectual Product|Hospital Course|7602,7605|false|false|false|C2129066||NEC
Event|Event|Hospital Course|7610,7619|false|false|false|||recommend
Event|Event|Hospital Course|7623,7627|false|false|false|||take
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7632,7636|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|7632,7636|false|false|false|C1742913|REST protein, human|rest
Event|Event|Hospital Course|7632,7636|false|false|false|||rest
Finding|Daily or Recreational Activity|Hospital Course|7632,7636|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|7632,7636|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|7632,7636|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Functional Concept|Hospital Course|7660,7667|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|7660,7667|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|7660,7667|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|7660,7667|false|false|false|C0199168|Medical service|medical
Event|Activity|Hospital Course|7668,7673|false|false|false|C1706081||leave
Event|Event|Hospital Course|7668,7673|false|false|false|||leave
Finding|Functional Concept|Hospital Course|7668,7673|false|false|false|C5401409|Leave from Employment|leave
Event|Activity|Hospital Course|7687,7694|false|false|false|C0556656|Meetings|meeting
Event|Event|Hospital Course|7687,7694|false|false|false|||meeting
Finding|Intellectual Product|Hospital Course|7710,7718|false|false|false|C3242376|Academic title|academic
Finding|Body Substance|Hospital Course|7740,7747|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7740,7747|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7740,7747|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7766,7772|false|false|false|||agreed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7802,7806|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|7802,7806|false|false|false|C1742913|REST protein, human|rest
Event|Event|Hospital Course|7802,7806|false|false|false|||rest
Finding|Daily or Recreational Activity|Hospital Course|7802,7806|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|7802,7806|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|7802,7806|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Functional Concept|Hospital Course|7830,7837|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|7830,7837|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|7830,7837|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|7830,7837|false|false|false|C0199168|Medical service|medical
Finding|Finding|Hospital Course|7830,7854|false|false|false|C3841833|Medical leave of absence|medical leave of absence
Event|Activity|Hospital Course|7838,7843|false|false|false|C1706081||leave
Event|Event|Hospital Course|7838,7843|false|false|false|||leave
Finding|Functional Concept|Hospital Course|7838,7843|false|false|false|C5401409|Leave from Employment|leave
Finding|Intellectual Product|Hospital Course|7838,7854|false|false|false|C1549079|Leave of Absence - Inactive Reason Code|leave of absence
Procedure|Health Care Activity|Hospital Course|7838,7854|false|false|false|C1555555|Leave of Absence Supply|leave of absence
Disorder|Anatomical Abnormality|Hospital Course|7847,7854|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|Hospital Course|7847,7854|false|false|false|||absence
Finding|Functional Concept|Hospital Course|7847,7854|false|false|false|C0332197|Absent|absence
Event|Event|Hospital Course|7880,7889|false|false|false|||returning
Finding|Idea or Concept|Hospital Course|7890,7894|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Idea or Concept|Hospital Course|7895,7899|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|7895,7899|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Body Substance|Hospital Course|7905,7912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7905,7912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7905,7912|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7913,7919|false|false|false|||stated
Event|Event|Hospital Course|7928,7936|false|false|false|||speaking
Finding|Classification|Hospital Course|7946,7952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|7946,7952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|7946,7952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|7946,7952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Hospital Course|7968,7974|false|false|false|||return
Event|Event|Hospital Course|8005,8010|false|false|false|||close
Finding|Finding|Hospital Course|8005,8010|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|8005,8010|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Classification|Hospital Course|8018,8024|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|8018,8024|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|8018,8024|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|8018,8024|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Attribute|Clinical Attribute|Hospital Course|8037,8044|false|false|false|C1317973|Support - dental|support
Drug|Organic Chemical|Hospital Course|8037,8044|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Pharmacologic Substance|Hospital Course|8037,8044|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Vitamin|Hospital Course|8037,8044|false|false|false|C1171411|Support brand of multivitamin|support
Event|Event|Hospital Course|8037,8044|false|false|false|||support
Finding|Conceptual Entity|Hospital Course|8037,8044|false|false|false|C1521721|Supportive assistance|support
Procedure|Health Care Activity|Hospital Course|8037,8044|false|false|false|C0344211|Supportive care|support
Finding|Finding|Hospital Course|8058,8062|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|8058,8062|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|8058,8062|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Functional Concept|Hospital Course|8066,8073|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|8066,8073|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|8066,8073|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|8066,8073|false|false|false|C0199168|Medical service|medical
Event|Event|Hospital Course|8074,8080|false|false|false|||leave.
Event|Event|Hospital Course|8093,8099|false|false|false|||agreed
Event|Event|Hospital Course|8109,8115|false|false|false|||needed
Event|Event|Hospital Course|8119,8127|false|false|false|||continue
Event|Event|Hospital Course|8128,8134|false|false|false|||taking
Attribute|Clinical Attribute|Hospital Course|8139,8150|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|8139,8150|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|8139,8150|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|8139,8150|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|8161,8169|false|false|false|||followup
Procedure|Health Care Activity|Hospital Course|8161,8169|false|false|false|C1522577|follow-up|followup
Finding|Finding|Hospital Course|8176,8187|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|Hospital Course|8176,8187|false|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8176,8187|false|false|false|C3526598|Psychiatric service|psychiatric
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8176,8192|false|false|false|C0204523|Psychiatric therapeutic procedure|psychiatric care
Event|Activity|Hospital Course|8188,8192|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|8188,8192|false|false|false|||care
Finding|Finding|Hospital Course|8188,8192|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8188,8192|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Hospital Course|8234,8243|false|false|false|||satisfied
Finding|Intellectual Product|Hospital Course|8234,8243|false|false|false|C0242428;C4084799|Satisfaction;Satisfied|satisfied
Finding|Mental Process|Hospital Course|8234,8243|false|false|false|C0242428;C4084799|Satisfaction;Satisfied|satisfied
Finding|Mental Process|Hospital Course|8253,8259|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Hospital Course|8253,8266|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Hospital Course|8253,8266|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Hospital Course|8260,8266|false|false|false|C5889824||status
Event|Event|Hospital Course|8260,8266|false|false|false|||status
Finding|Idea or Concept|Hospital Course|8260,8266|false|false|false|C1546481|What subject filter - Status|status
Anatomy|Body Space or Junction|Hospital Course|8275,8280|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|Hospital Course|8275,8280|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|Hospital Course|8275,8280|false|false|false|C0575044|Joint problem|joint
Event|Activity|Hospital Course|8281,8288|false|false|false|C0556656|Meetings|meeting
Event|Event|Hospital Course|8294,8298|false|false|false|||felt
Event|Event|Hospital Course|8306,8310|true|false|false|||safe
Finding|Intellectual Product|Hospital Course|8306,8310|true|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|Hospital Course|8332,8341|true|false|false|||continued
Event|Activity|Hospital Course|8345,8349|false|false|false|C2700401|Deny (action)|deny
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8351,8361|true|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|8351,8361|true|false|false|||depression
Finding|Functional Concept|Hospital Course|8351,8361|true|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|8351,8361|true|false|false|C0460137;C1579931|Depression - motion|depression
Event|Event|Hospital Course|8367,8370|true|false|false|||SIB
Event|Event|Hospital Course|8383,8391|false|false|false|||oriented
Finding|Idea or Concept|Hospital Course|8396,8400|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|8396,8400|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|Hospital Course|8401,8409|false|false|false|||oriented
Event|Event|Hospital Course|8419,8425|false|false|false|||deemed
Event|Event|Hospital Course|8426,8430|false|false|false|||safe
Finding|Intellectual Product|Hospital Course|8426,8430|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|Hospital Course|8435,8444|false|false|false|||discharge
Finding|Body Substance|Hospital Course|8435,8444|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8435,8444|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8435,8444|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8435,8444|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|8457,8464|false|false|false|||Medical
Finding|Functional Concept|Hospital Course|8457,8464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|Hospital Course|8457,8464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|Hospital Course|8457,8464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|Hospital Course|8457,8464|false|false|false|C0199168|Medical service|Medical
Event|Event|Hospital Course|8476,8482|true|false|false|||issues
Finding|Idea or Concept|Hospital Course|8490,8498|true|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|8499,8503|true|false|false|||stay
Finding|Idea or Concept|Hospital Course|8509,8515|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|Groups
Finding|Intellectual Product|Hospital Course|8509,8515|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|Groups
Finding|Behavior|Hospital Course|8516,8526|false|false|false|C0004927|Behavior|Behavioral
Event|Event|Hospital Course|8540,8546|false|false|false|||groups
Finding|Idea or Concept|Hospital Course|8540,8546|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Finding|Intellectual Product|Hospital Course|8540,8546|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Event|Event|Hospital Course|8548,8556|false|false|false|||remained
Event|Event|Hospital Course|8557,8564|false|false|false|||visible
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8570,8574|false|false|false|C1366910|Calmodulin 1|calm
Drug|Biologically Active Substance|Hospital Course|8570,8574|false|false|false|C1366910|Calmodulin 1|calm
Event|Event|Hospital Course|8570,8574|false|false|false|||calm
Finding|Gene or Genome|Hospital Course|8570,8574|false|false|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Finding|Mental Process|Hospital Course|8570,8574|false|false|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8570,8574|false|false|false|C5552882|Cancer and Living Meaningfully Therapy|calm
Finding|Individual Behavior|Hospital Course|8610,8630|true|false|false|C0562573|Threatening behavior|threatening behavior
Attribute|Clinical Attribute|Hospital Course|8622,8630|true|false|false|C2707008||behavior
Event|Event|Hospital Course|8622,8630|true|false|false|||behavior
Finding|Behavior|Hospital Course|8622,8630|true|false|false|C0004927|Behavior|behavior
Event|Event|Hospital Course|8653,8659|false|false|false|||sitter
Event|Event|Hospital Course|8661,8669|true|false|false|||physical
Finding|Finding|Hospital Course|8661,8669|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|8661,8669|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|8661,8669|true|false|false|C0031809|Physical Examination|physical
Drug|Chemical|Hospital Course|8673,8681|true|false|false|C0220806|Chemicals|chemical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8673,8692|true|false|false|C1320374|Chemical restraint (procedure)|chemical restraints
Attribute|Clinical Attribute|Hospital Course|8682,8692|true|false|false|C2708180||restraints
Event|Event|Hospital Course|8682,8692|true|false|false|||restraints
Event|Event|Hospital Course|8693,8699|true|false|false|||needed
Finding|Finding|Hospital Course|8707,8711|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|8707,8711|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|8707,8711|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Conceptual Entity|Hospital Course|8717,8722|false|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|Legal
Finding|Functional Concept|Hospital Course|8717,8722|false|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|Legal
Finding|Intellectual Product|Hospital Course|8717,8722|false|false|false|C1301860;C1550438;C1550727|Entity Name Use - Legal;Legal;Organization Name Type - Legal|Legal
Attribute|Clinical Attribute|Hospital Course|8728,8739|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8728,8739|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8728,8739|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8728,8739|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8728,8752|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8743,8752|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8743,8752|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Hospital Course|8761,8770|true|false|false|||Discharge
Finding|Body Substance|Hospital Course|8761,8770|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8761,8770|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8761,8770|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8761,8770|true|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8761,8782|true|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8771,8782|true|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8771,8782|true|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8771,8782|true|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8771,8782|true|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8787,8797|false|false|false|C0008845|citalopram|Citalopram
Drug|Pharmacologic Substance|Hospital Course|8787,8797|false|false|false|C0008845|citalopram|Citalopram
Drug|Biomedical or Dental Material|Hospital Course|8804,8810|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8824,8830|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8824,8830|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|8858,8864|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|8869,8876|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8884,8894|false|false|false|C0009011|clonazepam|Clonazepam
Drug|Pharmacologic Substance|Hospital Course|8884,8894|false|false|false|C0009011|clonazepam|Clonazepam
Drug|Biomedical or Dental Material|Hospital Course|8902,8908|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8902,8908|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|8922,8928|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8922,8928|false|false|false|||Tablet
Event|Event|Hospital Course|8932,8935|false|false|false|||QAM
Event|Event|Hospital Course|8940,8943|false|false|false|||QHS
Drug|Biomedical or Dental Material|Hospital Course|8954,8960|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|8965,8972|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|8980,8989|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8980,8989|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8980,8989|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8980,8989|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8980,8989|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8980,9001|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8980,9001|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8990,9001|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8990,9001|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8990,9001|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|9003,9007|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|9003,9007|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9003,9007|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9003,9007|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|9010,9019|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9010,9019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9010,9019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9010,9019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9010,9019|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9010,9029|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9020,9029|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9020,9029|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9020,9029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9020,9029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9020,9029|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9031,9035|false|false|false|C0004457|Axis vertebra|Axis
Disorder|Injury or Poisoning|Hospital Course|9031,9035|false|false|false|C0349013|Fracture of second cervical vertebra|Axis
Finding|Classification|Hospital Course|9031,9037|false|false|false|C0221443|axis i|Axis I
Finding|Classification|Hospital Course|9039,9044|true|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9039,9064|true|false|false|C0041696;C1269683|Major Depressive Disorder;Unipolar Depression|Major depressive disorder
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9045,9064|true|false|false|C0011581|Depressive disorder|depressive disorder
Disorder|Disease or Syndrome|Hospital Course|9056,9064|true|false|false|C0012634|Disease|disorder
Event|Event|Hospital Course|9056,9064|true|false|false|||disorder
Finding|Finding|Hospital Course|9066,9072|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|9066,9072|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9082,9091|true|false|false|C0033975|Psychotic Disorders|psychotic
Event|Event|Hospital Course|9082,9091|true|false|false|||psychotic
Finding|Finding|Hospital Course|9082,9091|true|false|false|C0459435|Psychotic symptom present|psychotic
Finding|Finding|Hospital Course|9082,9100|true|false|false|C5436702|Psychotic features|psychotic features
Event|Event|Hospital Course|9092,9100|true|false|false|||features
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9101,9108|true|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|9101,9108|true|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|9101,9108|true|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9101,9117|true|false|false|C0003469|Anxiety Disorders|Anxiety disorder
Disorder|Disease or Syndrome|Hospital Course|9109,9117|true|false|false|C0012634|Disease|disorder
Event|Event|Hospital Course|9109,9117|true|false|false|||disorder
Event|Event|Hospital Course|9132,9141|true|false|false|||specified
Event|Event|Hospital Course|9146,9154|true|false|false|||deferred
Finding|Functional Concept|Hospital Course|9146,9154|true|false|false|C1554180;C1697785;C2347710|Protocol Deferred;Query Priority - Deferred;deferred - ResponseMode|deferred
Finding|Intellectual Product|Hospital Course|9146,9154|true|false|false|C1554180;C1697785;C2347710|Protocol Deferred;Query Priority - Deferred;deferred - ResponseMode|deferred
Attribute|Clinical Attribute|Hospital Course|9160,9166|false|false|false|C5889824||status
Event|Event|Hospital Course|9160,9166|false|false|false|||status
Finding|Idea or Concept|Hospital Course|9160,9166|false|false|false|C1546481|What subject filter - Status|status
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9172,9180|false|false|false|C0224498|Meniscus structure of joint|meniscus
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9172,9187|false|false|false|C0407887|Repair of meniscus|meniscus repair
Event|Event|Hospital Course|9181,9187|false|false|false|||repair
Finding|Functional Concept|Hospital Course|9181,9187|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Hospital Course|9181,9187|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Hospital Course|9181,9187|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9181,9187|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Anatomy|Body Location or Region|Hospital Course|9189,9193|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9189,9193|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Hospital Course|9189,9193|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Hospital Course|9189,9193|false|false|false|C0562271|Examination of knee joint|knee
Finding|Finding|Hospital Course|9199,9209|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Finding|Finding|Hospital Course|9210,9216|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|9210,9216|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9217,9229|false|false|false|C0740697|Psychosocial problem|psychosocial
Event|Event|Hospital Course|9217,9229|false|false|false|||psychosocial
Finding|Functional Concept|Hospital Course|9217,9229|false|false|false|C0542298|Psychosocial|psychosocial
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9217,9239|false|false|false|C0748073|psychosocial stressor|psychosocial stressors
Event|Event|Hospital Course|9230,9239|false|false|false|||stressors
Finding|Idea or Concept|Hospital Course|9230,9239|false|false|false|C0597530|Stressor|stressors
Event|Event|Hospital Course|9240,9250|false|false|false|||identified
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9254,9257|false|false|false|C1565805|FGF9 protein, human|GAF
Drug|Biologically Active Substance|Hospital Course|9254,9257|false|false|false|C1565805|FGF9 protein, human|GAF
Event|Event|Hospital Course|9254,9257|false|false|false|||GAF
Finding|Gene or Genome|Hospital Course|9254,9257|false|false|false|C1333540;C1708018|FGF9 gene;FGF9 wt Allele|GAF
Event|Event|Hospital Course|9263,9272|false|false|false|||discharge
Finding|Body Substance|Hospital Course|9263,9272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9263,9272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9263,9272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9263,9272|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Discharge Condition|9301,9304|false|false|false|||MSE
Finding|Gene or Genome|Discharge Condition|9301,9304|false|false|false|C1414405;C3537320|ENO3 gene;MYELINATING SCHWANN CELL ELEMENT|MSE
Event|Event|Discharge Condition|9305,9312|false|false|false|||general
Finding|Classification|Discharge Condition|9305,9312|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|Discharge Condition|9305,9312|false|false|false|C3812897|General medical service|general
Event|Event|Discharge Condition|9333,9339|false|false|false|||seated
Disorder|Disease or Syndrome|Discharge Condition|9341,9344|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Discharge Condition|9341,9344|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Discharge Condition|9341,9344|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Discharge Condition|9341,9344|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Discharge Condition|9341,9344|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Discharge Condition|9341,9344|true|false|false|||NAD
Finding|Finding|Discharge Condition|9341,9344|true|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Attribute|Clinical Attribute|Discharge Condition|9345,9353|true|false|false|C2707008||behavior
Event|Event|Discharge Condition|9345,9353|true|false|false|||behavior
Finding|Behavior|Discharge Condition|9345,9353|true|false|false|C0004927|Behavior|behavior
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|9355,9359|true|false|false|C1366910|Calmodulin 1|calm
Drug|Biologically Active Substance|Discharge Condition|9355,9359|true|false|false|C1366910|Calmodulin 1|calm
Event|Event|Discharge Condition|9355,9359|true|false|false|||calm
Finding|Gene or Genome|Discharge Condition|9355,9359|true|false|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Finding|Mental Process|Discharge Condition|9355,9359|true|false|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|9355,9359|true|false|false|C5552882|Cancer and Living Meaningfully Therapy|calm
Event|Event|Discharge Condition|9364,9371|true|false|false|||tremors
Finding|Sign or Symptom|Discharge Condition|9364,9371|true|false|false|C0040822|Tremor|tremors
Disorder|Disease or Syndrome|Discharge Condition|9376,9379|true|false|false|C0917981|Progressive Muscular Atrophy|PMA
Drug|Hazardous or Poisonous Substance|Discharge Condition|9376,9379|true|false|false|C0039654;C0048451|4-methoxyamphetamine;Tetradecanoylphorbol Acetate|PMA
Drug|Organic Chemical|Discharge Condition|9376,9379|true|false|false|C0039654;C0048451|4-methoxyamphetamine;Tetradecanoylphorbol Acetate|PMA
Drug|Pharmacologic Substance|Discharge Condition|9376,9379|true|false|false|C0039654;C0048451|4-methoxyamphetamine;Tetradecanoylphorbol Acetate|PMA
Event|Event|Discharge Condition|9376,9379|true|false|false|||PMA
Finding|Intellectual Product|Discharge Condition|9376,9379|true|false|false|C2825188|Premarket Device Application|PMA
Event|Event|Discharge Condition|9380,9386|true|false|false|||speech
Finding|Organism Function|Discharge Condition|9380,9386|true|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Discharge Condition|9380,9386|true|false|false|C0846595|Speech assessment|speech
Finding|Finding|Discharge Condition|9380,9394|true|false|false|C0395017||speech- normal
Event|Event|Discharge Condition|9388,9394|true|false|false|||normal
Event|Event|Discharge Condition|9400,9409|true|false|false|||pressured
Event|Event|Discharge Condition|9411,9417|true|false|false|||affect
Finding|Mental Process|Discharge Condition|9411,9417|true|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Discharge Condition|9411,9417|true|false|false|C2237113|assessment of affect|affect
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|9437,9445|false|false|false|C4722408|Reactive Therapy|reactive
Event|Event|Discharge Condition|9458,9464|false|false|false|||smiles
Finding|Finding|Discharge Condition|9458,9464|false|false|false|C0517048;C1883032|Simplified Molecular Input Line Entry Specification;Smiles (finding)|smiles
Finding|Intellectual Product|Discharge Condition|9458,9464|false|false|false|C0517048;C1883032|Simplified Molecular Input Line Entry Specification;Smiles (finding)|smiles
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|9505,9514|true|false|false|C0011253|Delusions|delusions
Event|Event|Discharge Condition|9505,9514|true|false|false|||delusions
Event|Event|Discharge Condition|9519,9522|true|false|false|||AVH
Finding|Idea or Concept|Discharge Condition|9538,9542|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Discharge Condition|9538,9542|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|Discharge Condition|9543,9551|false|false|false|||directed
Phenomenon|Human-caused Phenomenon or Process|Discharge Condition|9553,9559|true|false|false|C0036043|Safety|safety
Event|Event|Discharge Condition|9561,9567|false|false|false|||denies
Event|Event|Discharge Condition|9572,9575|true|false|false|||SIB
Event|Event|Discharge Condition|9577,9583|true|false|false|||intent
Finding|Idea or Concept|Discharge Condition|9577,9583|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|Discharge Condition|9577,9583|true|false|false|C0162425;C1550453|Act Mood - intent|intent
Disorder|Disease or Syndrome|Discharge Condition|9585,9589|true|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Discharge Condition|9585,9589|true|false|false|||plan
Finding|Functional Concept|Discharge Condition|9585,9589|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Discharge Condition|9585,9589|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Discharge Condition|9585,9589|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Gene or Genome|Discharge Condition|9591,9594|false|false|false|C1516685|Clusters of Orthologous Groups of Genes|cog
Attribute|Clinical Attribute|Discharge Instructions|9655,9666|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9655,9666|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9655,9666|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9655,9666|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9670,9680|false|false|false|||prescribed
Finding|Classification|Discharge Instructions|9696,9706|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|9696,9706|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Activity|Discharge Instructions|9707,9719|false|false|false|C0003629|Appointments|appointments
Event|Event|Discharge Instructions|9707,9719|false|false|false|||appointments
Event|Event|Discharge Instructions|9723,9732|false|false|false|||scheduled
Event|Event|Discharge Instructions|9745,9752|false|false|false|||feeling
Finding|Finding|Discharge Instructions|9745,9759|false|false|false|C5973924|feeling unsafe|feeling unsafe
Event|Event|Discharge Instructions|9753,9759|false|false|false|||unsafe
Attribute|Clinical Attribute|Discharge Instructions|9773,9782|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|9773,9782|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|9773,9782|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|9773,9782|false|false|false|C1705253|Logical Condition|condition
Event|Event|Discharge Instructions|9786,9795|false|false|false|||worsening
Finding|Idea or Concept|Discharge Instructions|9786,9795|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|Discharge Instructions|9798,9802|false|false|false|||call
Finding|Functional Concept|Discharge Instructions|9798,9802|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Discharge Instructions|9798,9802|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Discharge Instructions|9798,9802|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Discharge Instructions|9798,9802|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Event|Event|Discharge Instructions|9810,9812|false|false|false|||go
Procedure|Health Care Activity|Discharge Instructions|9835,9843|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9844,9856|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9844,9856|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9844,9856|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

