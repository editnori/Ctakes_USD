 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|45,54|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|79,88|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Organic Chemical|Allergies|182,189|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|182,189|false|false|false|C0009214|codeine|Codeine
Drug|Antibiotic|Allergies|192,201|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|192,201|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|204,211|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|Allergies|204,211|false|false|false|C0723778|Topamax|Topamax
Event|Event|Allergies|214,223|false|false|false|||Attending
Finding|Functional Concept|Allergies|214,223|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|249,252|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Chief Complaint|249,252|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Sign or Symptom|Chief Complaint|249,262|false|true|false|C0024031|Low Back Pain|Low back pain
Finding|Sign or Symptom|Chief Complaint|253,262|false|true|false|C0004604|Back Pain|back pain
Finding|Sign or Symptom|Chief Complaint|253,277|false|false|false|C0740363|Back Pain with Radiation|back pain with radiation
Attribute|Clinical Attribute|Chief Complaint|258,262|false|false|false|C2598155||pain
Event|Event|Chief Complaint|258,262|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|258,262|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|258,262|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Chief Complaint|268,277|false|false|false|||radiation
Phenomenon|Natural Phenomenon or Process|Chief Complaint|268,277|false|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|Chief Complaint|268,277|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|268,277|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Finding|Functional Concept|Chief Complaint|287,292|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|287,296|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|293,296|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Classification|Chief Complaint|300,305|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|306,314|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|306,314|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|318,336|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|327,336|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|327,336|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|327,336|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|327,336|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|327,336|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|338,351|false|false|false|||DECOMPRESSION
Finding|Functional Concept|Chief Complaint|338,351|false|false|false|C1965697|Decompression - action (qualifier value)|DECOMPRESSION
Phenomenon|Phenomenon or Process|Chief Complaint|338,351|false|false|false|C0011117|external decompression|DECOMPRESSION
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|338,351|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|DECOMPRESSION
Event|Event|Chief Complaint|359,365|false|false|false|||FUSION
Finding|Functional Concept|Chief Complaint|359,365|false|false|false|C0332466|Fused structure|FUSION
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|359,365|false|false|false|C1293131|Fusion procedure|FUSION
Event|Event|Chief Complaint|373,383|false|false|false|||DURAPLASTY
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|373,383|false|false|false|C0546551|Duraplasty|DURAPLASTY
Event|Event|History of Present Illness|457,464|false|false|false|||medical
Finding|Functional Concept|History of Present Illness|457,464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|457,464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|457,464|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|457,464|false|false|false|C0199168|Medical service|medical
Event|Event|History of Present Illness|466,473|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|466,473|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|466,473|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|466,473|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|474,485|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|474,485|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|490,498|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|History of Present Illness|490,507|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Event|Event|History of Present Illness|499,507|false|false|false|||aneurysm
Finding|Pathologic Function|History of Present Illness|499,507|false|false|false|C0002940|Aneurysm|aneurysm
Disorder|Anatomical Abnormality|History of Present Illness|499,525|false|false|false|C0162871|Aortic Aneurysm, Abdominal|aneurysm, abdominal aortic
Anatomy|Body Location or Region|History of Present Illness|509,518|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|519,525|false|false|false|C0003483|Aorta|aortic
Event|Event|History of Present Illness|527,535|false|false|false|||aneurysm
Finding|Pathologic Function|History of Present Illness|527,535|false|false|false|C0002940|Aneurysm|aneurysm
Disorder|Disease or Syndrome|History of Present Illness|537,562|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid syndrome
Disorder|Disease or Syndrome|History of Present Illness|554,562|false|false|false|C0039082|Syndrome|syndrome
Event|Event|History of Present Illness|554,562|false|false|false|||syndrome
Disorder|Disease or Syndrome|History of Present Illness|554,564|false|false|false|C0796110|Pallister W syndrome|syndrome w
Disorder|Disease or Syndrome|History of Present Illness|575,579|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|History of Present Illness|575,579|false|false|false|||DVTs
Event|Event|History of Present Illness|589,594|false|false|false|C0441471|Event|event
Finding|Gene or Genome|History of Present Illness|608,613|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|614,617|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|History of Present Illness|614,617|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|History of Present Illness|614,617|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|618,629|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|History of Present Illness|621,629|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|History of Present Illness|621,629|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|History of Present Illness|621,629|false|false|false|C0043031|warfarin|warfarin
Event|Event|History of Present Illness|621,629|false|false|false|||warfarin
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|631,636|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|History of Present Illness|631,636|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Event|Event|History of Present Illness|631,636|false|false|false|||BRCA1
Finding|Gene or Genome|History of Present Illness|631,636|false|false|false|C0376571|BRCA1 gene|BRCA1
Disorder|Cell or Molecular Dysfunction|History of Present Illness|631,645|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 mutation
Disorder|Cell or Molecular Dysfunction|History of Present Illness|637,645|false|false|false|C1705285|Mutation Abnormality|mutation
Event|Event|History of Present Illness|637,645|false|false|false|||mutation
Finding|Genetic Function|History of Present Illness|637,645|false|false|false|C0026882|Mutation|mutation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|658,664|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|658,664|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|History of Present Illness|658,664|false|false|false|||breast
Finding|Finding|History of Present Illness|658,664|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|658,664|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|History of Present Illness|658,671|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|History of Present Illness|665,671|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|665,671|false|false|false|||cancer
Event|Event|History of Present Illness|676,686|false|false|false|||lumpectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|676,686|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Event|Event|History of Present Illness|692,700|false|false|false|||presents
Event|Event|History of Present Illness|716,721|false|false|false|||month
Finding|Idea or Concept|History of Present Illness|716,721|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|716,721|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Functional Concept|History of Present Illness|725,730|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Sign or Symptom|History of Present Illness|725,746|false|true|false|C2219286|right-sided low back pain|right lower back pain
Anatomy|Body Location or Region|History of Present Illness|731,736|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|731,736|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|History of Present Illness|731,741|false|false|false|C0230102;C2939142|Lower back (surface region);Lower back structure|lower back
Finding|Sign or Symptom|History of Present Illness|731,746|false|true|false|C0024031|Low Back Pain|lower back pain
Finding|Sign or Symptom|History of Present Illness|737,746|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|History of Present Illness|742,746|false|true|false|C2598155||pain
Event|Event|History of Present Illness|742,746|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|742,746|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|742,746|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|752,766|false|false|false|C0278147|Radicular pain|radicular pain
Attribute|Clinical Attribute|History of Present Illness|762,766|false|false|false|C2598155||pain
Event|Event|History of Present Illness|762,766|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|762,766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|762,766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|History of Present Illness|777,782|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|777,786|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Finding|Sign or Symptom|History of Present Illness|777,791|false|true|false|C5848135|Pain in right leg|right leg pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|783,786|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|History of Present Illness|783,791|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|History of Present Illness|787,791|false|false|false|C2598155||pain
Event|Event|History of Present Illness|787,791|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|787,791|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|787,791|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|808,817|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|808,817|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Intellectual Product|History of Present Illness|826,831|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|833,842|false|false|false|||worsening
Finding|Idea or Concept|History of Present Illness|833,842|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Attribute|Clinical Attribute|History of Present Illness|850,854|false|false|false|C2598155||pain
Event|Event|History of Present Illness|850,854|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|850,854|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|850,854|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|859,867|false|false|false|||swelling
Finding|Finding|History of Present Illness|859,867|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|859,867|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Conceptual Entity|History of Present Illness|871,881|false|false|false|C1706907|Background|background
Finding|Functional Concept|History of Present Illness|901,906|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|901,910|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Finding|Sign or Symptom|History of Present Illness|901,915|false|true|false|C5848135|Pain in right leg|right leg pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|907,910|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|History of Present Illness|907,915|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|History of Present Illness|911,915|false|false|false|C2598155||pain
Event|Event|History of Present Illness|911,915|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|911,915|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|911,915|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|932,936|false|false|false|||show
Event|Event|History of Present Illness|937,945|false|false|false|||evidence
Finding|Idea or Concept|History of Present Illness|937,945|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|History of Present Illness|937,948|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Location or Region|History of Present Illness|949,952|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|949,952|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|949,952|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|History of Present Illness|949,952|false|false|false|||DVT
Event|Event|History of Present Illness|954,958|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|954,958|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|954,958|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|969,979|false|false|false|||consistent
Finding|Idea or Concept|History of Present Illness|969,979|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|History of Present Illness|969,984|false|false|false|C0332290|Consistent with|consistent with
Finding|Functional Concept|History of Present Illness|985,990|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|History of Present Illness|985,1012|false|false|false|C3862456|right trochanteric bursitis|right trochanteric bursitis
Disorder|Disease or Syndrome|History of Present Illness|991,1012|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|History of Present Illness|1004,1012|false|false|false|C0006444|Bursitis|bursitis
Event|Event|History of Present Illness|1004,1012|false|false|false|||bursitis
Drug|Organic Chemical|History of Present Illness|1032,1039|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|History of Present Illness|1032,1039|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1032,1049|false|false|false|C1261311|Injection of steroid|steroid injection
Drug|Biomedical or Dental Material|History of Present Illness|1040,1049|false|false|false|C1272883|Injection|injection
Event|Event|History of Present Illness|1040,1049|false|false|false|||injection
Finding|Functional Concept|History of Present Illness|1040,1049|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1040,1049|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Functional Concept|History of Present Illness|1055,1060|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1055,1066|false|false|false|C0817321|Right tibia|right tibia
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1061,1066|false|false|false|C0040184|Bone structure of tibia|tibia
Finding|Sign or Symptom|History of Present Illness|1061,1071|false|false|false|C0740426|Tibia pain|tibia pain
Attribute|Clinical Attribute|History of Present Illness|1067,1071|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1067,1071|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1067,1071|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1067,1071|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1076,1080|false|false|false|||felt
Disorder|Disease or Syndrome|History of Present Illness|1099,1113|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1108,1113|false|false|false|C0042449|Veins|veins
Event|Event|History of Present Illness|1108,1113|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1108,1113|false|false|false|C0398102|Procedure on vein|veins
Event|Event|History of Present Illness|1123,1132|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|1123,1132|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|History of Present Illness|1133,1140|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1133,1140|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|1141,1148|false|false|false|||notable
Event|Event|History of Present Illness|1156,1162|false|false|false|||Normal
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1163,1167|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Drug|Enzyme|History of Present Illness|1163,1167|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Event|Event|History of Present Illness|1166,1167|false|false|false|||A
Disorder|Disease or Syndrome|History of Present Illness|1182,1197|false|false|false|C0392525|Nephrolithiasis|nephrolithiasis
Event|Event|History of Present Illness|1182,1197|false|false|false|||nephrolithiasis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1206,1211|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|History of Present Illness|1206,1211|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|History of Present Illness|1206,1211|false|false|false|C0150920|Spine Problem|spine
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1218,1222|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|History of Present Illness|1218,1222|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|History of Present Illness|1218,1222|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|History of Present Illness|1218,1222|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|History of Present Illness|1218,1222|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Event|Event|History of Present Illness|1223,1228|false|false|false|||bulge
Finding|Finding|History of Present Illness|1223,1228|false|false|false|C0038999|Swelling|bulge
Event|Event|History of Present Illness|1247,1252|false|false|false|||cause
Finding|Conceptual Entity|History of Present Illness|1247,1252|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|History of Present Illness|1247,1252|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Finding|History of Present Illness|1253,1259|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|1253,1259|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Anatomical Abnormality|History of Present Illness|1260,1269|false|false|false|C3854333|Narrowing|narrowing
Event|Event|History of Present Illness|1260,1269|false|false|false|||narrowing
Anatomy|Body Space or Junction|History of Present Illness|1278,1290|false|false|false|C0037922|Spinal Canal|spinal canal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1285,1290|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Anatomy|Body Space or Junction|History of Present Illness|1285,1290|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Event|Event|History of Present Illness|1296,1304|false|false|false|||crowding
Finding|Finding|History of Present Illness|1296,1304|false|false|false|C0010383;C0040433|Crowding;Tooth Crowding|crowding
Finding|Social Behavior|History of Present Illness|1296,1304|false|false|false|C0010383;C0040433|Crowding;Tooth Crowding|crowding
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1323,1335|false|false|false|C0007458|Cauda Equina|cauda equina
Disorder|Neoplastic Process|History of Present Illness|1323,1335|false|false|false|C0349017|Malignant neoplasm of cauda equina|cauda equina
Disorder|Disease or Syndrome|History of Present Illness|1329,1335|false|false|false|C0017589|Glanders|equina
Disorder|Disease or Syndrome|Past Medical History|1362,1374|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Past Medical History|1362,1374|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|1377,1391|false|false|false|C0042345|Varicosity|Varicose veins
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1386,1391|false|false|false|C0042449|Veins|veins
Event|Event|Past Medical History|1386,1391|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1386,1391|false|false|false|C0398102|Procedure on vein|veins
Event|Event|Past Medical History|1402,1410|false|false|false|||ligation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1402,1410|false|false|false|C0023690|Ligation|ligation
Disorder|Disease or Syndrome|Past Medical History|1413,1417|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1413,1417|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1413,1417|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1413,1417|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|1420,1423|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1420,1423|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Past Medical History|1420,1423|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|Past Medical History|1420,1423|false|false|false|||OSA
Event|Event|Past Medical History|1426,1430|false|false|false|||CPap
Finding|Gene or Genome|Past Medical History|1426,1430|false|false|false|C1424863|CENPJ gene|CPap
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1426,1430|false|false|false|C0199451|Continuous Positive Airway Pressure|CPap
Finding|Finding|Past Medical History|1434,1444|false|false|false|C2169609|recent upper respiratory infection|recent URI
Disorder|Disease or Syndrome|Past Medical History|1441,1444|false|false|false|C0041912|Upper Respiratory Infections|URI
Event|Event|Past Medical History|1441,1444|false|false|false|||URI
Finding|Gene or Genome|Past Medical History|1441,1444|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|Past Medical History|1441,1444|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Event|Event|Past Medical History|1455,1461|false|false|false|||course
Drug|Antibiotic|Past Medical History|1465,1474|false|false|false|C0678143|Zithromax|Zithromax
Drug|Organic Chemical|Past Medical History|1465,1474|false|false|false|C0678143|Zithromax|Zithromax
Event|Event|Past Medical History|1465,1474|false|false|false|||Zithromax
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1488,1491|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|Past Medical History|1488,1491|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|Past Medical History|1488,1491|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1500,1525|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Drug|Immunologic Factor|Past Medical History|1500,1525|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Finding|Finding|Past Medical History|1500,1525|false|false|false|C4019436|Antiphospholipid antibody positivity|antiphospholipid antibody
Disorder|Disease or Syndrome|Past Medical History|1500,1534|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid antibody syndrome
Anatomy|Cell Component|Past Medical History|1517,1525|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1517,1525|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Past Medical History|1517,1525|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Past Medical History|1517,1525|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Event|Event|Past Medical History|1517,1525|false|false|false|||antibody
Procedure|Laboratory Procedure|Past Medical History|1517,1525|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Past Medical History|1526,1534|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Past Medical History|1526,1534|false|false|false|||syndrome
Event|Event|Past Medical History|1549,1564|false|false|false|||anticoagulation
Finding|Finding|Past Medical History|1549,1564|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Past Medical History|1549,1564|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1549,1564|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Past Medical History|1579,1582|false|false|false|||A1C
Finding|Classification|Past Medical History|1579,1582|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|Past Medical History|1579,1582|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1596,1604|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|Past Medical History|1596,1613|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Event|Event|Past Medical History|1605,1613|false|false|false|||aneurysm
Finding|Pathologic Function|Past Medical History|1605,1613|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|Past Medical History|1636,1645|false|false|false|||unchanged
Finding|Finding|Past Medical History|1636,1645|false|false|false|C0442739||unchanged
Disorder|Disease or Syndrome|Past Medical History|1649,1653|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1649,1653|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|1656,1670|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|Past Medical History|1656,1670|false|false|false|||diverticulosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1677,1682|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Past Medical History|1677,1682|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Past Medical History|1677,1682|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Past Medical History|1677,1682|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Anatomical Abnormality|Past Medical History|1677,1689|false|false|false|C0009376|Colonic Polyps|colon polyps
Disorder|Anatomical Abnormality|Past Medical History|1683,1689|false|false|false|C0032584|polyps|polyps
Event|Event|Past Medical History|1683,1689|false|false|false|||polyps
Finding|Intellectual Product|Past Medical History|1683,1689|false|false|false|C1546747||polyps
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1692,1702|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Past Medical History|1692,1702|false|false|false|||depression
Finding|Functional Concept|Past Medical History|1692,1702|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|1692,1702|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Functional Concept|Past Medical History|1709,1714|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Cell|Past Medical History|1715,1718|false|false|false|C3890599|Circulating Melanoma Cell|CMC
Disorder|Congenital Abnormality|Past Medical History|1715,1718|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Disorder|Disease or Syndrome|Past Medical History|1715,1718|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1715,1718|false|false|false|C0065772|MCC protocol|CMC
Anatomy|Body Space or Junction|Past Medical History|1719,1724|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|Past Medical History|1719,1724|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|Past Medical History|1719,1724|false|false|false|C0575044|Joint problem|joint
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1719,1737|false|false|false|C0003893|Arthroplasty|joint arthroplasty
Event|Event|Past Medical History|1725,1737|false|false|false|||arthroplasty
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1725,1737|false|false|false|C0003893;C0700235;C5887062|Arthroplasty;Reconstruction of joint;Temporomandibular joint arthroplasty by dentist|arthroplasty
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1744,1756|false|false|false|C0085515|Rotator Cuff|rotator cuff
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1744,1763|false|false|false|C0186666|Repair of musculotendinous cuff of shoulder|rotator cuff repair
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1752,1756|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|Past Medical History|1752,1756|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Event|Event|Past Medical History|1757,1763|false|false|false|||repair
Finding|Functional Concept|Past Medical History|1757,1763|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Past Medical History|1757,1763|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Past Medical History|1757,1763|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1757,1763|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|Past Medical History|1766,1774|false|false|false|||excision
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1766,1774|false|false|false|C0015252;C0728940|Excision;removal technique|excision
Finding|Functional Concept|Past Medical History|1775,1780|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1785,1790|false|false|false|C0582802|Digit structure|digit
Finding|Gene or Genome|Past Medical History|1785,1790|false|false|false|C4761764|GSC-DT gene|digit
Event|Event|Past Medical History|1791,1795|false|false|false|||mass
Finding|Finding|Past Medical History|1791,1795|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Past Medical History|1791,1795|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Past Medical History|1791,1795|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Past Medical History|1798,1801|false|false|false|||CCY
Event|Event|Past Medical History|1804,1809|false|false|false|||stone
Finding|Body Substance|Past Medical History|1804,1809|false|false|false|C0006736|Calculi|stone
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1812,1822|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1812,1822|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|Past Medical History|1812,1822|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|Past Medical History|1812,1822|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1812,1827|false|false|false|C0030288;C4482304|Abdomen>Pancreatic duct;Pancreatic duct|pancreatic duct
Disorder|Neoplastic Process|Past Medical History|1812,1827|false|false|false|C0153461|Malignant neoplasm of pancreatic duct|pancreatic duct
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1823,1827|false|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Event|Event|Past Medical History|1828,1839|false|false|false|||exploration
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1828,1839|false|false|false|C1280903|Exploration procedure|exploration
Event|Event|Past Medical History|1848,1860|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|1848,1860|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1848,1860|false|false|false|C0020699|Hysterectomy|hysterectomy
Event|Event|Past Medical History|1863,1876|false|false|false|||tonsillectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1863,1876|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Finding|Idea or Concept|Family Medical History|1917,1923|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1932,1939|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|1932,1946|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|1940,1946|false|false|false|C0006826|Malignant Neoplasms|CANCER
Attribute|Clinical Attribute|Family Medical History|1940,1949|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Family Medical History|1950,1953|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|1950,1953|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|1950,1953|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|1950,1953|false|false|false|||age
Finding|Conceptual Entity|Family Medical History|1959,1965|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1959,1965|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1974,1979|false|false|false|C0006104;C4266577|Brain;Head>Brain|BRAIN
Disorder|Disease or Syndrome|Family Medical History|1974,1979|false|false|false|C0006111|Brain Diseases|BRAIN
Disorder|Neoplastic Process|Family Medical History|1974,1986|false|false|false|C0006118;C0153633|Brain Neoplasms;Malignant neoplasm of brain|BRAIN CANCER
Disorder|Neoplastic Process|Family Medical History|1980,1986|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Family Medical History|1980,1986|false|false|false|||CANCER
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1988,1991|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Drug|Enzyme|Family Medical History|1988,1991|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Drug|Inorganic Chemical|Family Medical History|1988,1991|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Event|Event|Family Medical History|1988,1991|false|false|false|||PGM
Finding|Molecular Function|Family Medical History|1988,1991|false|false|false|C1150365|phosphoglycerate mutase activity|PGM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1992,1999|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|1992,2006|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|2000,2006|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Family Medical History|2000,2006|false|false|false|||CANCER
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2013,2020|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|2013,2027|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|2021,2027|false|false|false|C0006826|Malignant Neoplasms|CANCER
Disorder|Neoplastic Process|Family Medical History|2056,2074|false|false|false|C0007103;C0476089|Endometrial Carcinoma;Malignant neoplasm of endometrium|ENDOMETRIAL CANCER
Disorder|Neoplastic Process|Family Medical History|2068,2074|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Family Medical History|2068,2074|false|false|false|||CANCER
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2076,2079|false|false|false|C1366394;C3712803;C3887684|IGF1 protein, human;Kit Ligand, human;STAT5A protein, human|MGF
Drug|Biologically Active Substance|Family Medical History|2076,2079|false|false|false|C1366394;C3712803;C3887684|IGF1 protein, human;Kit Ligand, human;STAT5A protein, human|MGF
Finding|Gene or Genome|Family Medical History|2076,2079|false|false|false|C1335875;C1366480;C1704887;C1705050|KITLG gene;KITLG wt Allele;STAT5A gene;STAT5A wt Allele|MGF
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2080,2088|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|PROSTATE
Disorder|Disease or Syndrome|Family Medical History|2080,2088|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|PROSTATE
Disorder|Neoplastic Process|Family Medical History|2080,2088|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|PROSTATE
Disorder|Neoplastic Process|Family Medical History|2080,2095|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|PROSTATE CANCER
Disorder|Neoplastic Process|Family Medical History|2089,2095|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Family Medical History|2089,2095|false|false|false|||CANCER
Finding|Conceptual Entity|Family Medical History|2097,2104|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2097,2104|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2113,2119|false|false|false|C0022646;C0227665|Both kidneys;Kidney|KIDNEY
Disorder|Neoplastic Process|Family Medical History|2113,2119|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|KIDNEY
Event|Event|Family Medical History|2113,2119|false|false|false|||KIDNEY
Finding|Sign or Symptom|Family Medical History|2113,2119|false|false|false|C0812426|Kidney problem|KIDNEY
Procedure|Diagnostic Procedure|Family Medical History|2113,2119|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2113,2119|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Disorder|Neoplastic Process|Family Medical History|2113,2126|false|false|false|C0740457;C1378703|Malignant neoplasm of kidney;Renal carcinoma|KIDNEY CANCER
Disorder|Neoplastic Process|Family Medical History|2120,2126|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Family Medical History|2120,2126|false|false|false|||CANCER
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2129,2134|false|false|false|C0022646|Kidney|RENAL
Disorder|Disease or Syndrome|Family Medical History|2129,2134|false|false|false|C0042075|Urologic Diseases|RENAL
Disorder|Disease or Syndrome|Family Medical History|2129,2142|false|false|false|C0035078|Kidney Failure|RENAL FAILURE
Event|Event|Family Medical History|2135,2142|false|false|false|||FAILURE
Finding|Functional Concept|Family Medical History|2135,2142|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Family Medical History|2135,2142|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Family Medical History|2135,2142|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2156,2161|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|2156,2161|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|Family Medical History|2156,2161|false|false|false|||HEART
Finding|Sign or Symptom|Family Medical History|2156,2161|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|Family Medical History|2164,2171|false|false|false|||FAILURE
Finding|Functional Concept|Family Medical History|2164,2171|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Family Medical History|2164,2171|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Family Medical History|2164,2171|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Disorder|Disease or Syndrome|Family Medical History|2174,2182|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|DIABETES
Disorder|Disease or Syndrome|Family Medical History|2174,2191|false|false|false|C0011849|Diabetes Mellitus|DIABETES MELLITUS
Event|Event|Family Medical History|2183,2191|false|false|false|||MELLITUS
Drug|Hazardous or Poisonous Substance|Family Medical History|2194,2201|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Family Medical History|2194,2201|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Family Medical History|2194,2201|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Family Medical History|2194,2201|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2194,2207|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2202,2207|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Family Medical History|2202,2207|false|false|false|||ABUSE
Event|Event|Family Medical History|2202,2207|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Family Medical History|2202,2207|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Conceptual Entity|Substance Abuse Treatment|2225,2231|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|Sister
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|2240,2247|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Substance Abuse Treatment|2240,2254|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|2248,2254|false|false|false|C0006826|Malignant Neoplasms|CANCER
Attribute|Clinical Attribute|Substance Abuse Treatment|2248,2257|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Substance Abuse Treatment|2258,2261|false|false|false|C1114365||age
Drug|Biologically Active Substance|Substance Abuse Treatment|2258,2261|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Substance Abuse Treatment|2258,2261|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Substance Abuse Treatment|2258,2261|false|false|false|||age
Finding|Conceptual Entity|Substance Abuse Treatment|2267,2274|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Substance Abuse Treatment|2267,2274|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Anatomy|Body Location or Region|Substance Abuse Treatment|2279,2285|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|THROAT
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|2279,2285|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|THROAT
Drug|Pharmacologic Substance|Substance Abuse Treatment|2279,2285|false|false|false|C1950455|Throat Homeopathic Medication|THROAT
Finding|Body Substance|Substance Abuse Treatment|2279,2285|false|false|false|C1547926;C1550663|Specimen Type - Throat|THROAT
Finding|Intellectual Product|Substance Abuse Treatment|2279,2285|false|false|false|C1547926;C1550663|Specimen Type - Throat|THROAT
Disorder|Neoplastic Process|Substance Abuse Treatment|2279,2292|false|false|false|C0740339|Throat cancer|THROAT CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|2286,2292|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Substance Abuse Treatment|2286,2292|false|false|false|||CANCER
Attribute|Clinical Attribute|Substance Abuse Treatment|2286,2295|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Substance Abuse Treatment|2296,2299|false|false|false|C1114365||age
Drug|Biologically Active Substance|Substance Abuse Treatment|2296,2299|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Substance Abuse Treatment|2296,2299|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Substance Abuse Treatment|2296,2299|false|false|false|||age
Event|Event|Substance Abuse Treatment|2305,2309|false|false|false|||died
Event|Event|Substance Abuse Treatment|2320,2326|false|false|false|||Sister
Finding|Conceptual Entity|Substance Abuse Treatment|2320,2326|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|Sister
Drug|Amino Acid, Peptide, or Protein|Substance Abuse Treatment|2327,2332|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|Substance Abuse Treatment|2327,2332|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Finding|Gene or Genome|Substance Abuse Treatment|2327,2332|false|false|false|C0376571|BRCA1 gene|BRCA1
Disorder|Cell or Molecular Dysfunction|Substance Abuse Treatment|2327,2341|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 MUTATION
Disorder|Cell or Molecular Dysfunction|Substance Abuse Treatment|2333,2341|false|false|false|C1705285|Mutation Abnormality|MUTATION
Event|Event|Substance Abuse Treatment|2333,2341|false|false|false|||MUTATION
Finding|Genetic Function|Substance Abuse Treatment|2333,2341|false|false|false|C0026882|Mutation|MUTATION
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|2343,2349|false|false|false|C0006141|Breast|BREAST
Disorder|Neoplastic Process|Substance Abuse Treatment|2343,2349|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|BREAST
Event|Event|Substance Abuse Treatment|2343,2349|false|false|false|||BREAST
Finding|Finding|Substance Abuse Treatment|2343,2349|false|false|false|C0567499|Breast problem|BREAST
Procedure|Therapeutic or Preventive Procedure|Substance Abuse Treatment|2343,2349|false|false|false|C0191838|Procedures on breast|BREAST
Disorder|Neoplastic Process|Substance Abuse Treatment|2343,2356|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|BREAST CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|2350,2356|false|false|false|C0006826|Malignant Neoplasms|CANCER
Event|Event|Substance Abuse Treatment|2350,2356|false|false|false|||CANCER
Event|Event|Substance Abuse Treatment|2367,2373|false|false|false|||Living
Finding|Finding|Substance Abuse Treatment|2377,2385|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Idea or Concept|Substance Abuse Treatment|2377,2385|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Finding|Substance Abuse Treatment|2377,2395|false|false|false|C0476427|Abnormal cervical smear|ABNORMAL PAP SMEAR
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|2386,2389|false|false|false|C3496568|pars anterior of the paramedian lobule|PAP
Drug|Amino Acid, Peptide, or Protein|Substance Abuse Treatment|2386,2389|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Drug|Enzyme|Substance Abuse Treatment|2386,2389|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Drug|Immunologic Factor|Substance Abuse Treatment|2386,2389|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Finding|Finding|Substance Abuse Treatment|2386,2389|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Finding|Gene or Genome|Substance Abuse Treatment|2386,2389|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Finding|Molecular Function|Substance Abuse Treatment|2386,2389|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Procedure|Diagnostic Procedure|Substance Abuse Treatment|2386,2395|false|false|false|C0079104;C3541459|Pap smear;Papanicolaou Test|PAP SMEAR
Procedure|Laboratory Procedure|Substance Abuse Treatment|2386,2395|false|false|false|C0079104;C3541459|Pap smear;Papanicolaou Test|PAP SMEAR
Event|Activity|Substance Abuse Treatment|2390,2395|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Event|Event|Substance Abuse Treatment|2390,2395|false|false|false|||SMEAR
Finding|Functional Concept|Substance Abuse Treatment|2390,2395|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|Substance Abuse Treatment|2390,2395|false|false|false|C0444186|Smear test|SMEAR
Event|Event|Substance Abuse Treatment|2418,2421|false|false|false|||Son
Finding|Gene or Genome|Substance Abuse Treatment|2418,2421|false|false|false|C1420310|SON gene|Son
Attribute|Clinical Attribute|Substance Abuse Treatment|2431,2440|false|false|false|C5889933||SUBSTANCE
Drug|Substance|Substance Abuse Treatment|2431,2440|false|false|false|C0439861|Substance|SUBSTANCE
Finding|Intellectual Product|Substance Abuse Treatment|2431,2440|false|false|false|C5887067|administrative information regarding test substance|SUBSTANCE
Disorder|Mental or Behavioral Dysfunction|Substance Abuse Treatment|2431,2446|false|false|false|C0740858;C5967394|Harmful pattern of substance use;Substance Abuse Problems|SUBSTANCE ABUSE
Disorder|Mental or Behavioral Dysfunction|Substance Abuse Treatment|2441,2446|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Substance Abuse Treatment|2441,2446|false|false|false|||ABUSE
Event|Event|Substance Abuse Treatment|2441,2446|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Substance Abuse Treatment|2441,2446|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Disorder|Injury or Poisoning|Substance Abuse Treatment|2453,2459|false|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|Substance Abuse Treatment|2453,2459|false|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|Substance Abuse Treatment|2453,2459|false|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|Substance Abuse Treatment|2453,2459|false|false|false|C0011892|heroin|heroin
Disorder|Injury or Poisoning|Substance Abuse Treatment|2453,2468|false|false|false|C0572070|Heroin overdose|heroin overdose
Disorder|Injury or Poisoning|Substance Abuse Treatment|2460,2468|false|false|false|C0029944|Drug Overdose|overdose
Event|Event|Substance Abuse Treatment|2460,2468|false|false|false|||overdose
Finding|Finding|Substance Abuse Treatment|2460,2468|false|false|false|C1546941;C4018909|Event Qualification - Overdose;Overdose|overdose
Finding|Idea or Concept|Substance Abuse Treatment|2460,2468|false|false|false|C1546941;C4018909|Event Qualification - Overdose;Overdose|overdose
Finding|Finding|General Exam|2494,2502|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|General Exam|2494,2502|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|General Exam|2494,2502|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|General Exam|2494,2507|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|General Exam|2494,2507|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|General Exam|2503,2507|false|false|false|||Exam
Finding|Functional Concept|General Exam|2503,2507|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|2503,2507|false|false|false|C0582103|Medical Examination|Exam
Event|Event|General Exam|2511,2520|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|2511,2520|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|General Exam|2522,2528|false|false|false|||VITALS
Event|Event|General Exam|2540,2544|false|false|false|||Temp
Finding|Gene or Genome|General Exam|2540,2544|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|2540,2544|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Individual Behavior|General Exam|2567,2572|false|false|false|C0600261|Telling untruths|Lying
Event|Event|General Exam|2573,2575|false|false|false|||HR
Event|Event|General Exam|2602,2610|false|false|false|||delivery
Finding|Finding|General Exam|2602,2610|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|2602,2610|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|2602,2610|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|2602,2610|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|2617,2624|false|false|false|||General
Finding|Classification|General Exam|2617,2624|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|2617,2624|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|2626,2633|false|false|false|C0424109|Weepiness|Tearful
Event|Event|General Exam|2635,2645|false|false|false|||expressing
Finding|Functional Concept|General Exam|2646,2651|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|2652,2656|false|false|false|||back
Anatomy|Body Part, Organ, or Organ Component|General Exam|2661,2664|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|General Exam|2661,2669|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|General Exam|2665,2669|false|false|false|C2598155||pain
Event|Event|General Exam|2665,2669|false|false|false|||pain
Finding|Functional Concept|General Exam|2665,2669|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|2665,2669|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|2675,2681|false|false|false|||spasms
Finding|Sign or Symptom|General Exam|2675,2681|false|false|false|C0037763|Spasm|spasms
Anatomy|Body Location or Region|General Exam|2685,2690|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|2685,2690|false|false|false|C0741025|Chest problem|Chest
Anatomy|Body Part, Organ, or Organ Component|General Exam|2694,2700|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|2694,2700|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|General Exam|2694,2700|false|false|false|||breast
Finding|Finding|General Exam|2694,2700|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|2694,2700|false|false|false|C0191838|Procedures on breast|breast
Event|Event|General Exam|2701,2710|false|false|false|||incisions
Procedure|Therapeutic or Preventive Procedure|General Exam|2701,2710|false|false|false|C0184898|Surgical incisions|incisions
Finding|Finding|General Exam|2711,2715|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2716,2722|false|false|false|||healed
Finding|Functional Concept|General Exam|2716,2722|false|false|false|C0205249|Healed|healed
Anatomy|Body Location or Region|General Exam|2730,2736|false|false|false|C0004454|Axilla|axilla
Event|Event|General Exam|2737,2745|false|false|false|||surgical
Procedure|Health Care Activity|General Exam|2737,2745|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|General Exam|2737,2745|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Drug|Substance|General Exam|2746,2751|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|General Exam|2746,2751|false|false|false|||drain
Finding|Intellectual Product|General Exam|2746,2751|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|General Exam|2746,2759|false|false|false|C0411815|Removal of drain|drain removal
Event|Activity|General Exam|2752,2759|false|false|false|C1883720|Removing (action)|removal
Event|Event|General Exam|2752,2759|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|General Exam|2752,2759|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Activity|General Exam|2773,2777|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|2773,2777|false|false|false|||rate
Finding|Idea or Concept|General Exam|2773,2777|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|2782,2788|false|false|false|||rhythm
Finding|Finding|General Exam|2782,2788|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2782,2788|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|2809,2816|false|false|false|||murmurs
Finding|Finding|General Exam|2809,2816|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2817,2822|false|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|2824,2829|false|false|false|||Clear
Finding|Idea or Concept|General Exam|2824,2829|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|2833,2845|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|2833,2845|false|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|2862,2869|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|2862,2869|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|2873,2881|false|false|false|||crackles
Finding|Finding|General Exam|2873,2881|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|2882,2889|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2882,2889|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|2882,2889|false|false|false|||Abdomen
Finding|Finding|General Exam|2882,2889|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2891,2895|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|2891,2895|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|2924,2929|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|2924,2936|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|2930,2936|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|2930,2936|false|false|false|C0037709||sounds
Finding|Finding|General Exam|2937,2944|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|2937,2944|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Congenital Abnormality|General Exam|2945,2948|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|2945,2948|false|false|false|||Ext
Finding|Gene or Genome|General Exam|2945,2948|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|2950,2954|false|false|false|||Warm
Finding|Finding|General Exam|2950,2954|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2950,2954|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2956,2960|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2961,2969|false|false|false|||perfused
Finding|Functional Concept|General Exam|2971,2976|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|2971,2992|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|General Exam|2977,2982|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|2977,2982|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|2977,2992|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|2983,2992|false|false|false|C0015385|Limb structure|extremity
Event|Event|General Exam|2996,3002|false|false|false|||tender
Event|Event|General Exam|3006,3015|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|3006,3015|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|3020,3028|false|false|false|||movement
Finding|Organism Function|General Exam|3020,3028|false|false|false|C0026649|Movement|movement
Event|Event|General Exam|3029,3036|false|false|false|||limited
Attribute|Clinical Attribute|General Exam|3040,3044|false|false|false|C2598155||pain
Event|Event|General Exam|3040,3044|false|false|false|||pain
Finding|Functional Concept|General Exam|3040,3044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|3040,3044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|3046,3054|false|false|false|||Swelling
Finding|Finding|General Exam|3046,3054|false|false|false|C0013604;C0038999|Edema;Swelling|Swelling
Finding|Pathologic Function|General Exam|3046,3054|false|false|false|C0013604;C0038999|Edema;Swelling|Swelling
Event|Event|General Exam|3058,3061|false|false|false|||RLE
Event|Event|General Exam|3064,3067|false|false|false|||LLE
Drug|Food|General Exam|3085,3091|false|false|false|C5890763||pulses
Event|Event|General Exam|3085,3091|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3085,3091|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3085,3091|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body System|General Exam|3105,3109|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|3105,3109|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|3105,3109|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|3105,3109|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|3105,3109|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|3111,3115|false|false|false|||Warm
Finding|Finding|General Exam|3111,3115|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3111,3115|false|false|false|C0687712|warming process|Warm
Disorder|Disease or Syndrome|General Exam|3122,3136|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|3131,3136|false|false|false|C0042449|Veins|veins
Event|Event|General Exam|3131,3136|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|General Exam|3131,3136|false|false|false|C0398102|Procedure on vein|veins
Event|Event|General Exam|3137,3142|false|false|false|||noted
Anatomy|Body Location or Region|General Exam|3146,3151|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|3146,3151|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|3146,3163|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3152,3163|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|3181,3189|false|false|false|||oriented
Finding|Finding|General Exam|3181,3189|false|false|false|C1961028|Oriented to place|oriented
Disorder|Congenital Abnormality|General Exam|3190,3193|false|false|false|C0022681|Medullary sponge kidney|MSK
Disorder|Disease or Syndrome|General Exam|3190,3193|false|false|false|C0022681|Medullary sponge kidney|MSK
Event|Event|General Exam|3190,3193|false|false|false|||MSK
Finding|Gene or Genome|General Exam|3190,3193|false|false|false|C1420279|SIK1 gene|MSK
Event|Event|General Exam|3194,3198|false|false|false|||exam
Finding|Functional Concept|General Exam|3194,3198|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3194,3198|false|false|false|C0582103|Medical Examination|exam
Finding|Functional Concept|General Exam|3200,3205|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Space or Junction|General Exam|3206,3214|false|false|false|C5453012|SI joint|SI Joint
Anatomy|Body Space or Junction|General Exam|3209,3214|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Anatomy|Body System|General Exam|3209,3214|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Finding|Finding|General Exam|3209,3214|false|false|false|C0575044|Joint problem|Joint
Finding|Sign or Symptom|General Exam|3209,3225|false|false|false|C0240094|Joint tenderness|Joint tenderness
Event|Event|General Exam|3215,3225|false|false|false|||tenderness
Finding|Mental Process|General Exam|3215,3225|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3215,3225|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3227,3241|false|false|false|C0278147|Radicular pain|Radicular pain
Attribute|Clinical Attribute|General Exam|3237,3241|false|false|false|C2598155||pain
Event|Event|General Exam|3237,3241|false|false|false|||pain
Finding|Functional Concept|General Exam|3237,3241|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|3237,3241|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|3242,3250|false|false|false|||worsened
Attribute|Clinical Attribute|General Exam|3262,3269|false|false|false|C1525443|W flexion|flexion
Event|Event|General Exam|3262,3269|false|false|false|||flexion
Finding|Organ or Tissue Function|General Exam|3262,3269|false|false|false|C0231452||flexion
Event|Event|General Exam|3274,3282|false|false|false|||relieved
Event|Event|General Exam|3288,3297|false|false|false|||extension
Finding|Conceptual Entity|General Exam|3288,3297|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Finding|Functional Concept|General Exam|3288,3297|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Event|Event|General Exam|3303,3311|false|false|false|||strength
Finding|Idea or Concept|General Exam|3303,3311|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|3327,3330|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|3327,3330|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|3327,3330|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|3327,3330|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|3327,3330|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|3327,3330|false|false|false|C1292890|Procedure on hip|hip
Finding|Finding|General Exam|3327,3338|false|false|false|C2237371|Hip flexion|hip flexion
Attribute|Clinical Attribute|General Exam|3331,3338|false|false|false|C1525443|W flexion|flexion
Event|Event|General Exam|3331,3338|false|false|false|||flexion
Finding|Organ or Tissue Function|General Exam|3331,3338|false|false|false|C0231452||flexion
Event|Event|General Exam|3343,3352|false|false|false|||extension
Finding|Conceptual Entity|General Exam|3343,3352|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Finding|Functional Concept|General Exam|3343,3352|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Anatomy|Body Location or Region|General Exam|3354,3358|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|3354,3358|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|3354,3358|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|3354,3358|false|false|false|C0562271|Examination of knee joint|knee
Finding|Finding|General Exam|3354,3366|false|false|false|C0240114|Knee flexion|knee flexion
Attribute|Clinical Attribute|General Exam|3359,3366|false|false|false|C1525443|W flexion|flexion
Event|Event|General Exam|3359,3366|false|false|false|||flexion
Finding|Organ or Tissue Function|General Exam|3359,3366|false|false|false|C0231452||flexion
Event|Event|General Exam|3371,3380|false|false|false|||extension
Finding|Conceptual Entity|General Exam|3371,3380|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Finding|Functional Concept|General Exam|3371,3380|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Anatomy|Body Part, Organ, or Organ Component|General Exam|3382,3386|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|General Exam|3382,3386|false|false|false|C0555980|Foot problem|foot
Anatomy|Body Location or Region|General Exam|3387,3394|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|plantar
Event|Event|General Exam|3399,3411|false|false|false|||dorsiflexion
Event|Event|General Exam|3413,3422|false|false|false|||sensation
Finding|Finding|General Exam|3413,3422|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3413,3422|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3413,3422|false|false|false|C2229507|sensory exam|sensation
Drug|Amino Acid, Peptide, or Protein|General Exam|3426,3430|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Element, Ion, or Isotope|General Exam|3426,3430|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Immunologic Factor|General Exam|3426,3430|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Pharmacologic Substance|General Exam|3426,3430|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Finding|Idea or Concept|General Exam|3449,3454|false|false|false|C0812371|Ortho-|Ortho
Anatomy|Body Part, Organ, or Organ Component|General Exam|3455,3460|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|Spine
Anatomy|Cell Component|General Exam|3455,3460|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|Spine
Finding|Finding|General Exam|3455,3460|false|false|false|C0150920|Spine Problem|Spine
Event|Event|General Exam|3461,3465|false|false|false|||Exam
Finding|Functional Concept|General Exam|3461,3465|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|3461,3465|false|false|false|C0582103|Medical Examination|Exam
Event|Event|General Exam|3483,3487|false|false|false|||Temp
Finding|Gene or Genome|General Exam|3483,3487|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|3483,3487|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Individual Behavior|General Exam|3510,3515|false|false|false|C0600261|Telling untruths|Lying
Event|Event|General Exam|3516,3518|false|false|false|||HR
Event|Event|General Exam|3545,3553|false|false|false|||delivery
Finding|Finding|General Exam|3545,3553|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|3545,3553|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|3545,3553|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|3545,3553|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|3567,3571|false|false|false|||Temp
Finding|Gene or Genome|General Exam|3567,3571|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|3567,3571|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Individual Behavior|General Exam|3594,3599|false|false|false|C0600261|Telling untruths|Lying
Event|Event|General Exam|3600,3602|false|false|false|||HR
Event|Event|General Exam|3629,3637|false|false|false|||delivery
Finding|Finding|General Exam|3629,3637|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|3629,3637|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|3629,3637|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|3629,3637|false|false|false|C0011209|Obstetric Delivery|delivery
Disorder|Disease or Syndrome|General Exam|3644,3647|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3644,3647|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3644,3647|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3644,3647|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3644,3647|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|3644,3647|false|false|false|||NAD
Finding|Finding|General Exam|3644,3647|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|3649,3650|false|false|false|||A
Attribute|Clinical Attribute|General Exam|3658,3662|false|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|General Exam|3658,3662|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Attribute|Clinical Attribute|General Exam|3658,3669|false|false|false|C4050166||resp effort
Event|Event|General Exam|3663,3669|false|false|false|||effort
Finding|Organism Function|General Exam|3663,3669|false|false|false|C0015264|Exertion|effort
Event|Event|General Exam|3670,3673|false|false|false|||RRR
Drug|Amino Acid, Peptide, or Protein|General Exam|3753,3756|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Biologically Active Substance|General Exam|3753,3756|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Immunologic Factor|General Exam|3753,3756|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Finding|Gene or Genome|General Exam|3753,3756|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|lat
Anatomy|Body Part, Organ, or Organ Component|General Exam|3757,3760|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|3757,3760|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|General Exam|3757,3760|false|false|false|||arm
Finding|Gene or Genome|General Exam|3757,3760|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|3757,3760|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|3757,3760|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|3757,3760|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|General Exam|3764,3769|false|false|false|C0040067|Thumb structure|thumb
Anatomy|Body Part, Organ, or Organ Component|General Exam|3790,3796|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Disorder|Congenital Abnormality|General Exam|3800,3803|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|General Exam|3800,3803|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|General Exam|3800,3803|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Anatomy|Body Part, Organ, or Organ Component|General Exam|3804,3807|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|3804,3807|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|General Exam|3804,3807|false|false|false|||arm
Finding|Gene or Genome|General Exam|3804,3807|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|3804,3807|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|3804,3807|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|3804,3807|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|General Exam|3826,3830|false|false|false|||SILT
Event|Event|General Exam|3863,3867|false|false|false|||SILT
Event|Event|General Exam|3885,3889|false|false|false|||SILT
Event|Event|General Exam|3922,3926|false|false|false|||SILT
Anatomy|Body Location or Region|General Exam|3935,3940|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Body Part, Organ, or Organ Component|General Exam|3935,3940|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Cell Component|General Exam|3935,3940|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Body Location or Region|General Exam|4024,4029|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|Groin
Anatomy|Body Location or Region|General Exam|4032,4036|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|4032,4036|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|General Exam|4032,4036|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|General Exam|4032,4036|false|false|false|C0562271|Examination of knee joint|Knee
Disorder|Congenital Abnormality|General Exam|4039,4042|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|Med
Finding|Gene or Genome|General Exam|4039,4042|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Finding|Intellectual Product|General Exam|4039,4042|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Anatomy|Body Location or Region|General Exam|4043,4047|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|4043,4047|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|4050,4053|false|false|false|C0228547|Clava structure (body structure)|Grt
Anatomy|Body Part, Organ, or Organ Component|General Exam|4054,4057|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Part, Organ, or Organ Component|General Exam|4063,4066|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Location or Region|General Exam|4074,4079|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|Thigh
Event|Event|General Exam|4093,4097|false|false|false|||SILT
Event|Event|General Exam|4132,4136|false|false|false|||SILT
Event|Event|General Exam|4150,4154|false|false|false|||SILT
Event|Event|General Exam|4189,4193|false|false|false|||SILT
Event|Event|General Exam|4196,4201|false|false|false|||Motor
Finding|Functional Concept|General Exam|4196,4201|false|false|false|C1513492|motor movement|Motor
Finding|Gene or Genome|General Exam|4208,4211|false|false|false|C1413248;C3273706|CDAN1 gene;CDAN1 wt Allele|Dlt
Anatomy|Body Part, Organ, or Organ Component|General Exam|4216,4219|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|General Exam|4216,4219|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|General Exam|4216,4219|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|General Exam|4216,4219|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|General Exam|4216,4219|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|General Exam|4231,4234|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|4231,4234|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Event|Event|General Exam|4542,4550|false|false|false|||Reflexes
Finding|Finding|General Exam|4542,4550|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|General Exam|4542,4550|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|General Exam|4542,4550|false|false|false|C0436145|Examination of reflexes|Reflexes
Anatomy|Body Part, Organ, or Organ Component|General Exam|4556,4559|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|General Exam|4556,4559|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|General Exam|4556,4559|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|General Exam|4556,4559|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|General Exam|4556,4559|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|General Exam|4577,4580|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|4577,4580|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Disorder|Disease or Syndrome|General Exam|4588,4591|false|false|false|C0030587|Paroxysmal atrial tachycardia|Pat
Drug|Organic Chemical|General Exam|4588,4591|false|false|false|C2825250|Fenamole|Pat
Drug|Pharmacologic Substance|General Exam|4588,4591|false|false|false|C2825250|Fenamole|Pat
Event|Event|General Exam|4588,4591|false|false|false|||Pat
Finding|Molecular Function|General Exam|4588,4591|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|Pat
Procedure|Diagnostic Procedure|General Exam|4588,4591|false|false|false|C3897364|Thermoacoustic Computed Tomography|Pat
Disorder|Congenital Abnormality|General Exam|4599,4602|false|false|false|C0001080|Achondroplasia|Ach
Drug|Biologically Active Substance|General Exam|4599,4602|false|false|false|C0001041|acetylcholine|Ach
Drug|Organic Chemical|General Exam|4599,4602|false|false|false|C0001041|acetylcholine|Ach
Drug|Pharmacologic Substance|General Exam|4599,4602|false|false|false|C0001041|acetylcholine|Ach
Event|Event|General Exam|4599,4602|false|false|false|||Ach
Finding|Gene or Genome|General Exam|4599,4602|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Finding|Sign or Symptom|General Exam|4599,4602|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Event|Event|General Exam|4736,4744|false|false|false|||Negative
Finding|Classification|General Exam|4736,4744|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|General Exam|4736,4744|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|General Exam|4736,4744|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|General Exam|4745,4753|false|false|false|C0034935|Babinski Reflex|Babinski
Event|Event|General Exam|4766,4772|false|false|false|||Clonus
Finding|Sign or Symptom|General Exam|4766,4772|false|false|false|C0009024|Clonus|Clonus
Event|Event|General Exam|4805,4812|false|false|false|||IMAGING
Finding|Finding|General Exam|4805,4812|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4805,4812|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Attribute|Clinical Attribute|General Exam|4814,4831|false|false|false|C0882557||MR THORACIC SPINE
Anatomy|Body Location or Region|General Exam|4817,4825|false|false|false|C0817096|Chest|THORACIC
Disorder|Disease or Syndrome|General Exam|4817,4825|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|THORACIC
Anatomy|Body Part, Organ, or Organ Component|General Exam|4817,4831|false|false|false|C0581269|Thoracic spine structure|THORACIC SPINE
Anatomy|Body Part, Organ, or Organ Component|General Exam|4826,4831|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|SPINE
Anatomy|Cell Component|General Exam|4826,4831|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|SPINE
Finding|Finding|General Exam|4826,4831|false|false|false|C0150920|Spine Problem|SPINE
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4836,4844|false|true|false|C0009924|Contrast Media|CONTRAST
Anatomy|Body Part, Organ, or Organ Component|General Exam|4853,4858|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|SPINE
Anatomy|Cell Component|General Exam|4853,4858|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|SPINE
Finding|Finding|General Exam|4853,4858|false|false|false|C0150920|Spine Problem|SPINE
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4863,4871|false|false|false|C0009924|Contrast Media|CONTRAST
Finding|Finding|Impression|4891,4897|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Impression|4891,4897|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Pharmacologic Substance|Impression|4898,4905|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Impression|4898,4905|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Impression|4898,4905|false|false|false|||central
Procedure|Laboratory Procedure|Impression|4898,4905|false|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|Impression|4898,4911|false|false|false|C0459414|Central cord canal structure|central canal
Anatomy|Body Part, Organ, or Organ Component|Impression|4906,4911|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Anatomy|Body Space or Junction|Impression|4906,4911|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Disorder|Anatomical Abnormality|Impression|4912,4921|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|4912,4921|false|false|false|||narrowing
Finding|Functional Concept|Impression|4942,4954|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|Impression|4942,4954|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|Impression|4942,4962|false|false|false|C0011164|Abnormal degeneration|degenerative changes
Event|Event|Impression|4955,4962|false|false|false|||changes
Finding|Functional Concept|Impression|4955,4962|false|false|false|C0392747|Changing|changes
Finding|Gene or Genome|Impression|4967,4972|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|Large
Finding|Functional Concept|Impression|4973,4978|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|5000,5004|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|Impression|5000,5004|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|Impression|5000,5004|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|Impression|5000,5004|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|Impression|5000,5004|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Event|Event|Impression|5005,5014|false|false|false|||extrusion
Finding|Finding|Impression|5005,5014|false|false|false|C0443213|Extrusion|extrusion
Event|Event|Impression|5028,5035|false|false|false|||extends
Finding|Functional Concept|Impression|5041,5046|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Impression|5058,5064|false|false|false|||recess
Event|Event|Impression|5066,5070|false|false|false|||mass
Finding|Finding|Impression|5066,5070|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|5066,5070|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|5066,5070|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Impression|5066,5077|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|Impression|5071,5077|false|false|false|||effect
Event|Event|Impression|5081,5088|false|false|false|||exiting
Finding|Functional Concept|Impression|5089,5094|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|5114,5120|false|false|false|C0027740|Nerve|nerves
Finding|Finding|Impression|5122,5128|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Impression|5122,5128|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|Impression|5129,5134|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Anatomical Abnormality|Impression|5150,5159|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|5150,5159|false|false|false|||narrowing
Finding|Functional Concept|Impression|5174,5186|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|Impression|5174,5186|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|Impression|5174,5194|false|false|false|C0011164|Abnormal degeneration|degenerative changes
Event|Event|Impression|5187,5194|false|false|false|||changes
Finding|Functional Concept|Impression|5187,5194|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|Impression|5195,5201|false|false|false|C0024090|Lumbar Region|lumbar
Anatomy|Body Location or Region|Impression|5195,5207|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Impression|5195,5207|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Impression|5202,5207|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Impression|5202,5207|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Impression|5202,5207|false|false|false|C0150920|Spine Problem|spine
Finding|Finding|Impression|5212,5220|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Impression|5212,5220|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Pharmacologic Substance|Impression|5221,5228|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Impression|5221,5228|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Impression|5221,5228|false|false|false|||central
Procedure|Laboratory Procedure|Impression|5221,5228|false|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|Impression|5221,5234|false|false|false|C0459414|Central cord canal structure|central canal
Anatomy|Body Part, Organ, or Organ Component|Impression|5229,5234|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Anatomy|Body Space or Junction|Impression|5229,5234|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Disorder|Anatomical Abnormality|Impression|5235,5244|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|5235,5244|false|false|false|||narrowing
Event|Event|Impression|5252,5260|false|false|false|||moderate
Finding|Finding|Impression|5252,5260|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Impression|5252,5260|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|Impression|5264,5270|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Impression|5264,5270|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Impression|5281,5287|false|false|false|||levels
Finding|Idea or Concept|Impression|5303,5314|false|false|false|C0750502|Significant|significant
Disorder|Anatomical Abnormality|Impression|5325,5334|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|5325,5334|false|false|false|||narrowing
Anatomy|Body Location or Region|Impression|5335,5341|false|false|false|C0024090|Lumbar Region|lumbar
Anatomy|Body Location or Region|Impression|5335,5347|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Impression|5335,5347|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Impression|5342,5347|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Impression|5342,5347|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Impression|5342,5347|false|false|false|C0150920|Spine Problem|spine
Finding|Idea or Concept|Impression|5353,5358|false|false|false|C1552828|Table Frame - above|above
Finding|Functional Concept|Impression|5363,5375|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degenerative
Finding|Pathologic Function|Impression|5363,5375|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degenerative
Finding|Pathologic Function|Impression|5363,5383|false|false|false|C0011164|Abnormal degeneration|Degenerative changes
Event|Event|Impression|5376,5383|false|false|false|||changes
Finding|Functional Concept|Impression|5376,5383|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|Impression|5384,5392|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Impression|5384,5392|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|Impression|5384,5398|false|false|false|C0581269|Thoracic spine structure|thoracic spine
Anatomy|Body Part, Organ, or Organ Component|Impression|5393,5398|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Impression|5393,5398|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Impression|5393,5398|false|false|false|C0150920|Spine Problem|spine
Finding|Intellectual Product|Impression|5400,5404|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Impression|5408,5416|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Impression|5408,5416|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Drug|Pharmacologic Substance|Impression|5417,5424|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Impression|5417,5424|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Impression|5417,5424|false|false|false|||central
Procedure|Laboratory Procedure|Impression|5417,5424|false|false|false|C1879652|Central Minus|central
Anatomy|Body Part, Organ, or Organ Component|Impression|5426,5431|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Anatomy|Body Space or Junction|Impression|5426,5431|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Disorder|Anatomical Abnormality|Impression|5432,5441|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|5432,5441|false|false|false|||narrowing
Disorder|Anatomical Abnormality|Impression|5453,5462|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Impression|5453,5462|false|false|false|||narrowing
Attribute|Clinical Attribute|Impression|5465,5471|false|false|false|C1644645||CT ABD
Anatomy|Body Location or Region|Impression|5468,5471|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|Impression|5468,5471|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|Impression|5468,5471|false|false|false|||ABD
Anatomy|Body Part, Organ, or Organ Component|Impression|5474,5480|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|Impression|5474,5480|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|Impression|5474,5480|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|Impression|5474,5480|false|false|false|||PELVIS
Finding|Finding|Impression|5474,5480|false|false|false|C0812455|Pelvis problem|PELVIS
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5486,5494|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|Impression|5486,5494|false|false|false|||CONTRAST
Finding|Intellectual Product|Impression|5519,5524|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|Impression|5528,5536|false|false|false|C2926606||findings
Event|Event|Impression|5528,5536|false|false|false|||findings
Finding|Functional Concept|Impression|5528,5536|false|false|false|C2607943|findings aspects|findings
Anatomy|Body Location or Region|Impression|5544,5551|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Impression|5544,5551|true|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Impression|5544,5551|true|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|Impression|5555,5561|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Impression|5555,5561|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Impression|5555,5561|true|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|Impression|5555,5561|false|false|false|||pelvis
Finding|Finding|Impression|5555,5561|true|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Impression|5565,5574|false|false|false|||correlate
Finding|Body Substance|Impression|5581,5588|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|5581,5588|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|5581,5588|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|5600,5608|false|false|false|||symptoms
Finding|Functional Concept|Impression|5600,5608|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Impression|5600,5608|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Impression|5628,5636|false|false|false|||evidence
Finding|Idea or Concept|Impression|5628,5636|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5628,5639|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Impression|5640,5651|false|false|false|||obstructive
Finding|Functional Concept|Impression|5640,5651|true|false|false|C0549186|Obstructed|obstructive
Anatomy|Body Part, Organ, or Organ Component|Impression|5653,5658|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Impression|5653,5658|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Impression|5653,5664|false|false|false|C0392525|Nephrolithiasis|renal stone
Finding|Body Substance|Impression|5653,5664|false|false|false|C0022650;C1458136|Kidney Calculi;Renal stone (substance)|renal stone
Event|Event|Impression|5659,5664|false|false|false|||stone
Finding|Body Substance|Impression|5659,5664|false|false|false|C0006736|Calculi|stone
Disorder|Disease or Syndrome|Impression|5668,5682|false|false|false|C0034186|Pyelonephritis|pyelonephritis
Event|Event|Impression|5668,5682|false|false|false|||pyelonephritis
Anatomy|Body Part, Organ, or Organ Component|Impression|5687,5694|false|false|false|C0227391|Sigmoid colon|Sigmoid
Disorder|Disease or Syndrome|Impression|5687,5709|false|false|false|C0012818|Diverticulosis of sigmoid colon|Sigmoid diverticulosis
Disorder|Disease or Syndrome|Impression|5695,5709|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|Impression|5695,5709|false|false|false|||diverticulosis
Event|Event|Impression|5720,5728|false|false|false|||evidence
Finding|Idea or Concept|Impression|5720,5728|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5720,5731|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Impression|5732,5737|false|false|false|||acute
Finding|Intellectual Product|Impression|5732,5737|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Impression|5739,5753|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|Impression|5739,5753|false|false|false|||diverticulitis
Procedure|Health Care Activity|Impression|5756,5765|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Impression|5766,5770|false|false|false|||Labs
Lab|Laboratory or Test Result|Impression|5766,5770|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|Impression|5784,5789|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|5784,5789|false|false|false|||BLOOD
Finding|Body Substance|Impression|5784,5789|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|5790,5793|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|5798,5801|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|5798,5801|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|5798,5801|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|5807,5810|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|5807,5810|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|5807,5810|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|5807,5810|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|5816,5819|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|5816,5819|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|5825,5828|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Impression|5825,5828|false|false|false|||MCV
Lab|Laboratory or Test Result|Impression|5825,5828|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|5825,5828|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|5825,5828|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|5833,5836|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|5833,5836|false|false|false|C0600370|methacholine|MCH
Event|Event|Impression|5833,5836|false|false|false|||MCH
Finding|Gene or Genome|Impression|5833,5836|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|5833,5836|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|5833,5836|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Impression|5842,5846|false|false|false|||MCHC
Procedure|Laboratory Procedure|Impression|5842,5846|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|5873,5876|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|5893,5898|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|5893,5898|false|false|false|||BLOOD
Finding|Body Substance|Impression|5893,5898|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Impression|5903,5906|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Impression|5903,5906|false|false|false|||PTT
Procedure|Laboratory Procedure|Impression|5903,5906|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Impression|5928,5933|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|5928,5933|false|false|false|||BLOOD
Finding|Body Substance|Impression|5928,5933|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|5928,5941|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|5928,5941|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|5928,5941|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|5934,5941|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|5934,5941|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|5934,5941|false|false|false|C0017725|glucose|Glucose
Event|Event|Impression|5934,5941|false|false|false|||Glucose
Lab|Laboratory or Test Result|Impression|5934,5941|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|5934,5941|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|5987,5991|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|5987,5991|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|5987,5991|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6017,6022|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6017,6022|false|false|false|||BLOOD
Finding|Body Substance|Impression|6017,6022|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|6023,6026|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|6031,6034|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|6031,6034|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|6031,6034|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|6041,6044|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|6041,6044|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|6041,6044|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|6041,6044|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|6050,6053|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|6050,6053|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|6061,6064|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Impression|6061,6064|false|false|false|||MCV
Lab|Laboratory or Test Result|Impression|6061,6064|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|6061,6064|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|6061,6064|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|6068,6071|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|6068,6071|false|false|false|C0600370|methacholine|MCH
Event|Event|Impression|6068,6071|false|false|false|||MCH
Finding|Gene or Genome|Impression|6068,6071|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|6068,6071|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|6068,6071|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Impression|6077,6081|false|false|false|||MCHC
Procedure|Laboratory Procedure|Impression|6077,6081|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|6108,6111|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|6128,6133|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6128,6133|false|false|false|||BLOOD
Finding|Body Substance|Impression|6128,6133|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|6134,6137|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|6142,6145|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|6142,6145|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|6142,6145|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|6152,6155|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|6152,6155|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|6152,6155|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|6152,6155|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|6161,6164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|6161,6164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|6172,6175|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Impression|6172,6175|false|false|false|||MCV
Lab|Laboratory or Test Result|Impression|6172,6175|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|6172,6175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|6172,6175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|6179,6182|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|6179,6182|false|false|false|C0600370|methacholine|MCH
Event|Event|Impression|6179,6182|false|false|false|||MCH
Finding|Gene or Genome|Impression|6179,6182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|6179,6182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|6179,6182|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Impression|6188,6192|false|false|false|||MCHC
Procedure|Laboratory Procedure|Impression|6188,6192|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|6219,6222|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|6239,6244|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6239,6244|false|false|false|||BLOOD
Finding|Body Substance|Impression|6239,6244|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|6245,6248|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|6253,6256|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|6253,6256|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|6253,6256|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|6263,6266|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|6263,6266|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|6263,6266|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|6263,6266|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|6273,6276|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|6273,6276|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|6284,6287|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Impression|6284,6287|false|false|false|||MCV
Lab|Laboratory or Test Result|Impression|6284,6287|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|6284,6287|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|6284,6287|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|6291,6294|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|6291,6294|false|false|false|C0600370|methacholine|MCH
Event|Event|Impression|6291,6294|false|false|false|||MCH
Finding|Gene or Genome|Impression|6291,6294|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|6291,6294|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|6291,6294|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Impression|6300,6304|false|false|false|||MCHC
Procedure|Laboratory Procedure|Impression|6300,6304|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|6332,6335|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|6352,6357|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|6352,6357|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|6358,6361|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|6378,6383|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6378,6383|false|false|false|||BLOOD
Finding|Body Substance|Impression|6378,6383|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|6378,6391|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|6378,6391|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|6378,6391|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|6384,6391|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|6384,6391|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|6384,6391|false|false|false|C0017725|glucose|Glucose
Event|Event|Impression|6384,6391|false|false|false|||Glucose
Lab|Laboratory or Test Result|Impression|6384,6391|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|6384,6391|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|6437,6441|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|6437,6441|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|6437,6441|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6466,6471|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6466,6471|false|false|false|||BLOOD
Finding|Body Substance|Impression|6466,6471|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|6466,6479|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|6466,6479|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|6466,6479|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|6472,6479|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|6472,6479|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|6472,6479|false|false|false|C0017725|glucose|Glucose
Event|Event|Impression|6472,6479|false|false|false|||Glucose
Lab|Laboratory or Test Result|Impression|6472,6479|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|6472,6479|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|6524,6528|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|6524,6528|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|6524,6528|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6553,6558|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6553,6558|false|false|false|||BLOOD
Finding|Body Substance|Impression|6553,6558|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|6553,6566|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|6553,6566|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|6553,6566|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|6559,6566|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|6559,6566|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|6559,6566|false|false|false|C0017725|glucose|Glucose
Event|Event|Impression|6559,6566|false|false|false|||Glucose
Lab|Laboratory or Test Result|Impression|6559,6566|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|6559,6566|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|6612,6616|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|6612,6616|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|6612,6616|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6641,6646|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6641,6646|false|false|false|||BLOOD
Finding|Body Substance|Impression|6641,6646|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|6641,6654|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|6647,6654|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|6647,6654|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|6647,6654|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|6647,6654|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|6647,6654|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Impression|6647,6654|false|false|false|||Calcium
Finding|Physiologic Function|Impression|6647,6654|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|6647,6654|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|Impression|6688,6693|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6688,6693|false|false|false|||BLOOD
Finding|Body Substance|Impression|6688,6693|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|6688,6701|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|6694,6701|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|6694,6701|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|6694,6701|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|6694,6701|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|6694,6701|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Impression|6694,6701|false|false|false|||Calcium
Finding|Physiologic Function|Impression|6694,6701|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|6694,6701|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|Impression|6734,6739|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6734,6739|false|false|false|||BLOOD
Finding|Body Substance|Impression|6734,6739|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|6734,6747|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|6740,6747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|6740,6747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|6740,6747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|6740,6747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|6740,6747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Impression|6740,6747|false|false|false|||Calcium
Finding|Physiologic Function|Impression|6740,6747|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|6740,6747|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Idea or Concept|Hospital Course|6794,6801|false|false|false|C1555582|Initial (abbreviation)|Initial
Event|Event|Hospital Course|6802,6811|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|6802,6811|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Hospital Course|6821,6827|false|false|false|||ISSUES
Finding|Finding|Hospital Course|6852,6855|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Hospital Course|6852,6855|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Sign or Symptom|Hospital Course|6852,6865|false|false|false|C0024031|Low Back Pain|Low Back pain
Finding|Sign or Symptom|Hospital Course|6856,6865|false|true|false|C0004604|Back Pain|Back pain
Attribute|Clinical Attribute|Hospital Course|6861,6865|false|false|false|C2598155||pain
Event|Event|Hospital Course|6861,6865|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6861,6865|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6861,6865|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6870,6873|false|false|false|C0023216;C1140621|Leg;Lower Extremity|Leg
Finding|Sign or Symptom|Hospital Course|6870,6878|false|true|false|C0023222|Pain in lower limb|Leg Pain
Attribute|Clinical Attribute|Hospital Course|6874,6878|false|false|false|C2598155||Pain
Event|Event|Hospital Course|6874,6878|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|6874,6878|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|6874,6878|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|Hospital Course|6881,6894|false|false|false|C0700594|Radiculopathy|Radiculopathy
Event|Event|Hospital Course|6881,6894|false|false|false|||Radiculopathy
Finding|Body Substance|Hospital Course|6895,6902|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6895,6902|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6895,6902|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6903,6911|false|false|false|||presents
Finding|Finding|Hospital Course|6917,6923|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6917,6923|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|Hospital Course|6924,6929|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Sign or Symptom|Hospital Course|6924,6945|false|true|false|C2219286|right-sided low back pain|right lower back pain
Anatomy|Body Location or Region|Hospital Course|6930,6935|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|6930,6935|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|Hospital Course|6930,6940|false|false|false|C0230102;C2939142|Lower back (surface region);Lower back structure|lower back
Finding|Sign or Symptom|Hospital Course|6930,6945|false|true|false|C0024031|Low Back Pain|lower back pain
Finding|Sign or Symptom|Hospital Course|6936,6945|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Hospital Course|6941,6945|false|true|false|C2598155||pain
Event|Event|Hospital Course|6941,6945|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6941,6945|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6941,6945|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6962,6973|false|false|false|||lancinating
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6974,6983|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|6974,6983|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|6974,6983|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|6974,6983|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|6974,6983|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|6974,6983|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6985,6989|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Drug|Enzyme|Hospital Course|6985,6989|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Event|Event|Hospital Course|6988,6989|false|false|false|||A
Event|Event|Hospital Course|7000,7008|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|7000,7008|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|7000,7011|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Hospital Course|7012,7020|false|false|false|||visceral
Event|Event|Hospital Course|7021,7030|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|7021,7030|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|7021,7030|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|7021,7030|false|false|false|C0919386|Pathology procedure|pathology
Disorder|Disease or Syndrome|Hospital Course|7034,7049|false|false|false|C0392525|Nephrolithiasis|nephrolithiasis
Event|Event|Hospital Course|7034,7049|false|false|false|||nephrolithiasis
Event|Event|Hospital Course|7051,7054|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|7051,7054|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|7051,7054|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|7051,7054|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Location or Region|Hospital Course|7055,7062|false|false|false|C3887615|Lumbar spine structure|L spine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7057,7062|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Hospital Course|7057,7062|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Hospital Course|7057,7062|false|false|false|C0150920|Spine Problem|spine
Finding|Idea or Concept|Hospital Course|7068,7079|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7080,7084|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|Hospital Course|7080,7084|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|Hospital Course|7080,7084|false|false|false|C0993608|Disk Drug Form|disc
Event|Event|Hospital Course|7080,7084|false|false|false|||disc
Finding|Finding|Hospital Course|7080,7084|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|Hospital Course|7080,7084|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Event|Event|Hospital Course|7085,7090|false|false|false|||bulge
Finding|Finding|Hospital Course|7085,7090|false|false|false|C0038999|Swelling|bulge
Event|Event|Hospital Course|7109,7114|false|false|false|||cause
Finding|Conceptual Entity|Hospital Course|7109,7114|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Hospital Course|7109,7114|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Finding|Hospital Course|7115,7121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|7115,7121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Anatomical Abnormality|Hospital Course|7122,7131|false|false|false|C3854333|Narrowing|narrowing
Event|Event|Hospital Course|7122,7131|false|false|false|||narrowing
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7146,7151|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Anatomy|Body Space or Junction|Hospital Course|7146,7151|false|false|false|C0086881;C1550227|Pulp Canals;canal [body parts]|canal
Event|Event|Hospital Course|7156,7165|false|false|false|||extrusion
Finding|Finding|Hospital Course|7156,7165|false|false|false|C0443213|Extrusion|extrusion
Finding|Idea or Concept|Hospital Course|7179,7190|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7191,7199|false|false|false|C0501792|Fourth lumbar nerve|L4 nerve
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7194,7199|false|false|false|C0027740|Nerve|nerve
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7194,7204|false|false|false|C0228084|Nerve root structure|nerve root
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7200,7204|false|false|false|C0040452;C1318154|Root body part;Tooth root structure|root
Finding|Idea or Concept|Hospital Course|7200,7204|false|false|false|C1705917|Tree Root (hierarchy)|root
Event|Event|Hospital Course|7205,7216|false|false|false|||compression
Finding|Functional Concept|Hospital Course|7205,7216|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|7205,7216|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|7205,7216|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7205,7216|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Finding|Hospital Course|7218,7224|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|7218,7224|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|7229,7234|false|false|false|||cause
Finding|Conceptual Entity|Hospital Course|7229,7234|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Hospital Course|7229,7234|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Body Substance|Hospital Course|7238,7245|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7238,7245|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7238,7245|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|7248,7252|false|false|false|C2598155||pain
Event|Event|Hospital Course|7248,7252|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7248,7252|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7248,7252|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|7272,7280|false|false|false|||admitted
Finding|Functional Concept|Hospital Course|7286,7291|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7286,7295|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Finding|Sign or Symptom|Hospital Course|7286,7300|false|false|false|C5848135|Pain in right leg|right leg pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7292,7295|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|7292,7300|false|false|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Hospital Course|7296,7300|false|false|false|C2598155||pain
Event|Event|Hospital Course|7296,7300|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7296,7300|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7296,7300|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|7307,7311|false|false|false|||exam
Finding|Functional Concept|Hospital Course|7307,7311|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|7307,7311|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|7312,7319|false|false|false|||notable
Event|Event|Hospital Course|7324,7336|false|false|false|||trochanteric
Disorder|Disease or Syndrome|Hospital Course|7337,7345|false|false|false|C0006444|Bursitis|bursitis
Event|Event|Hospital Course|7337,7345|false|false|false|||bursitis
Drug|Biomedical or Dental Material|Hospital Course|7355,7364|false|false|false|C1272883|Injection|injection
Event|Event|Hospital Course|7355,7364|false|false|false|||injection
Finding|Functional Concept|Hospital Course|7355,7364|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7355,7364|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Drug|Hormone|Hospital Course|7368,7382|false|false|false|C0001617;C3536709|Adrenal Cortex Hormones;Corticosteroid [EPC]|corticosteroid
Drug|Organic Chemical|Hospital Course|7368,7382|false|false|false|C0001617;C3536709|Adrenal Cortex Hormones;Corticosteroid [EPC]|corticosteroid
Drug|Pharmacologic Substance|Hospital Course|7368,7382|false|false|false|C0001617;C3536709|Adrenal Cortex Hormones;Corticosteroid [EPC]|corticosteroid
Event|Event|Hospital Course|7368,7382|false|false|false|||corticosteroid
Event|Event|Hospital Course|7410,7416|false|false|false|||intact
Finding|Finding|Hospital Course|7410,7416|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|Hospital Course|7426,7434|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|7426,7434|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|7426,7437|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7438,7442|false|false|false|C1550235|Cord - Body Parts|cord
Disorder|Disease or Syndrome|Hospital Course|7438,7442|false|false|false|C3489532|Cone-Rod Dystrophy 2|cord
Disorder|Disease or Syndrome|Hospital Course|7438,7454|true|false|false|C0037926;C0266798|Compression of spinal cord;Compression of umbilical cord|cord compression
Event|Event|Hospital Course|7443,7454|false|false|false|||compression
Finding|Functional Concept|Hospital Course|7443,7454|true|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|7443,7454|true|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|7443,7454|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7443,7454|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|Hospital Course|7458,7465|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|7458,7465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7458,7465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7458,7465|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|Hospital Course|7472,7476|false|false|false|||exam
Finding|Functional Concept|Hospital Course|7472,7476|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|7472,7476|false|false|false|C0582103|Medical Examination|exam
Finding|Idea or Concept|Hospital Course|7482,7487|false|false|false|C0812371|Ortho-|ortho
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7488,7493|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Hospital Course|7488,7493|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Hospital Course|7488,7493|false|false|false|C0150920|Spine Problem|spine
Event|Event|Hospital Course|7501,7508|false|false|false|||benefit
Event|Event|Hospital Course|7514,7527|false|false|false|||decompression
Finding|Functional Concept|Hospital Course|7514,7527|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|Hospital Course|7514,7527|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7514,7527|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Event|Event|Hospital Course|7539,7552|false|false|false|||DECOMPRESSION
Finding|Functional Concept|Hospital Course|7539,7552|false|false|false|C1965697|Decompression - action (qualifier value)|DECOMPRESSION
Phenomenon|Phenomenon or Process|Hospital Course|7539,7552|false|false|false|C0011117|external decompression|DECOMPRESSION
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7539,7552|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|DECOMPRESSION
Event|Event|Hospital Course|7560,7566|false|false|false|||FUSION
Finding|Functional Concept|Hospital Course|7560,7566|false|false|false|C0332466|Fused structure|FUSION
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7560,7566|false|false|false|C1293131|Fusion procedure|FUSION
Event|Event|Hospital Course|7575,7585|false|false|false|||DURAPLASTY
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7575,7585|false|false|false|C0546551|Duraplasty|DURAPLASTY
Attribute|Clinical Attribute|Hospital Course|7617,7620|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|Hospital Course|7617,7620|false|false|false|||INR
Procedure|Laboratory Procedure|Hospital Course|7617,7620|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7617,7620|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|Hospital Course|7639,7646|false|false|false|||started
Drug|Biologically Active Substance|Hospital Course|7652,7659|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7652,7659|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|7652,7659|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|7660,7666|false|false|false|||bridge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7660,7666|false|false|false|C0399080|Fixation of dental bridge|bridge
Attribute|Clinical Attribute|Hospital Course|7683,7686|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|Hospital Course|7683,7686|false|false|false|||INR
Procedure|Laboratory Procedure|Hospital Course|7683,7686|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7683,7686|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|Hospital Course|7687,7694|false|false|false|||dropped
Event|Event|Hospital Course|7710,7722|false|false|false|||transitioned
Drug|Organic Chemical|Hospital Course|7726,7733|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|7726,7733|false|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|7734,7740|false|false|false|||bridge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7734,7740|false|false|false|C0399080|Fixation of dental bridge|bridge
Drug|Organic Chemical|Hospital Course|7744,7752|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|7744,7752|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Hospital Course|7744,7752|false|false|false|||coumadin
Event|Event|Hospital Course|7764,7771|false|false|false|||Dysuria
Finding|Sign or Symptom|Hospital Course|7764,7771|false|false|false|C0013428|Dysuria|Dysuria
Event|Event|Hospital Course|7773,7781|false|false|false|||resolved
Disorder|Disease or Syndrome|Hospital Course|7785,7788|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7785,7788|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|7785,7788|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|7785,7788|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|7785,7788|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|Hospital Course|7789,7795|false|false|false|||States
Finding|Sign or Symptom|Hospital Course|7816,7823|false|false|false|C0085624|Burning sensation|burning
Finding|Sign or Symptom|Hospital Course|7816,7828|false|false|false|C0234230|Pain, Burning|burning pain
Attribute|Clinical Attribute|Hospital Course|7824,7828|false|false|false|C2598155||pain
Event|Event|Hospital Course|7824,7828|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7824,7828|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7824,7828|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7824,7843|false|false|false|C0013428|Dysuria|pain with urination
Event|Event|Hospital Course|7834,7843|false|false|false|||urination
Finding|Organism Function|Hospital Course|7834,7843|false|false|false|C0042034|Urination|urination
Event|Event|Hospital Course|7863,7868|false|false|false|||feels
Event|Event|Hospital Course|7878,7883|false|false|false|||needs
Event|Event|Hospital Course|7887,7891|false|false|false|||push
Anatomy|Body Location or Region|Hospital Course|7899,7906|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|7899,7906|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|7899,7906|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|Hospital Course|7910,7917|false|false|false|||urinate
Event|Event|Hospital Course|7924,7934|false|false|false|||concerning
Disorder|Disease or Syndrome|Hospital Course|7939,7942|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7939,7942|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|7939,7942|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|7939,7942|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|7939,7942|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|Hospital Course|7947,7960|false|false|false|||demonstrating
Finding|Gene or Genome|Hospital Course|7961,7966|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Cell|Hospital Course|7967,7977|false|false|false|C0023516|Leukocytes|leukocytes
Finding|Body Substance|Hospital Course|7967,7977|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Finding|Intellectual Product|Hospital Course|7967,7977|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Anatomy|Cell|Hospital Course|7984,7987|false|false|false|C0023516|Leukocytes|WBC
Finding|Body Substance|Hospital Course|7998,8003|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|7998,8003|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|7998,8003|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Procedure|Laboratory Procedure|Hospital Course|7998,8011|false|false|false|C0430404|Urine culture|urine culture
Drug|Biomedical or Dental Material|Hospital Course|8004,8011|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|8004,8011|false|false|false|||culture
Finding|Functional Concept|Hospital Course|8004,8011|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|8004,8011|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|8004,8011|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|Hospital Course|8012,8019|false|false|false|||showing
Event|Event|Hospital Course|8042,8052|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|8042,8052|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|8042,8057|false|false|false|C0332290|Consistent with|consistent with
Event|Event|Hospital Course|8058,8071|false|false|false|||contamination
Finding|Idea or Concept|Hospital Course|8058,8071|false|false|false|C2349974|Contamination|contamination
Phenomenon|Human-caused Phenomenon or Process|Hospital Course|8058,8071|false|false|false|C0259846|adulteration|contamination
Event|Event|Hospital Course|8078,8083|false|false|false|||treat
Event|Event|Hospital Course|8090,8098|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|8090,8098|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|8090,8098|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body Location or Region|Hospital Course|8100,8109|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Hospital Course|8100,8114|false|true|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Hospital Course|8110,8114|false|true|false|C2598155||pain
Event|Event|Hospital Course|8110,8114|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8110,8114|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8110,8114|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8134,8146|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|8134,8146|false|true|false|C0009806|Constipation|constipation
Finding|Mental Process|Hospital Course|8154,8161|false|false|false|C0542559|contextual factors|setting
Drug|Hazardous or Poisonous Substance|Hospital Course|8165,8171|false|false|false|C0242402|Opioids|opioid
Drug|Organic Chemical|Hospital Course|8165,8171|false|false|false|C0242402|Opioids|opioid
Drug|Pharmacologic Substance|Hospital Course|8165,8171|false|false|false|C0242402|Opioids|opioid
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8165,8175|false|false|false|C0240602|opioid use|opioid use
Event|Event|Hospital Course|8172,8175|false|false|false|||use
Finding|Functional Concept|Hospital Course|8172,8175|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|8172,8175|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Hospital Course|8177,8184|false|false|false|||Reports
Finding|Intellectual Product|Hospital Course|8177,8184|false|false|false|C0684224|Report (document)|Reports
Procedure|Health Care Activity|Hospital Course|8177,8184|false|false|false|C0700287|Reporting|Reports
Event|Event|Hospital Course|8185,8195|false|false|false|||resolution
Finding|Conceptual Entity|Hospital Course|8185,8195|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|8185,8195|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Event|Event|Hospital Course|8199,8207|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|8199,8207|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|8199,8207|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|8220,8227|false|false|false|||treated
Drug|Organic Chemical|Hospital Course|8234,8241|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|Hospital Course|8234,8241|false|false|false|C0591139|Bactrim|bactrim
Event|Event|Hospital Course|8234,8241|false|false|false|||bactrim
Drug|Organic Chemical|Hospital Course|8234,8244|false|false|false|C1154231|Bactrim DS|bactrim DS
Drug|Pharmacologic Substance|Hospital Course|8234,8244|false|false|false|C1154231|Bactrim DS|bactrim DS
Event|Event|Hospital Course|8242,8244|false|false|false|||DS
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8245,8248|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8245,8248|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8245,8248|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8245,8248|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8245,8248|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|8260,8268|false|false|false|||starting
Event|Event|Hospital Course|8291,8298|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|8291,8298|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|8291,8298|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Event|Event|Hospital Course|8329,8336|false|false|false|||History
Finding|Conceptual Entity|Hospital Course|8329,8336|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|8329,8336|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|8329,8336|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|8329,8339|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|8340,8343|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|8340,8343|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|8340,8343|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|8340,8343|false|false|false|||DVT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8349,8374|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Drug|Immunologic Factor|Hospital Course|8349,8374|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Finding|Finding|Hospital Course|8349,8374|false|false|false|C4019436|Antiphospholipid antibody positivity|Antiphospholipid antibody
Disorder|Disease or Syndrome|Hospital Course|8349,8383|false|false|false|C0085278|Antiphospholipid Syndrome|Antiphospholipid antibody syndrome
Anatomy|Cell Component|Hospital Course|8366,8374|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8366,8374|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Hospital Course|8366,8374|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Hospital Course|8366,8374|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Hospital Course|8366,8374|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Hospital Course|8375,8383|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|8375,8383|false|false|false|||syndrome
Disorder|Disease or Syndrome|Hospital Course|8385,8390|false|false|false|C0024131;C0024138;C0024141;C0409974;C5574816|Chronic discoid lupus erythematosus;Discoid lupus erythematosus;Lupus Erythematosus;Lupus Erythematosus, Systemic;Lupus Vulgaris|Lupus
Disorder|Disease or Syndrome|Hospital Course|8385,8404|false|false|false|C0311370|Lupus anticoagulant disorder|Lupus anticoagulant
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8385,8404|false|false|false|C0085240|Lupus Coagulation Inhibitor|Lupus anticoagulant
Drug|Immunologic Factor|Hospital Course|8385,8404|false|false|false|C0085240|Lupus Coagulation Inhibitor|Lupus anticoagulant
Finding|Finding|Hospital Course|8385,8404|false|false|false|C4321325||Lupus anticoagulant
Procedure|Laboratory Procedure|Hospital Course|8385,8404|false|false|false|C1142517|Lupus anticoagulant assay|Lupus anticoagulant
Lab|Laboratory or Test Result|Hospital Course|8385,8413|false|false|false|C1142516|Lupus anticoagulant positive|Lupus anticoagulant positive
Drug|Pharmacologic Substance|Hospital Course|8391,8404|false|false|false|C0003280;C3536711|Anti-coagulant [EPC];Anticoagulants|anticoagulant
Event|Event|Hospital Course|8391,8404|false|false|false|||anticoagulant
Event|Event|Hospital Course|8460,8466|false|false|false|||taking
Finding|Idea or Concept|Hospital Course|8471,8475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8471,8475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8471,8475|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8476,8480|false|false|false|||dose
Drug|Hazardous or Poisonous Substance|Hospital Course|8484,8492|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|8484,8492|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|8484,8492|false|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|8484,8492|false|false|false|||warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|8528,8536|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|8528,8536|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|8528,8536|false|false|false|C0043031|warfarin|Warfarin
Event|Event|Hospital Course|8537,8541|false|false|false|||held
Event|Event|Hospital Course|8545,8554|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8545,8554|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Attribute|Clinical Attribute|Hospital Course|8559,8568|false|false|false|C0945766||procedure
Event|Event|Hospital Course|8559,8568|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|8559,8568|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|8559,8568|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8559,8568|false|false|false|C0184661|Interventional procedure|procedure
Drug|Biologically Active Substance|Hospital Course|8575,8582|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8575,8582|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8575,8582|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|8583,8587|false|false|false|||drip
Attribute|Clinical Attribute|Hospital Course|8594,8603|false|false|false|C0945766||procedure
Event|Event|Hospital Course|8594,8603|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|8594,8603|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|8594,8603|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8594,8603|false|false|false|C0184661|Interventional procedure|procedure
Disorder|Anatomical Abnormality|Hospital Course|8609,8612|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Hospital Course|8609,8612|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8609,8612|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Hospital Course|8609,8612|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Hospital Course|8609,8612|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Hospital Course|8609,8612|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|Hospital Course|8609,8612|false|false|false|||AAA
Finding|Gene or Genome|Hospital Course|8609,8612|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|Hospital Course|8628,8635|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|8628,8635|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8628,8635|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|8628,8635|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8628,8638|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|Hospital Course|8639,8642|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Hospital Course|8639,8642|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8639,8642|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Hospital Course|8639,8642|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Hospital Course|8639,8642|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Hospital Course|8639,8642|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|Hospital Course|8639,8642|false|false|false|||AAA
Finding|Gene or Genome|Hospital Course|8639,8642|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|Hospital Course|8646,8651|false|false|false|||chart
Finding|Intellectual Product|Hospital Course|8646,8651|false|false|false|C0684240|Charts (publication)|chart
Event|Event|Hospital Course|8666,8672|false|false|false|||follow
Event|Event|Hospital Course|8692,8704|false|false|false|||surveillance
Event|Occupational Activity|Hospital Course|8692,8704|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|Hospital Course|8692,8704|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|Hospital Course|8692,8704|false|false|false|C0733511|Medical Surveillance|surveillance
Attribute|Clinical Attribute|Hospital Course|8709,8715|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|Hospital Course|8712,8715|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|Hospital Course|8712,8715|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8716,8722|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|8716,8722|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|8716,8722|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|8716,8722|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|Hospital Course|8731,8735|false|false|false|||show
Anatomy|Body Location or Region|Hospital Course|8739,8748|false|false|false|C0000726|Abdomen|abdominal
Attribute|Clinical Attribute|Hospital Course|8739,8764|false|false|false|C2926614||abdominal aortic aneurysm
Disorder|Anatomical Abnormality|Hospital Course|8739,8764|false|false|false|C0162871|Aortic Aneurysm, Abdominal|abdominal aortic aneurysm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8749,8755|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|Hospital Course|8749,8764|false|false|false|C0003486;C0340629|Aortic Aneurysm|aortic aneurysm
Event|Event|Hospital Course|8756,8764|false|false|false|||aneurysm
Finding|Pathologic Function|Hospital Course|8756,8764|false|false|false|C0002940|Aneurysm|aneurysm
Drug|Organic Chemical|Hospital Course|8769,8776|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|8769,8776|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|8769,8776|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|8769,8778|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|8769,8778|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|8769,8778|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|8769,8778|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|8769,8778|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Disorder|Disease or Syndrome|Hospital Course|8769,8789|false|false|false|C0042870|Vitamin D Deficiency|Vitamin D deficiency
Finding|Finding|Hospital Course|8769,8789|false|false|false|C5886864|Decreased circulating vitamin D concentration|Vitamin D deficiency
Disorder|Disease or Syndrome|Hospital Course|8779,8789|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Hospital Course|8779,8789|false|false|false|||deficiency
Finding|Functional Concept|Hospital Course|8779,8789|false|false|false|C0011155|Deficiency|deficiency
Event|Event|Hospital Course|8793,8802|false|false|false|||Continued
Drug|Organic Chemical|Hospital Course|8803,8810|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|8803,8810|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|8803,8810|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|8803,8812|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|8803,8812|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|8803,8812|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|8803,8812|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|8803,8812|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|8811,8812|false|false|false|||D
Disorder|Disease or Syndrome|Hospital Course|8826,8829|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8826,8829|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Hospital Course|8826,8829|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|Hospital Course|8826,8829|false|false|false|||OSA
Event|Event|Hospital Course|8832,8840|false|false|false|||Remained
Event|Event|Hospital Course|8844,8848|false|false|false|||CPAP
Finding|Gene or Genome|Hospital Course|8844,8848|false|false|false|C1424863|CENPJ gene|CPAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8844,8848|false|false|false|C0199451|Continuous Positive Airway Pressure|CPAP
Event|Event|Hospital Course|8858,8862|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|8858,8862|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8858,8862|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8858,8862|false|false|false|C1553498|home health encounter|Home
Disorder|Disease or Syndrome|Hospital Course|8863,8867|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Meds
Event|Event|Hospital Course|8863,8867|false|false|false|||Meds
Finding|Intellectual Product|Hospital Course|8863,8867|false|false|false|C4284232|Medications|Meds
Drug|Organic Chemical|Hospital Course|8881,8891|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|8881,8891|false|false|false|C0028978|omeprazole|omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8897,8900|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8897,8900|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8897,8900|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8897,8900|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8897,8900|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|8905,8909|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Hospital Course|8905,8909|false|false|false|||GERD
Drug|Organic Chemical|Hospital Course|8922,8932|false|false|false|C0074393|sertraline|sertraline
Drug|Pharmacologic Substance|Hospital Course|8922,8932|false|false|false|C0074393|sertraline|sertraline
Event|Event|Hospital Course|8922,8932|false|false|false|||sertraline
Event|Event|Hospital Course|8939,8941|false|false|false|||PO
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8952,8962|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|8952,8962|false|false|false|||depression
Finding|Functional Concept|Hospital Course|8952,8962|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|8952,8962|false|false|false|C0460137;C1579931|Depression - motion|depression
Event|Event|Hospital Course|8965,8974|false|false|false|||Continued
Drug|Organic Chemical|Hospital Course|8975,8984|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8975,8984|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8992,8995|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8992,8995|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8992,8995|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|8992,8995|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8992,8995|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9003,9006|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|9003,9006|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|9003,9006|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|9003,9006|false|false|false|||NEB
Finding|Cell Function|Hospital Course|9003,9006|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9003,9006|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9014,9017|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|9018,9023|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|9018,9023|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|9018,9023|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|9018,9023|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|9025,9031|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|9025,9031|false|false|false|C0043144|Wheezing|wheeze
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9034,9038|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|Hospital Course|9034,9038|false|false|false|C0675390|ARID1A protein, human|Held
Event|Event|Hospital Course|9034,9038|false|false|false|||Held
Finding|Gene or Genome|Hospital Course|9034,9038|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|Hospital Course|9034,9038|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Drug|Organic Chemical|Hospital Course|9039,9045|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|9039,9045|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Event|Event|Hospital Course|9039,9045|false|false|false|||ProAir
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9048,9052|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|Hospital Course|9048,9052|false|false|false|C0675390|ARID1A protein, human|Held
Event|Event|Hospital Course|9048,9052|false|false|false|||Held
Finding|Gene or Genome|Hospital Course|9048,9052|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|Hospital Course|9048,9052|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Event|Event|Hospital Course|9053,9062|false|false|false|||trazadone
Drug|Hazardous or Poisonous Substance|Hospital Course|9077,9084|false|false|false|C0002772;C0242402|Analgesics, Opioid;Opioids|opioids
Drug|Organic Chemical|Hospital Course|9077,9084|false|false|false|C0002772;C0242402|Analgesics, Opioid;Opioids|opioids
Drug|Pharmacologic Substance|Hospital Course|9077,9084|false|false|false|C0002772;C0242402|Analgesics, Opioid;Opioids|opioids
Event|Event|Hospital Course|9077,9084|false|false|false|||opioids
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9087,9091|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|Hospital Course|9087,9091|false|false|false|C0675390|ARID1A protein, human|Held
Finding|Gene or Genome|Hospital Course|9087,9091|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|Hospital Course|9087,9091|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Drug|Organic Chemical|Hospital Course|9092,9102|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|9092,9102|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|9117,9120|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|9117,9120|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|9142,9152|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|9142,9152|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|Hospital Course|9142,9152|false|false|false|||gabapentin
Event|Event|Hospital Course|9158,9165|false|false|false|||helping
Event|Event|Hospital Course|9174,9180|false|false|false|||taking
Drug|Antibiotic|Hospital Course|9187,9199|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|Hospital Course|9187,9199|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|Hospital Course|9187,9199|false|false|false|||erythromycin
Event|Event|Hospital Course|9211,9217|false|false|false|||taking
Event|Event|Hospital Course|9219,9228|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|9219,9228|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Idea or Concept|Hospital Course|9232,9237|false|false|false|C0812371|Ortho-|Ortho
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9238,9243|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Hospital Course|9238,9243|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Hospital Course|9238,9243|false|false|false|C0150920|Spine Problem|spine
Event|Event|Hospital Course|9282,9289|false|false|false|||medical
Finding|Functional Concept|Hospital Course|9282,9289|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|9282,9289|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|9282,9289|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|9282,9289|false|false|false|C0199168|Medical service|medical
Event|Event|Hospital Course|9291,9298|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|9291,9298|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|9291,9298|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|9291,9298|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|Hospital Course|9299,9310|false|false|false|||significant
Finding|Idea or Concept|Hospital Course|9299,9310|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Hospital Course|9315,9318|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9315,9318|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Hospital Course|9315,9318|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|Hospital Course|9315,9318|false|false|false|||OSA
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9320,9328|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|Hospital Course|9320,9337|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Event|Event|Hospital Course|9329,9337|false|false|false|||aneurysm
Finding|Pathologic Function|Hospital Course|9329,9337|false|false|false|C0002940|Aneurysm|aneurysm
Disorder|Anatomical Abnormality|Hospital Course|9329,9355|false|false|false|C0162871|Aortic Aneurysm, Abdominal|aneurysm, abdominal aortic
Anatomy|Body Location or Region|Hospital Course|9339,9348|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9349,9355|false|false|false|C0003483|Aorta|aortic
Event|Event|Hospital Course|9357,9365|false|false|false|||aneurysm
Finding|Pathologic Function|Hospital Course|9357,9365|false|false|false|C0002940|Aneurysm|aneurysm
Disorder|Disease or Syndrome|Hospital Course|9367,9392|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid syndrome
Disorder|Disease or Syndrome|Hospital Course|9384,9392|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|9384,9392|false|false|false|||syndrome
Disorder|Disease or Syndrome|Hospital Course|9384,9394|false|false|false|C0796110|Pallister W syndrome|syndrome w
Disorder|Disease or Syndrome|Hospital Course|9405,9409|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|Hospital Course|9405,9409|false|false|false|||DVTs
Event|Event|Hospital Course|9419,9424|false|false|false|C0441471|Event|event
Finding|Gene or Genome|Hospital Course|9438,9443|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9444,9447|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|Hospital Course|9444,9447|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|Hospital Course|9444,9447|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9448,9459|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|9451,9459|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|9451,9459|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|9451,9459|false|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|9451,9459|false|false|false|||warfarin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9461,9466|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|Hospital Course|9461,9466|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Event|Event|Hospital Course|9461,9466|false|false|false|||BRCA1
Finding|Gene or Genome|Hospital Course|9461,9466|false|false|false|C0376571|BRCA1 gene|BRCA1
Disorder|Cell or Molecular Dysfunction|Hospital Course|9461,9475|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 mutation
Disorder|Cell or Molecular Dysfunction|Hospital Course|9467,9475|false|false|false|C1705285|Mutation Abnormality|mutation
Event|Event|Hospital Course|9467,9475|false|false|false|||mutation
Finding|Genetic Function|Hospital Course|9467,9475|false|false|false|C0026882|Mutation|mutation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9487,9493|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|9487,9493|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Hospital Course|9487,9493|false|false|false|||breast
Finding|Finding|Hospital Course|9487,9493|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9487,9493|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|Hospital Course|9487,9500|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|Hospital Course|9494,9500|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|9494,9500|false|false|false|||cancer
Event|Event|Hospital Course|9505,9515|false|false|false|||lumpectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9505,9515|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Event|Event|Hospital Course|9521,9529|false|false|false|||presents
Event|Event|Hospital Course|9545,9550|false|false|false|||month
Finding|Idea or Concept|Hospital Course|9545,9550|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|9545,9550|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Functional Concept|Hospital Course|9554,9559|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Sign or Symptom|Hospital Course|9554,9575|false|true|false|C2219286|right-sided low back pain|right lower back pain
Anatomy|Body Location or Region|Hospital Course|9560,9565|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|9560,9565|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|Hospital Course|9560,9570|false|false|false|C0230102;C2939142|Lower back (surface region);Lower back structure|lower back
Finding|Sign or Symptom|Hospital Course|9560,9575|false|true|false|C0024031|Low Back Pain|lower back pain
Finding|Sign or Symptom|Hospital Course|9566,9575|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Hospital Course|9571,9575|false|true|false|C2598155||pain
Event|Event|Hospital Course|9571,9575|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9571,9575|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9571,9575|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9581,9595|false|false|false|C0278147|Radicular pain|radicular pain
Attribute|Clinical Attribute|Hospital Course|9591,9595|false|false|false|C2598155||pain
Event|Event|Hospital Course|9591,9595|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9591,9595|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9591,9595|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|9606,9611|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9606,9615|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Finding|Sign or Symptom|Hospital Course|9606,9620|false|true|false|C5848135|Pain in right leg|right leg pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9612,9615|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|9612,9620|false|false|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Hospital Course|9616,9620|false|false|false|C2598155||pain
Event|Event|Hospital Course|9616,9620|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9616,9620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9616,9620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9621,9626|false|false|false|||found
Finding|Idea or Concept|Hospital Course|9635,9646|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9647,9651|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|Hospital Course|9647,9651|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|Hospital Course|9647,9651|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|Hospital Course|9647,9651|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|Hospital Course|9647,9651|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Disorder|Disease or Syndrome|Hospital Course|9647,9663|false|false|false|C0021818|Intervertebral Disk Displacement|disc herniations
Disorder|Anatomical Abnormality|Hospital Course|9652,9663|false|false|false|C0019270|Hernia|herniations
Event|Event|Hospital Course|9652,9663|false|false|false|||herniations
Event|Event|Hospital Course|9707,9717|false|false|false|||discectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9707,9717|false|false|false|C0206078|Diskectomy|discectomy
Event|Event|Hospital Course|9741,9747|false|false|false|||fusion
Finding|Functional Concept|Hospital Course|9741,9747|false|false|false|C0332466|Fused structure|fusion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9741,9747|false|false|false|C1293131|Fusion procedure|fusion
Event|Event|Hospital Course|9752,9760|false|false|false|||durotomy
Finding|Gene or Genome|Hospital Course|9777,9781|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|Post
Finding|Body Substance|Hospital Course|9794,9801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9794,9801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9794,9801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9806,9814|false|false|false|||admitted
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9826,9831|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|Spine
Anatomy|Cell Component|Hospital Course|9826,9831|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|Spine
Finding|Finding|Hospital Course|9826,9831|false|false|false|C0150920|Spine Problem|Spine
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9826,9839|false|false|false|C0920347;C2608059|Operation on spinal cord (procedure);Procedure on spinal cord (procedure)|Spine Surgery
Finding|Finding|Hospital Course|9832,9839|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Hospital Course|9832,9839|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Hospital Course|9832,9839|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9832,9839|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Occupational Activity|Hospital Course|9840,9847|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|9840,9847|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|9853,9858|false|false|false|||taken
Finding|Finding|Hospital Course|9866,9875|false|false|false|C4738506|Operating|Operating
Finding|Idea or Concept|Hospital Course|9889,9894|false|false|false|C1552828|Table Frame - above|above
Attribute|Clinical Attribute|Hospital Course|9895,9904|false|false|false|C0945766||procedure
Event|Event|Hospital Course|9895,9904|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|9895,9904|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|9895,9904|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9895,9904|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Hospital Course|9919,9927|false|false|false|||dictated
Attribute|Clinical Attribute|Hospital Course|9928,9942|false|false|false|C0551628||operative note
Event|Event|Hospital Course|9938,9942|false|false|false|||note
Event|Event|Hospital Course|9955,9962|false|false|false|||details
Event|Event|Hospital Course|9967,9974|false|false|false|||surgery
Finding|Finding|Hospital Course|9967,9974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|9967,9974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|9967,9974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9967,9974|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Hospital Course|9988,10000|false|false|false|||complication
Finding|Idea or Concept|Hospital Course|9988,10000|false|false|false|C0009566;C2362589|Complication;Complication (attribute)|complication
Finding|Pathologic Function|Hospital Course|9988,10000|false|false|false|C0009566;C2362589|Complication;Complication (attribute)|complication
Finding|Body Substance|Hospital Course|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10009,10016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|10021,10032|false|false|false|||transferred
Event|Event|Hospital Course|10040,10044|false|false|false|||PACU
Finding|Intellectual Product|Hospital Course|10051,10057|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|10058,10067|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|10058,10067|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|10058,10067|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|10058,10067|false|false|false|C1705253|Logical Condition|condition
Disorder|Disease or Syndrome|Hospital Course|10070,10087|false|false|false|C0589110|Postoperative deep vein thrombosis|Postoperative DVT
Anatomy|Body Location or Region|Hospital Course|10084,10087|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|10084,10087|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|10084,10087|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|10084,10087|false|false|false|||DVT
Finding|Gene or Genome|Hospital Course|10097,10101|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Event|Event|Hospital Course|10121,10125|false|false|false|||back
Drug|Organic Chemical|Hospital Course|10129,10136|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|10129,10136|false|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|10137,10143|false|false|false|||bridge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10137,10143|false|false|false|C0399080|Fixation of dental bridge|bridge
Drug|Organic Chemical|Hospital Course|10147,10155|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|10147,10155|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Hospital Course|10147,10155|false|false|false|||coumadin
Event|Activity|Hospital Course|10165,10173|false|false|false|C0441655|Activities|Activity
Event|Event|Hospital Course|10165,10173|false|false|false|||Activity
Finding|Daily or Recreational Activity|Hospital Course|10165,10173|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Hospital Course|10165,10173|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Hospital Course|10174,10182|false|false|false|||remained
Event|Event|Hospital Course|10188,10195|false|false|false|||bedrest
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10188,10195|false|false|false|C0004910|Bed rest|bedrest
Disorder|Injury or Poisoning|Hospital Course|10200,10210|false|false|false|C1504340|Dural tear|dural tear
Disorder|Injury or Poisoning|Hospital Course|10206,10210|false|false|false|C0043246;C3203359|Laceration;Rupture|tear
Finding|Body Substance|Hospital Course|10206,10210|false|false|false|C0039409|Tears (substance)|tear
Event|Event|Hospital Course|10211,10222|false|false|false|||precautions
Finding|Conceptual Entity|Hospital Course|10211,10222|false|false|false|C1882442|Precaution|precautions
Event|Event|Hospital Course|10231,10236|false|false|false|||hours
Event|Activity|Hospital Course|10240,10248|false|false|false|C0441655|Activities|Activity
Event|Event|Hospital Course|10240,10248|false|false|false|||Activity
Finding|Daily or Recreational Activity|Hospital Course|10240,10248|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Hospital Course|10240,10248|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Hospital Course|10253,10261|false|false|false|||advanced
Finding|Functional Concept|Hospital Course|10278,10289|false|false|false|C1522726|Intravenous Route of Administration|Intravenous
Drug|Antibiotic|Hospital Course|10290,10301|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|10290,10301|false|false|false|||antibiotics
Event|Event|Hospital Course|10308,10317|false|false|false|||continued
Event|Event|Hospital Course|10339,10347|false|false|false|||standard
Finding|Idea or Concept|Hospital Course|10339,10347|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Finding|Intellectual Product|Hospital Course|10339,10347|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Procedure|Laboratory Procedure|Hospital Course|10339,10347|false|false|false|C3873211|Standard base excess calculation technique|standard
Event|Event|Hospital Course|10348,10356|false|false|false|||protocol
Finding|Finding|Hospital Course|10348,10356|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|Hospital Course|10348,10356|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Idea or Concept|Hospital Course|10359,10366|false|false|false|C1555582|Initial (abbreviation)|Initial
Finding|Sign or Symptom|Hospital Course|10367,10378|false|false|false|C0030201|Pain, Postoperative|postop pain
Attribute|Clinical Attribute|Hospital Course|10374,10378|false|false|false|C2598155||pain
Event|Event|Hospital Course|10374,10378|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10374,10378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10374,10378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|10383,10393|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|10399,10403|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|10399,10403|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|10399,10403|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|10399,10403|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|Hospital Course|10411,10415|false|false|false|C2598155||pain
Event|Event|Hospital Course|10411,10415|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10411,10415|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10411,10415|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|10417,10427|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|10417,10427|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|10417,10427|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Food|Hospital Course|10428,10432|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Event|Event|Hospital Course|10428,10432|false|false|false|||Diet
Finding|Functional Concept|Hospital Course|10428,10432|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|Hospital Course|10428,10432|false|false|false|C0012159|Diet therapy|Diet
Event|Event|Hospital Course|10437,10445|false|false|false|||advanced
Event|Event|Hospital Course|10449,10458|false|false|false|||tolerated
Event|Event|Hospital Course|10469,10476|false|false|false|||removed
Finding|Finding|Hospital Course|10488,10496|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Hospital Course|10488,10496|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Hospital Course|10488,10496|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Hospital Course|10488,10504|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10488,10504|false|false|false|C0949766|Physical therapy|Physical therapy
Event|Event|Hospital Course|10497,10504|false|false|false|||therapy
Finding|Finding|Hospital Course|10497,10504|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|10497,10504|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10497,10504|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Functional Concept|Hospital Course|10509,10521|false|false|false|C0521127|Occupational|Occupational
Finding|Intellectual Product|Hospital Course|10509,10529|false|false|false|C1547993|Diagnostic Service Section ID - Occupational Therapy|Occupational therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10509,10529|false|false|false|C1318464|Occupational therapy (procedure)|Occupational therapy
Event|Event|Hospital Course|10522,10529|false|false|false|||therapy
Finding|Finding|Hospital Course|10522,10529|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|10522,10529|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10522,10529|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Hospital Course|10535,10544|false|false|false|||consulted
Event|Event|Hospital Course|10550,10562|false|false|false|||mobilization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10550,10562|false|false|false|C0185112;C2080791|Mobilization (procedure);physical therapy mobilization (treatment)|mobilization
Event|Event|Hospital Course|10563,10566|false|false|false|||OOB
Event|Event|Hospital Course|10570,10578|false|false|false|||ambulate
Finding|Finding|Hospital Course|10570,10578|false|false|false|C4036205|Ambulate|ambulate
Disorder|Disease or Syndrome|Hospital Course|10583,10586|false|false|false|C5443983|VISCERAL LEIOMYOPATHY, AFRICAN DEGENERATIVE|ADL
Event|Event|Hospital Course|10583,10586|false|false|false|||ADL
Finding|Daily or Recreational Activity|Hospital Course|10583,10586|false|false|false|C0001288;C1420005;C5960776|Activity of daily living (function);SGCA gene;SGCA wt Allele|ADL
Finding|Gene or Genome|Hospital Course|10583,10586|false|false|false|C0001288;C1420005;C5960776|Activity of daily living (function);SGCA gene;SGCA wt Allele|ADL
Finding|Gene or Genome|Hospital Course|10591,10595|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|Post
Event|Event|Hospital Course|10599,10605|false|false|false|||course
Event|Event|Hospital Course|10610,10617|false|false|false|||notable
Finding|Intellectual Product|Hospital Course|10622,10627|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Hospital Course|10622,10638|false|false|false|C0333276|Acute hemorrhage|acute blood loss
Disorder|Disease or Syndrome|Hospital Course|10622,10645|false|false|false|C0154286;C0154298|Acute posthaemorrhagic anaemia;Iron deficiency anemia secondary to chronic blood loss|acute blood loss anemia
Disorder|Disease or Syndrome|Hospital Course|10628,10633|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|10628,10633|false|false|false|||blood
Finding|Body Substance|Hospital Course|10628,10633|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|10628,10638|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|Hospital Course|10628,10638|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Disorder|Disease or Syndrome|Hospital Course|10628,10645|false|false|false|C0154286;C0154298;C0948824|Acute posthaemorrhagic anaemia;Anemia due to blood loss;Iron deficiency anemia secondary to chronic blood loss|blood loss anemia
Finding|Finding|Hospital Course|10634,10638|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Hospital Course|10639,10645|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|10639,10645|false|false|false|||anemia
Event|Event|Hospital Course|10648,10660|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|10648,10660|false|false|false|C0009806|Constipation|constipation
Attribute|Clinical Attribute|Hospital Course|10662,10666|false|false|false|C2598155||pain
Event|Event|Hospital Course|10662,10666|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10662,10666|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10662,10666|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|10671,10682|false|false|false|||hypokalemia
Finding|Finding|Hospital Course|10671,10682|false|false|false|C0020621|Hypokalemia|hypokalemia
Finding|Intellectual Product|Hospital Course|10684,10689|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Pathologic Function|Hospital Course|10684,10700|false|false|false|C0333276|Acute hemorrhage|Acute blood loss
Disorder|Disease or Syndrome|Hospital Course|10684,10707|false|false|false|C0154286;C0154298|Acute posthaemorrhagic anaemia;Iron deficiency anemia secondary to chronic blood loss|Acute blood loss anemia
Disorder|Disease or Syndrome|Hospital Course|10690,10695|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|10690,10695|false|false|false|||blood
Finding|Body Substance|Hospital Course|10690,10695|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|10690,10700|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|Hospital Course|10690,10700|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Disorder|Disease or Syndrome|Hospital Course|10690,10707|false|false|false|C0154286;C0154298;C0948824|Acute posthaemorrhagic anaemia;Anemia due to blood loss;Iron deficiency anemia secondary to chronic blood loss|blood loss anemia
Finding|Finding|Hospital Course|10696,10700|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Hospital Course|10701,10707|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|10701,10707|false|false|false|||anemia
Event|Event|Hospital Course|10712,10718|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|10712,10718|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|10731,10738|false|false|false|||require
Event|Event|Hospital Course|10739,10751|false|false|false|||intervention
Procedure|Health Care Activity|Hospital Course|10739,10751|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10739,10751|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Event|Event|Hospital Course|10761,10768|false|false|false|||treated
Event|Event|Hospital Course|10775,10784|false|false|false|||Immediate
Finding|Idea or Concept|Hospital Course|10775,10784|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|10775,10784|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|10775,10792|false|false|false|C1708470|Immediate Release Dosage Form|Immediate release
Event|Event|Hospital Course|10785,10792|false|false|false|||release
Finding|Functional Concept|Hospital Course|10785,10792|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|10785,10792|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10785,10792|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Drug|Organic Chemical|Hospital Course|10793,10801|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Hospital Course|10793,10801|false|false|false|C0026549|morphine|morphine
Event|Event|Hospital Course|10793,10801|false|false|false|||morphine
Drug|Organic Chemical|Hospital Course|10803,10809|false|false|false|C0699187|Valium|Valium
Drug|Pharmacologic Substance|Hospital Course|10803,10809|false|false|false|C0699187|Valium|Valium
Event|Event|Hospital Course|10803,10809|false|false|false|||Valium
Drug|Organic Chemical|Hospital Course|10814,10821|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Hospital Course|10814,10821|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Hospital Course|10814,10821|false|false|false|||Tylenol
Attribute|Clinical Attribute|Hospital Course|10826,10830|false|false|false|C2598155||pain
Event|Event|Hospital Course|10826,10830|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10826,10830|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10826,10830|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|10826,10838|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10826,10838|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Hospital Course|10831,10838|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|10831,10838|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|10831,10838|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|10831,10838|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|10831,10838|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|10831,10838|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|10831,10838|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Space or Junction|Hospital Course|10841,10845|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|10841,10845|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|10841,10845|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|10841,10845|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Clinical Drug|Hospital Course|10841,10855|false|false|false|C0357141||Oral Potassium
Drug|Biologically Active Substance|Hospital Course|10846,10855|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|10846,10855|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|10846,10855|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|10846,10855|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|10846,10855|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|10846,10855|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|10846,10855|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|10846,10855|false|false|false|C0202194|Potassium measurement|Potassium
Event|Event|Hospital Course|10860,10865|false|false|false|||given
Event|Event|Hospital Course|10870,10881|false|false|false|||hypokalemia
Finding|Finding|Hospital Course|10870,10881|false|false|false|C0020621|Hypokalemia|hypokalemia
Event|Event|Hospital Course|10909,10913|false|false|false|||labs
Lab|Laboratory or Test Result|Hospital Course|10909,10913|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Hospital Course|10928,10934|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|10928,10934|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Idea or Concept|Hospital Course|10938,10946|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|Hospital Course|10938,10953|false|false|false|C0488549||Hospital course
Finding|Finding|Hospital Course|10938,10953|false|false|false|C0489547|Hospital course|Hospital course
Event|Event|Hospital Course|10947,10953|false|false|false|||course
Event|Event|Hospital Course|10968,10980|false|false|false|||unremarkable
Finding|Idea or Concept|Hospital Course|10988,10991|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10988,10991|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|10996,11005|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10996,11005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10996,11005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10996,11005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10996,11005|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|11010,11017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11010,11017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11010,11017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|11022,11030|false|false|false|||afebrile
Finding|Finding|Hospital Course|11022,11030|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|11036,11042|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|11036,11042|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|Hospital Course|11043,11048|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|11043,11054|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|11043,11054|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|11049,11054|false|false|false|||signs
Finding|Finding|Hospital Course|11049,11054|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|11049,11054|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|11057,11068|false|false|false|||comfortable
Finding|Finding|Hospital Course|11057,11068|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Space or Junction|Hospital Course|11072,11076|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|11072,11076|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|11072,11076|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|11072,11076|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|11072,11081|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|11077,11081|false|false|false|C2598155||pain
Event|Event|Hospital Course|11077,11081|false|false|false|||pain
Finding|Functional Concept|Hospital Course|11077,11081|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11077,11081|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|11077,11089|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11077,11089|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Hospital Course|11082,11089|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|11082,11089|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|11082,11089|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|11082,11089|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|11082,11089|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|11082,11089|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|11082,11089|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Hospital Course|11094,11104|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|11107,11119|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|11115,11119|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|11115,11119|false|false|false|||diet
Finding|Functional Concept|Hospital Course|11115,11119|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|11115,11119|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|Hospital Course|11124,11135|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11124,11135|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11124,11135|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11124,11135|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|11124,11148|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|11139,11148|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|11139,11148|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|11167,11177|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11167,11177|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|11167,11182|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|11178,11182|false|false|false|||list
Finding|Intellectual Product|Hospital Course|11178,11182|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|11186,11194|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|11199,11207|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|11199,11207|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|11199,11207|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|11199,11207|false|false|false|||complete
Finding|Functional Concept|Hospital Course|11199,11207|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11199,11207|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|11212,11225|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|11212,11225|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|11212,11225|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|11212,11225|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|11241,11244|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|11245,11249|false|false|false|C2598155||Pain
Event|Event|Hospital Course|11245,11249|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|11245,11249|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|11245,11249|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|11252,11256|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|11257,11262|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|11257,11262|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|11267,11276|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|11267,11276|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11284,11287|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|11284,11287|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|11284,11287|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|11284,11287|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|11284,11287|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11295,11298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|11295,11298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|11295,11298|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|11295,11298|false|false|false|||NEB
Finding|Cell Function|Hospital Course|11295,11298|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|11295,11298|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|11306,11309|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|11310,11315|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|11310,11315|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|11310,11315|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|11310,11315|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|11317,11323|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|11317,11323|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|11328,11340|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11328,11340|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|11350,11353|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|11358,11366|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|11358,11366|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|11358,11366|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|11358,11373|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|11358,11373|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|11367,11373|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|11367,11373|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|11367,11373|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|11367,11373|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|11367,11373|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|11367,11373|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11384,11387|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11384,11387|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11384,11387|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11384,11387|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11384,11387|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11392,11402|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|11392,11402|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11412,11415|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11412,11415|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11412,11415|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11412,11415|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11412,11415|false|false|false|C1332410|BID gene|BID
Drug|Biomedical or Dental Material|Hospital Course|11420,11432|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|11420,11432|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|11420,11432|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|11420,11439|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|11420,11439|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|11433,11439|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|11433,11439|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|11433,11439|false|false|false|||Glycol
Finding|Gene or Genome|Hospital Course|11454,11457|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|11458,11470|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|11458,11470|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|11480,11484|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|11480,11484|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|11480,11484|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|Hospital Course|11480,11484|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|11489,11494|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|11489,11494|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|11512,11522|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|11512,11522|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|11543,11552|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|Hospital Course|11543,11552|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|Hospital Course|11566,11569|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|11570,11575|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|11570,11575|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|11570,11575|false|false|false|||sleep
Finding|Organism Function|Hospital Course|11570,11575|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|11581,11588|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|11581,11588|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|11581,11588|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|11581,11590|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|11581,11590|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|11581,11590|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|11581,11590|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|11581,11590|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|11595,11599|false|false|false|||UNIT
Drug|Hazardous or Poisonous Substance|Hospital Course|11614,11622|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|11614,11622|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|11614,11622|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|11636,11640|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Organic Chemical|Hospital Course|11652,11661|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|11652,11661|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|Hospital Course|11652,11661|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|Hospital Course|11665,11670|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|11665,11670|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11673,11677|false|false|false|C4308013|PTCH1 protein, human|PTCH
Event|Event|Hospital Course|11673,11677|false|false|false|||PTCH
Finding|Gene or Genome|Hospital Course|11673,11677|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|Hospital Course|11673,11677|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Event|Event|Hospital Course|11681,11684|false|false|false|||QAM
Finding|Functional Concept|Hospital Course|11685,11690|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|11685,11694|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11691,11694|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11691,11694|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|11691,11694|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|11691,11694|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|Hospital Course|11691,11694|false|false|false|||hip
Finding|Gene or Genome|Hospital Course|11691,11694|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11691,11694|false|false|false|C1292890|Procedure on hip|hip
Drug|Organic Chemical|Hospital Course|11700,11710|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|11700,11710|false|false|false|C0016860|furosemide|Furosemide
Finding|Gene or Genome|Hospital Course|11726,11729|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11730,11733|false|false|false|C0023216;C1140621|Leg;Lower Extremity|Leg
Finding|Pathologic Function|Hospital Course|11730,11742|false|false|false|C0581394|Swelling of lower limb|Leg swelling
Event|Event|Hospital Course|11734,11742|false|false|false|||swelling
Finding|Finding|Hospital Course|11734,11742|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|11734,11742|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Hospital Course|11748,11754|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|11748,11754|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|11748,11758|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|11748,11758|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|11755,11758|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|11755,11758|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|11755,11758|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Organic Chemical|Hospital Course|11760,11769|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|11760,11769|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|11760,11777|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|11760,11777|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|11770,11777|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|11770,11777|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|11770,11777|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|11770,11777|false|false|false|||sulfate
Event|Event|Hospital Course|11796,11806|false|false|false|||inhalation
Finding|Functional Concept|Hospital Course|11796,11806|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|11796,11806|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|Hospital Course|11812,11815|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Hazardous or Poisonous Substance|Hospital Course|11821,11829|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|11821,11829|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|11821,11829|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|11841,11845|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Organic Chemical|Hospital Course|11857,11867|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|11857,11867|false|false|false|C0060926|gabapentin|Gabapentin
Event|Event|Hospital Course|11878,11881|false|false|false|||TID
Drug|Organic Chemical|Hospital Course|11887,11895|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|Hospital Course|11887,11895|false|false|false|C0040610|tramadol|TraMADol
Event|Event|Hospital Course|11887,11895|false|false|false|||TraMADol
Procedure|Laboratory Procedure|Hospital Course|11887,11895|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|Hospital Course|11909,11912|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|11913,11917|false|false|false|C2598155||Pain
Event|Event|Hospital Course|11913,11917|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|11913,11917|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|11913,11917|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|11920,11928|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|11920,11928|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|11933,11942|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11933,11942|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11933,11942|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11933,11942|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11933,11942|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11933,11954|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|11943,11954|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11943,11954|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11943,11954|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11943,11954|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|11960,11968|false|false|false|C0012010|diazepam|Diazepam
Drug|Pharmacologic Substance|Hospital Course|11960,11968|false|false|false|C0012010|diazepam|Diazepam
Finding|Gene or Genome|Hospital Course|11981,11984|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|11985,11989|false|false|false|C2598155||pain
Event|Event|Hospital Course|11985,11989|false|false|false|||pain
Finding|Functional Concept|Hospital Course|11985,11989|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11985,11989|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|Hospital Course|11990,11995|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|Hospital Course|11990,11995|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Event|Event|Hospital Course|12001,12006|false|false|false|||cause
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12007,12017|false|true|false|C2830004|Somnolence|drowsiness
Event|Event|Hospital Course|12007,12017|false|false|false|||drowsiness
Finding|Finding|Hospital Course|12007,12017|false|true|false|C0013144|Drowsiness|drowsiness
Event|Event|Hospital Course|12019,12021|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|12023,12031|false|false|false|C0012010|diazepam|diazepam
Drug|Pharmacologic Substance|Hospital Course|12023,12031|false|false|false|C0012010|diazepam|diazepam
Event|Event|Hospital Course|12023,12031|false|false|false|||diazepam
Drug|Biomedical or Dental Material|Hospital Course|12039,12045|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|12039,12045|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|12046,12054|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12049,12054|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12049,12054|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|12077,12081|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|12077,12081|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|12088,12094|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12095,12102|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12095,12102|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12111,12121|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|12111,12121|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|12111,12121|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|12111,12128|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|12111,12128|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|12122,12128|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12122,12128|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12122,12128|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12122,12128|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12122,12128|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12122,12128|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Disease or Syndrome|Hospital Course|12144,12169|false|false|false|C0085278|Antiphospholipid Syndrome|Antiphospholipid Syndrome
Disorder|Disease or Syndrome|Hospital Course|12161,12169|false|false|false|C0039082|Syndrome|Syndrome
Event|Event|Hospital Course|12161,12169|false|false|false|||Syndrome
Event|Event|Hospital Course|12171,12180|false|false|false|||Treatment
Finding|Conceptual Entity|Hospital Course|12171,12180|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Finding|Functional Concept|Hospital Course|12171,12180|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Procedure|Health Care Activity|Hospital Course|12171,12180|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12171,12180|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12181,12187|false|false|false|C0399080|Fixation of dental bridge|Bridge
Drug|Organic Chemical|Hospital Course|12201,12209|false|false|false|C0026549|morphine|Morphine
Drug|Pharmacologic Substance|Hospital Course|12201,12209|false|false|false|C0026549|morphine|Morphine
Event|Event|Hospital Course|12201,12209|false|false|false|||Morphine
Drug|Organic Chemical|Hospital Course|12201,12217|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Pharmacologic Substance|Hospital Course|12201,12217|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Finding|Gene or Genome|Hospital Course|12235,12238|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12239,12243|false|false|false|C2598155||Pain
Event|Event|Hospital Course|12239,12243|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|12239,12243|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|12239,12243|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|12246,12252|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Hospital Course|12246,12252|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Event|Event|Hospital Course|12268,12275|false|false|false|||operate
Disorder|Injury or Poisoning|Hospital Course|12282,12291|false|false|false|C0337246|Contact with machinery|machinery
Event|Event|Hospital Course|12282,12291|false|false|false|||machinery
Event|Event|Hospital Course|12293,12298|false|false|false|||drink
Drug|Organic Chemical|Hospital Course|12299,12306|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|12299,12306|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Hospital Course|12299,12306|false|false|false|||alcohol
Finding|Intellectual Product|Hospital Course|12299,12306|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|Hospital Course|12310,12315|false|false|false|||drive
Finding|Mental Process|Hospital Course|12310,12315|false|false|false|C0013126|Intrinsic drive|drive
Event|Event|Hospital Course|12317,12319|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|12321,12329|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Hospital Course|12321,12329|false|false|false|C0026549|morphine|morphine
Event|Event|Hospital Course|12321,12329|false|false|false|||morphine
Drug|Biomedical or Dental Material|Hospital Course|12338,12344|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|12348,12356|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12351,12356|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12351,12356|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|12377,12381|false|false|false|||Disp
Drug|Biomedical or Dental Material|Hospital Course|12388,12394|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12395,12402|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12395,12402|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12411,12421|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|12411,12421|false|false|false|C0016860|furosemide|Furosemide
Finding|Gene or Genome|Hospital Course|12437,12440|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12441,12444|false|false|false|C0023216;C1140621|Leg;Lower Extremity|Leg
Finding|Pathologic Function|Hospital Course|12441,12453|false|false|false|C0581394|Swelling of lower limb|Leg swelling
Event|Event|Hospital Course|12445,12453|false|false|false|||swelling
Finding|Finding|Hospital Course|12445,12453|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|12445,12453|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Hospital Course|12460,12473|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|12460,12473|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|12460,12473|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|12460,12473|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|12489,12492|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12493,12497|false|false|false|C2598155||Pain
Event|Event|Hospital Course|12493,12497|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|12493,12497|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|12493,12497|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|12500,12504|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|12505,12510|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|12505,12510|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|12517,12526|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|12517,12526|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12534,12537|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|12534,12537|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|12534,12537|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|12534,12537|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|12534,12537|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12545,12548|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|12545,12548|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|12545,12548|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|12545,12548|false|false|false|||NEB
Finding|Cell Function|Hospital Course|12545,12548|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|12545,12548|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|12556,12559|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|12560,12565|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|12560,12565|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|12560,12565|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|12560,12565|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|12567,12573|false|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|12567,12573|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|12580,12592|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12580,12592|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|12602,12605|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|12612,12620|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|12612,12620|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|12612,12620|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|12612,12627|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|12612,12627|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|12621,12627|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12621,12627|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12621,12627|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12621,12627|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12621,12627|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12621,12627|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12638,12641|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12638,12641|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12638,12641|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12638,12641|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12638,12641|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12648,12657|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|12648,12657|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|Hospital Course|12648,12657|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|Hospital Course|12661,12666|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|12661,12666|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12669,12673|false|false|false|C4308013|PTCH1 protein, human|PTCH
Event|Event|Hospital Course|12669,12673|false|false|false|||PTCH
Finding|Gene or Genome|Hospital Course|12669,12673|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|Hospital Course|12669,12673|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Event|Event|Hospital Course|12677,12680|false|false|false|||QAM
Finding|Functional Concept|Hospital Course|12681,12686|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|12681,12690|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12687,12690|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12687,12690|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|12687,12690|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|12687,12690|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|Hospital Course|12687,12690|false|false|false|||hip
Finding|Gene or Genome|Hospital Course|12687,12690|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12687,12690|false|false|false|C1292890|Procedure on hip|hip
Drug|Organic Chemical|Hospital Course|12698,12708|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|12698,12708|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12718,12721|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12718,12721|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12718,12721|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12718,12721|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12718,12721|false|false|false|C1332410|BID gene|BID
Drug|Biomedical or Dental Material|Hospital Course|12729,12741|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|12729,12741|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|12729,12741|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|12729,12748|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|12729,12748|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|12742,12748|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|12742,12748|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|12742,12748|false|false|false|||Glycol
Finding|Gene or Genome|Hospital Course|12763,12766|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|12767,12779|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|12767,12779|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|12789,12793|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|12789,12793|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|12789,12793|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|Hospital Course|12789,12793|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|12801,12807|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|12801,12807|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|12801,12811|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|12801,12811|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|12808,12811|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|12808,12811|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|12808,12811|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Organic Chemical|Hospital Course|12813,12822|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|12813,12822|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|12813,12830|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|12813,12830|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12823,12830|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|12823,12830|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|12823,12830|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|12823,12830|false|false|false|||sulfate
Event|Event|Hospital Course|12849,12859|false|false|false|||inhalation
Finding|Functional Concept|Hospital Course|12849,12859|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|12849,12859|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|Hospital Course|12865,12868|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|12876,12881|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|12876,12881|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|12902,12912|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|12902,12912|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|12936,12945|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|Hospital Course|12936,12945|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|Hospital Course|12959,12962|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|12963,12968|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|12963,12968|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|12963,12968|false|false|false|||sleep
Finding|Organism Function|Hospital Course|12963,12968|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|12976,12983|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12976,12983|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12976,12983|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12976,12985|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12976,12985|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12976,12985|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12976,12985|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12976,12985|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|12990,12994|false|false|false|||UNIT
Drug|Hazardous or Poisonous Substance|Hospital Course|13011,13019|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|13011,13019|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|13011,13019|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|13031,13035|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Hazardous or Poisonous Substance|Hospital Course|13049,13057|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|13049,13057|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|13049,13057|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|13071,13075|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Event|Event|Hospital Course|13087,13096|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13087,13096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13087,13096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13087,13096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13087,13096|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|13087,13108|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|13087,13108|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|13097,13108|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|13097,13108|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|13097,13108|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|13110,13118|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|13110,13118|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|13110,13123|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|13119,13123|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|13119,13123|false|false|false|||Care
Finding|Finding|Hospital Course|13119,13123|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|13119,13123|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|13126,13134|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|13126,13134|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|13142,13151|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13142,13151|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13142,13151|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13142,13151|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13142,13151|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13142,13161|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|13152,13161|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|13152,13161|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|13152,13161|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|13152,13161|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|13152,13161|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Location or Region|Hospital Course|13164,13170|false|false|false|C0024090|Lumbar Region|Lumbar
Disorder|Disease or Syndrome|Hospital Course|13164,13186|false|false|false|C0158288|Spinal stenosis of lumbar region|Lumbar spinal stenosis
Disorder|Acquired Abnormality|Hospital Course|13171,13186|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|spinal stenosis
Disorder|Anatomical Abnormality|Hospital Course|13171,13186|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|spinal stenosis
Event|Event|Hospital Course|13178,13186|false|false|false|||stenosis
Finding|Pathologic Function|Hospital Course|13178,13186|false|false|false|C1261287|Stenosis|stenosis
Disorder|Acquired Abnormality|Hospital Course|13189,13206|false|false|false|C0038016;C0038017;C2242765|Acquired spondylolisthesis;Congenital spondylolisthesis;Spondylolisthesis|Spondylolisthesis
Disorder|Congenital Abnormality|Hospital Course|13189,13206|false|false|false|C0038016;C0038017;C2242765|Acquired spondylolisthesis;Congenital spondylolisthesis;Spondylolisthesis|Spondylolisthesis
Disorder|Disease or Syndrome|Hospital Course|13189,13206|false|false|false|C0038016;C0038017;C2242765|Acquired spondylolisthesis;Congenital spondylolisthesis;Spondylolisthesis|Spondylolisthesis
Event|Event|Hospital Course|13189,13206|false|false|false|||Spondylolisthesis
Finding|Finding|Hospital Course|13189,13213|false|false|false|C5542839|Spondylolisthesis, L4-L5|Spondylolisthesis, L4-L5
Disorder|Disease or Syndrome|Hospital Course|13216,13219|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13216,13219|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|13216,13219|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|13216,13219|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|13216,13219|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|Hospital Course|13221,13233|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|13221,13233|false|false|false|C0009806|Constipation|Constipation
Disorder|Neoplastic Process|Hospital Course|13235,13244|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Hospital Course|13235,13244|false|false|false|||Secondary
Finding|Functional Concept|Hospital Course|13235,13244|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|Hospital Course|13245,13254|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|Hospital Course|13245,13254|false|false|false|C0011900|Diagnosis|Diagnoses
Event|Event|Hospital Course|13258,13265|false|false|false|||History
Finding|Conceptual Entity|Hospital Course|13258,13265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|13258,13265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|13258,13265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|13258,13268|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|13269,13272|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|13269,13272|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|13269,13272|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|13269,13272|false|false|false|||DVT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13278,13303|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Drug|Immunologic Factor|Hospital Course|13278,13303|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Finding|Finding|Hospital Course|13278,13303|false|false|false|C4019436|Antiphospholipid antibody positivity|Antiphospholipid antibody
Disorder|Disease or Syndrome|Hospital Course|13278,13312|false|false|false|C0085278|Antiphospholipid Syndrome|Antiphospholipid antibody syndrome
Anatomy|Cell Component|Hospital Course|13295,13303|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13295,13303|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Hospital Course|13295,13303|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Hospital Course|13295,13303|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Hospital Course|13295,13303|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Hospital Course|13304,13312|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|13304,13312|false|false|false|||syndrome
Disorder|Anatomical Abnormality|Hospital Course|13315,13318|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Hospital Course|13315,13318|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13315,13318|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Hospital Course|13315,13318|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Hospital Course|13315,13318|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Hospital Course|13315,13318|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|Hospital Course|13315,13318|false|false|false|||AAA
Finding|Gene or Genome|Hospital Course|13315,13318|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Disorder|Disease or Syndrome|Hospital Course|13321,13324|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13321,13324|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Hospital Course|13321,13324|false|false|false|C0764906|OSA protein, Drosophila|OSA
Event|Event|Hospital Course|13321,13324|false|false|false|||OSA
Event|Event|Hospital Course|13328,13332|false|false|false|||CPAP
Finding|Gene or Genome|Hospital Course|13328,13332|false|false|false|C1424863|CENPJ gene|CPAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13328,13332|false|false|false|C0199451|Continuous Positive Airway Pressure|CPAP
Finding|Mental Process|Discharge Condition|13358,13364|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13358,13371|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13358,13371|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13365,13371|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13365,13371|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13373,13378|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13373,13378|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13383,13391|false|false|false|||coherent
Finding|Finding|Discharge Condition|13383,13391|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13393,13398|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13393,13415|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13393,13415|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13402,13415|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13402,13415|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13402,13415|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13417,13422|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13417,13422|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13417,13422|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13417,13422|false|false|false|||Alert
Finding|Finding|Discharge Condition|13417,13422|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13417,13422|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13417,13422|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13427,13438|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13427,13438|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|13440,13448|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|13440,13448|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|13440,13448|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|13449,13455|false|false|false|C5889824||Status
Event|Event|Discharge Condition|13449,13455|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|13449,13455|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|13457,13467|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|13457,13467|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|13457,13467|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|13457,13467|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|13470,13478|false|false|false|||requires
Event|Event|Discharge Condition|13479,13489|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|13479,13489|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|13493,13496|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|13493,13496|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|13493,13496|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|13493,13496|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|13493,13496|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|13498,13504|false|false|false|||walker
Event|Event|Discharge Instructions|13552,13560|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|13552,13560|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|13552,13560|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|13564,13568|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|13564,13568|false|false|false|||care
Finding|Finding|Discharge Instructions|13564,13568|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13564,13568|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|13609,13613|false|false|false|||come
Finding|Idea or Concept|Discharge Instructions|13621,13629|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|13640,13644|false|false|false|||came
Finding|Idea or Concept|Discharge Instructions|13652,13660|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|13685,13694|false|false|false|||worsening
Finding|Idea or Concept|Discharge Instructions|13685,13694|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Finding|Sign or Symptom|Discharge Instructions|13696,13705|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Discharge Instructions|13701,13705|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|13701,13705|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|13701,13705|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13701,13705|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|13711,13715|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|13711,13715|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|13711,13715|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13711,13715|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|13716,13725|false|false|false|||radiating
Finding|Functional Concept|Discharge Instructions|13736,13741|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13736,13745|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13742,13745|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Attribute|Clinical Attribute|Discharge Instructions|13752,13756|false|true|false|C2598155||pain
Event|Event|Discharge Instructions|13752,13756|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|13752,13756|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13752,13756|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|13758,13765|false|false|false|||started
Finding|Idea or Concept|Discharge Instructions|13774,13779|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Discharge Instructions|13774,13779|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|Discharge Instructions|13780,13783|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Discharge Instructions|13806,13811|false|false|false|||worse
Finding|Finding|Discharge Instructions|13806,13811|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|13806,13811|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Event|Discharge Instructions|13813,13819|false|false|false|||making
Event|Event|Discharge Instructions|13824,13833|false|false|false|||difficult
Finding|Finding|Discharge Instructions|13824,13833|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|Discharge Instructions|13837,13841|false|false|false|||walk
Event|Event|Discharge Instructions|13856,13863|false|false|false|||burning
Finding|Sign or Symptom|Discharge Instructions|13856,13863|false|false|false|C0085624|Burning sensation|burning
Finding|Sign or Symptom|Discharge Instructions|13856,13868|false|false|false|C0234230|Pain, Burning|burning pain
Attribute|Clinical Attribute|Discharge Instructions|13864,13868|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|13864,13868|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|13864,13868|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13864,13868|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|13864,13883|false|false|false|C0013428|Dysuria|pain with urination
Event|Event|Discharge Instructions|13874,13883|false|false|false|||urination
Finding|Organism Function|Discharge Instructions|13874,13883|false|false|false|C0042034|Urination|urination
Event|Event|Discharge Instructions|13899,13906|false|false|false|||receive
Finding|Idea or Concept|Discharge Instructions|13914,13922|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|13939,13942|false|false|false|||MRI
Finding|Gene or Genome|Discharge Instructions|13939,13942|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Discharge Instructions|13939,13942|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Discharge Instructions|13939,13942|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Discharge Instructions|13948,13954|false|false|false|||showed
Finding|Idea or Concept|Discharge Instructions|13955,13966|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13967,13971|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|Discharge Instructions|13967,13971|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|Discharge Instructions|13967,13971|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|Discharge Instructions|13967,13971|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|Discharge Instructions|13967,13971|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Disorder|Disease or Syndrome|Discharge Instructions|13967,13982|false|false|false|C0021818|Intervertebral Disk Displacement|disc herniation
Disorder|Anatomical Abnormality|Discharge Instructions|13972,13982|false|false|false|C0019270|Hernia|herniation
Event|Event|Discharge Instructions|13972,13982|false|false|false|||herniation
Anatomy|Body Location or Region|Discharge Instructions|13992,13997|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Discharge Instructions|13992,13997|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|Discharge Instructions|13992,14002|false|false|false|C0230102;C2939142|Lower back (surface region);Lower back structure|lower back
Event|Event|Discharge Instructions|14018,14023|false|false|false|||cause
Finding|Conceptual Entity|Discharge Instructions|14018,14023|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Discharge Instructions|14018,14023|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Attribute|Clinical Attribute|Discharge Instructions|14032,14036|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|14032,14036|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|14032,14036|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14032,14036|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14042,14047|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Discharge Instructions|14042,14047|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Discharge Instructions|14042,14047|false|false|false|C0150920|Spine Problem|spine
Event|Event|Discharge Instructions|14048,14056|false|false|false|||surgeons
Event|Event|Discharge Instructions|14058,14062|false|false|false|||felt
Event|Event|Discharge Instructions|14078,14085|false|false|false|||benefit
Event|Event|Discharge Instructions|14091,14098|false|false|false|||surgery
Finding|Finding|Discharge Instructions|14091,14098|false|false|true|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|14091,14098|false|false|true|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|14091,14098|false|false|true|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14091,14098|false|false|true|C0543467|Operative Surgical Procedures|surgery
Attribute|Clinical Attribute|Discharge Instructions|14115,14119|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|14115,14119|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|14115,14119|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14115,14119|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|14125,14133|false|false|false|||constant
Finding|Intellectual Product|Discharge Instructions|14125,14133|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Event|Event|Discharge Instructions|14138,14147|false|false|false|||worsening
Finding|Idea or Concept|Discharge Instructions|14162,14167|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Discharge Instructions|14162,14167|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|Discharge Instructions|14172,14176|false|false|false|||gave
Attribute|Clinical Attribute|Discharge Instructions|14181,14185|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|14181,14185|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|14181,14185|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14181,14185|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|14187,14198|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|14187,14198|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|14187,14198|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|14187,14198|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|14203,14210|false|false|false|||stopped
Drug|Hazardous or Poisonous Substance|Discharge Instructions|14216,14224|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Discharge Instructions|14216,14224|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Discharge Instructions|14216,14224|false|false|false|C0043031|warfarin|warfarin
Event|Event|Discharge Instructions|14216,14224|false|false|false|||warfarin
Event|Event|Discharge Instructions|14238,14242|false|false|false|||safe
Finding|Intellectual Product|Discharge Instructions|14238,14242|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|Discharge Instructions|14260,14267|false|false|false|||surgery
Finding|Finding|Discharge Instructions|14260,14267|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|14260,14267|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|14260,14267|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14260,14267|false|false|false|C0543467|Operative Surgical Procedures|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14279,14299|false|false|false|C0022983;C0408670|Decompression of spinal cord;Laminectomy|spinal decompression
Event|Event|Discharge Instructions|14286,14299|false|false|false|||decompression
Finding|Functional Concept|Discharge Instructions|14286,14299|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|Discharge Instructions|14286,14299|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14286,14299|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Event|Event|Discharge Instructions|14317,14321|false|false|false|||gave
Drug|Antibiotic|Discharge Instructions|14326,14337|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|14326,14337|false|false|false|||antibiotics
Finding|Sign or Symptom|Discharge Instructions|14347,14354|false|false|false|C0085624|Burning sensation|burning
Finding|Sign or Symptom|Discharge Instructions|14347,14359|false|false|false|C0234230|Pain, Burning|burning pain
Attribute|Clinical Attribute|Discharge Instructions|14355,14359|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|14355,14359|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|14355,14359|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14355,14359|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14355,14374|false|false|false|C0013428|Dysuria|pain with urination
Event|Event|Discharge Instructions|14365,14374|false|false|false|||urination
Finding|Organism Function|Discharge Instructions|14365,14374|false|false|false|C0042034|Urination|urination
Event|Event|Discharge Instructions|14386,14393|false|false|false|||believe
Event|Event|Discharge Instructions|14398,14404|false|false|false|||caused
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14410,14417|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14410,14423|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|Discharge Instructions|14410,14423|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|Discharge Instructions|14410,14433|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14418,14423|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|Discharge Instructions|14424,14433|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|14424,14433|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|14424,14433|false|false|false|C3714514|Infection|infection
Finding|Intellectual Product|Discharge Instructions|14456,14460|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Discharge Instructions|14465,14470|false|false|false|||leave
Finding|Idea or Concept|Discharge Instructions|14475,14483|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|14488,14494|false|false|false|C0024090|Lumbar Region|Lumbar
Event|Event|Discharge Instructions|14495,14508|false|false|false|||Decompression
Finding|Functional Concept|Discharge Instructions|14495,14508|false|false|false|C1965697|Decompression - action (qualifier value)|Decompression
Phenomenon|Phenomenon or Process|Discharge Instructions|14495,14508|false|false|false|C0011117|external decompression|Decompression
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14495,14508|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|Decompression
Event|Event|Discharge Instructions|14514,14520|false|false|false|||Fusion
Finding|Functional Concept|Discharge Instructions|14514,14520|false|false|false|C0332466|Fused structure|Fusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14514,14520|false|false|false|C1293131|Fusion procedure|Fusion
Event|Event|Discharge Instructions|14532,14541|false|false|false|||undergone
Event|Activity|Discharge Instructions|14556,14565|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|14556,14565|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|14556,14565|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14556,14565|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Anatomy|Body Location or Region|Discharge Instructions|14567,14573|false|false|false|C0024090|Lumbar Region|Lumbar
Event|Event|Discharge Instructions|14574,14587|false|false|false|||Decompression
Finding|Functional Concept|Discharge Instructions|14574,14587|false|false|false|C1965697|Decompression - action (qualifier value)|Decompression
Phenomenon|Phenomenon or Process|Discharge Instructions|14574,14587|false|false|false|C0011117|external decompression|Decompression
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14574,14587|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|Decompression
Event|Event|Discharge Instructions|14594,14600|false|false|false|||Fusion
Finding|Functional Concept|Discharge Instructions|14594,14600|false|false|false|C0332466|Fused structure|Fusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14594,14600|false|false|false|C1293131|Fusion procedure|Fusion
Event|Activity|Discharge Instructions|14624,14633|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|14624,14633|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|14624,14633|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14624,14633|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Event|Activity|Discharge Instructions|14653,14661|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Instructions|14653,14661|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Instructions|14653,14661|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Discharge Instructions|14677,14681|false|false|false|||lift
Procedure|Laboratory Procedure|Discharge Instructions|14708,14711|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|14741,14752|false|false|false|||comfortable
Finding|Finding|Discharge Instructions|14741,14752|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|Discharge Instructions|14768,14771|false|false|false|||sit
Finding|Finding|Discharge Instructions|14768,14771|true|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Gene or Genome|Discharge Instructions|14768,14771|true|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Finding|Discharge Instructions|14775,14780|true|true|false|C0038137;C0596013|Does stand;standards characteristics|stand
Finding|Functional Concept|Discharge Instructions|14775,14780|true|true|false|C0038137;C0596013|Does stand;standards characteristics|stand
Event|Event|Discharge Instructions|14826,14833|false|false|false|||walking
Event|Event|Discharge Instructions|14860,14874|false|false|false|||Rehabilitation
Finding|Finding|Discharge Instructions|14860,14874|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Finding|Functional Concept|Discharge Instructions|14860,14874|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14860,14874|false|false|false|C0034991|Rehabilitation therapy|Rehabilitation
Event|Event|Discharge Instructions|14876,14884|false|false|false|||Physical
Finding|Finding|Discharge Instructions|14876,14884|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Discharge Instructions|14876,14884|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Discharge Instructions|14876,14884|false|false|false|C0031809|Physical Examination|Physical
Finding|Idea or Concept|Discharge Instructions|14898,14901|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|14898,14901|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|14922,14926|false|false|false|||walk
Finding|Daily or Recreational Activity|Discharge Instructions|14922,14926|false|false|false|C0080331|Walking (function)|walk
Finding|Idea or Concept|Discharge Instructions|14946,14950|false|false|false|C1552020|Role Class - part|part
Event|Activity|Discharge Instructions|14960,14968|false|false|false|C0237820||recovery
Event|Event|Discharge Instructions|14960,14968|false|false|false|||recovery
Finding|Organism Function|Discharge Instructions|14960,14968|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|Discharge Instructions|14977,14981|false|false|false|||walk
Finding|Finding|Discharge Instructions|14985,14989|false|false|false|C4281574|Much|much
Event|Event|Discharge Instructions|15001,15009|false|false|false|||tolerate
Event|Event|Discharge Instructions|15020,15024|false|false|false|||kind
Finding|Intellectual Product|Discharge Instructions|15020,15024|false|false|false|C1706124|Terminology Kind|kind
Event|Activity|Discharge Instructions|15029,15036|false|false|false|C0206244|Lifting|lifting
Drug|Food|Discharge Instructions|15056,15060|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Event|Event|Discharge Instructions|15056,15060|false|false|false|||Diet
Finding|Functional Concept|Discharge Instructions|15056,15060|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|Discharge Instructions|15056,15060|false|false|false|C0012159|Diet therapy|Diet
Finding|Gene or Genome|Discharge Instructions|15062,15065|false|false|false|C0013470;C1708811|Eating;MCL1 wt Allele|Eat
Finding|Organism Function|Discharge Instructions|15062,15065|false|false|false|C0013470;C1708811|Eating;MCL1 wt Allele|Eat
Finding|Finding|Discharge Instructions|15075,15087|false|false|false|C0452415|Diet, Healthy|healthy diet
Drug|Food|Discharge Instructions|15083,15087|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|15083,15087|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|15083,15087|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|15083,15087|false|false|false|C0012159|Diet therapy|diet
Event|Event|Discharge Instructions|15107,15119|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|15107,15119|false|false|false|C0009806|Constipation|constipation
Finding|Finding|Discharge Instructions|15120,15133|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|Discharge Instructions|15126,15133|false|false|false|||surgery
Finding|Finding|Discharge Instructions|15126,15133|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|15126,15133|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|15126,15133|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15126,15133|false|false|false|C0543467|Operative Surgical Procedures|surgery
Drug|Pharmacologic Substance|Discharge Instructions|15154,15164|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|15154,15164|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|15154,15164|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|15169,15173|false|false|false|||help
Event|Activity|Discharge Instructions|15184,15189|false|false|false|C5966184|Issue (action)|issue
Event|Event|Discharge Instructions|15184,15189|false|false|false|||issue
Finding|Finding|Discharge Instructions|15184,15189|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|Discharge Instructions|15184,15189|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|Discharge Instructions|15209,15214|false|false|false|||Brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15209,15214|false|false|false|C1828220|Application of brace (procedure)|Brace
Event|Event|Discharge Instructions|15241,15246|false|false|false|||brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15241,15246|false|false|false|C1828220|Application of brace (procedure)|brace
Event|Event|Discharge Instructions|15273,15278|false|false|false|||brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15273,15278|false|false|false|C1828220|Application of brace (procedure)|brace
Event|Event|Discharge Instructions|15284,15289|false|false|false|||brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15284,15289|false|false|false|C1828220|Application of brace (procedure)|brace
Event|Event|Discharge Instructions|15299,15303|false|false|false|||worn
Event|Event|Discharge Instructions|15318,15325|false|false|false|||walking
Finding|Daily or Recreational Activity|Discharge Instructions|15318,15325|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|Discharge Instructions|15318,15325|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|Discharge Instructions|15318,15325|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Event|Discharge Instructions|15334,15338|false|false|false|||take
Event|Event|Discharge Instructions|15351,15358|false|false|false|||sitting
Event|Event|Discharge Instructions|15380,15385|false|false|false|||lying
Disorder|Disease or Syndrome|Discharge Instructions|15389,15392|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|Discharge Instructions|15389,15392|false|false|false|||bed
Finding|Intellectual Product|Discharge Instructions|15389,15392|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Injury or Poisoning|Discharge Instructions|15412,15417|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|Discharge Instructions|15412,15417|false|false|false|||Wound
Finding|Body Substance|Discharge Instructions|15412,15417|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|Discharge Instructions|15412,15417|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|Discharge Instructions|15412,15417|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15412,15422|false|false|false|C0886052;C1272654|Wound care management;wound care|Wound Care
Event|Activity|Discharge Instructions|15418,15422|false|false|false|C1947933|care activity|Care
Event|Event|Discharge Instructions|15418,15422|false|false|false|||Care
Finding|Finding|Discharge Instructions|15418,15422|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|15418,15422|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Discharge Instructions|15430,15434|false|false|false|||keep
Anatomy|Body Location or Region|Discharge Instructions|15439,15447|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|15439,15447|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15439,15447|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|15448,15455|false|false|false|||covered
Drug|Biomedical or Dental Material|Discharge Instructions|15468,15476|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|Discharge Instructions|15468,15476|false|false|false|||dressing
Finding|Daily or Recreational Activity|Discharge Instructions|15468,15476|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Discharge Instructions|15468,15476|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Discharge Instructions|15468,15476|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15468,15476|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|Discharge Instructions|15491,15497|false|false|false|||follow
Event|Activity|Discharge Instructions|15501,15512|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|15501,15512|false|false|false|||appointment
Anatomy|Body Location or Region|Discharge Instructions|15531,15539|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|15531,15539|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|15531,15539|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15531,15539|false|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|Discharge Instructions|15545,15549|false|false|false|C0150141|Bathing|bath
Attribute|Clinical Attribute|Discharge Instructions|15553,15557|false|false|false|C1509144|Sample pool|pool
Event|Event|Discharge Instructions|15553,15557|false|false|false|||pool
Finding|Functional Concept|Discharge Instructions|15553,15557|false|false|false|C2349200|Pool (action)|pool
Anatomy|Body Location or Region|Discharge Instructions|15565,15573|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|15565,15573|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15565,15573|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|15574,15580|false|false|false|||starts
Event|Event|Discharge Instructions|15582,15590|false|false|false|||draining
Finding|Finding|Discharge Instructions|15602,15615|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|Discharge Instructions|15608,15615|false|false|false|||surgery
Finding|Finding|Discharge Instructions|15608,15615|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|15608,15615|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|15608,15615|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15608,15615|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|Discharge Instructions|15631,15639|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|15631,15639|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|15631,15639|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15631,15639|false|false|false|C0184898|Surgical incisions|incision
Finding|Idea or Concept|Discharge Instructions|15654,15660|false|false|false|C1549636|Address type - Office|office
Finding|Finding|Discharge Instructions|15669,15673|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|15669,15673|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|15669,15673|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|15704,15710|false|false|false|||resume
Event|Event|Discharge Instructions|15711,15717|false|false|false|||taking
Event|Event|Discharge Instructions|15730,15734|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|15730,15734|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|15730,15734|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|15730,15734|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|15736,15747|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|15736,15747|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|15736,15747|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|15736,15747|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|15792,15802|false|false|false|C1524062|Additional|Additional
Attribute|Clinical Attribute|Discharge Instructions|15803,15814|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Discharge Instructions|15803,15814|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Discharge Instructions|15803,15814|false|false|false|||Medications
Finding|Intellectual Product|Discharge Instructions|15803,15814|false|false|false|C4284232|Medications|Medications
Event|Event|Discharge Instructions|15819,15826|false|false|false|||control
Attribute|Clinical Attribute|Discharge Instructions|15832,15836|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|15832,15836|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|15832,15836|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|15832,15836|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|15844,15849|false|false|false|||allow
Finding|Idea or Concept|Discharge Instructions|15863,15869|false|false|false|C0807726|refill|refill
Drug|Hazardous or Poisonous Substance|Discharge Instructions|15874,15882|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|15874,15882|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|15874,15882|false|false|false|||narcotic
Attribute|Clinical Attribute|Discharge Instructions|15883,15896|false|false|false|C2741652||prescriptions
Event|Event|Discharge Instructions|15883,15896|false|false|false|||prescriptions
Procedure|Health Care Activity|Discharge Instructions|15883,15896|false|false|false|C0033080|Prescription (procedure)|prescriptions
Event|Event|Discharge Instructions|15907,15911|false|false|false|||plan
Event|Event|Discharge Instructions|15944,15950|false|false|false|||mailed
Event|Event|Discharge Instructions|15959,15963|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|15959,15963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|15959,15963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|15959,15963|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|15967,15971|false|false|false|||pick
Event|Event|Discharge Instructions|16021,16028|false|false|false|||allowed
Event|Event|Discharge Instructions|16032,16036|false|false|false|||call
Finding|Idea or Concept|Discharge Instructions|16043,16046|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|fax
Finding|Intellectual Product|Discharge Instructions|16043,16046|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|fax
Drug|Hazardous or Poisonous Substance|Discharge Instructions|16047,16055|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|16047,16055|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|16047,16055|false|false|false|||narcotic
Attribute|Clinical Attribute|Discharge Instructions|16057,16070|false|false|false|C2741652||prescriptions
Event|Event|Discharge Instructions|16057,16070|false|false|false|||prescriptions
Procedure|Health Care Activity|Discharge Instructions|16057,16070|false|false|false|C0033080|Prescription (procedure)|prescriptions
Drug|Organic Chemical|Discharge Instructions|16071,16080|false|false|false|C0722364|Oxycontin|oxycontin
Drug|Pharmacologic Substance|Discharge Instructions|16071,16080|false|false|false|C0722364|Oxycontin|oxycontin
Event|Event|Discharge Instructions|16071,16080|false|false|false|||oxycontin
Drug|Organic Chemical|Discharge Instructions|16081,16090|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Discharge Instructions|16081,16090|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Discharge Instructions|16081,16090|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Discharge Instructions|16081,16090|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Discharge Instructions|16091,16099|false|false|false|C0086787|Percocet|percocet
Drug|Pharmacologic Substance|Discharge Instructions|16091,16099|false|false|false|C0086787|Percocet|percocet
Event|Event|Discharge Instructions|16091,16099|false|false|false|||percocet
Event|Event|Discharge Instructions|16109,16117|false|false|false|||pharmacy
Finding|Intellectual Product|Discharge Instructions|16109,16117|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Discharge Instructions|16109,16117|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|Discharge Instructions|16122,16130|false|false|false|||addition
Finding|Functional Concept|Discharge Instructions|16122,16130|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Discharge Instructions|16143,16150|false|false|false|||allowed
Event|Event|Discharge Instructions|16154,16159|false|false|false|||write
Attribute|Clinical Attribute|Discharge Instructions|16164,16168|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|16164,16168|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|16164,16168|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|16169,16180|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|16169,16180|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|16169,16180|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|16169,16180|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|16211,16218|false|false|false|||surgery
Finding|Finding|Discharge Instructions|16211,16218|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|16211,16218|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|16211,16218|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16211,16218|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|Discharge Instructions|16238,16244|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Discharge Instructions|16238,16244|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Discharge Instructions|16238,16247|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Discharge Instructions|16238,16247|false|false|false|C1522577|follow-up|Follow up
Event|Event|Discharge Instructions|16245,16247|false|false|false|||up
Event|Event|Discharge Instructions|16272,16276|false|false|false|||Call
Event|Event|Discharge Instructions|16281,16287|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|16281,16287|false|false|false|C1549636|Address type - Office|office
Event|Event|Discharge Instructions|16292,16296|false|false|false|||make
Event|Activity|Discharge Instructions|16300,16311|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|16300,16311|false|false|false|||appointment
Finding|Idea or Concept|Discharge Instructions|16335,16338|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|16335,16338|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Discharge Instructions|16347,16356|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|16347,16356|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|16347,16356|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16347,16356|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Intellectual Product|Discharge Instructions|16418,16422|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Discharge Instructions|16423,16428|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|16423,16428|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|16437,16442|false|false|false|||check
Anatomy|Body Location or Region|Discharge Instructions|16449,16457|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|16449,16457|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|16449,16457|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16449,16457|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|16458,16462|false|false|false|||take
Drug|Biomedical or Dental Material|Discharge Instructions|16463,16471|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Discharge Instructions|16463,16471|false|false|false|||baseline
Finding|Idea or Concept|Discharge Instructions|16463,16471|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Pharmacologic Substance|Discharge Instructions|16472,16478|false|false|false|C0885876|X-rays, Homeopathic Preparations|X-rays
Event|Event|Discharge Instructions|16472,16478|false|false|false|||X-rays
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|16472,16478|false|false|false|C0043309|Roentgen Rays|X-rays
Procedure|Diagnostic Procedure|Discharge Instructions|16472,16478|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|X-rays
Event|Event|Discharge Instructions|16483,16489|false|false|false|||answer
Event|Event|Discharge Instructions|16494,16503|false|false|false|||questions
Finding|Finding|Discharge Instructions|16520,16524|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|16520,16524|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|16520,16524|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|16525,16530|false|false|false|||start
Finding|Finding|Discharge Instructions|16531,16539|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Discharge Instructions|16531,16539|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Discharge Instructions|16531,16539|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Discharge Instructions|16531,16547|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16531,16547|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Discharge Instructions|16540,16547|false|false|false|||therapy
Finding|Finding|Discharge Instructions|16540,16547|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Discharge Instructions|16540,16547|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16540,16547|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Intellectual Product|Discharge Instructions|16573,16577|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Discharge Instructions|16578,16581|false|false|false|||see
Finding|Idea or Concept|Discharge Instructions|16606,16609|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|16606,16609|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Discharge Instructions|16618,16627|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|16618,16627|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|16618,16627|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16618,16627|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Finding|Discharge Instructions|16640,16644|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|16640,16644|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|16640,16644|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|16645,16652|false|false|false|||release
Finding|Functional Concept|Discharge Instructions|16645,16652|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Discharge Instructions|16645,16652|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16645,16652|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Event|Activity|Discharge Instructions|16665,16673|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|16665,16673|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|16665,16673|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|16665,16673|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|16683,16687|false|false|false|||call
Event|Event|Discharge Instructions|16692,16698|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|16692,16698|false|false|false|C1549636|Address type - Office|office
Event|Event|Discharge Instructions|16713,16718|false|false|false|||fever
Finding|Finding|Discharge Instructions|16713,16718|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|16713,16718|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|16725,16732|false|false|false|||degrees
Finding|Intellectual Product|Discharge Instructions|16725,16732|false|false|false|C0542560|Academic degree|degrees
Event|Event|Discharge Instructions|16752,16760|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|16752,16760|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|16752,16760|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16752,16760|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Injury or Poisoning|Discharge Instructions|16771,16776|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|16771,16776|false|false|false|||wound
Finding|Body Substance|Discharge Instructions|16771,16776|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|16771,16776|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|16771,16776|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Discharge Instructions|16779,16787|false|false|false|||Physical
Finding|Finding|Discharge Instructions|16779,16787|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Discharge Instructions|16779,16787|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Discharge Instructions|16779,16787|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Discharge Instructions|16779,16795|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16779,16795|false|false|false|C0949766|Physical therapy|Physical Therapy
Event|Event|Discharge Instructions|16788,16795|false|false|false|||Therapy
Finding|Finding|Discharge Instructions|16788,16795|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|Discharge Instructions|16788,16795|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16788,16795|false|false|false|C0087111|Therapeutic procedure|Therapy
Attribute|Clinical Attribute|Discharge Instructions|16799,16805|false|false|false|C0944911||Weight
Event|Event|Discharge Instructions|16799,16805|false|false|false|||Weight
Finding|Finding|Discharge Instructions|16799,16805|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|Discharge Instructions|16799,16805|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|Discharge Instructions|16799,16805|false|false|false|C1305866|Weighing patient|Weight
Finding|Finding|Discharge Instructions|16829,16833|false|false|false|C0016928|Gait|Gait
Drug|Organic Chemical|Discharge Instructions|16834,16841|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|Discharge Instructions|16834,16841|false|false|false|C4319618|Balance (substance)|balance
Event|Event|Discharge Instructions|16834,16841|false|false|false|||balance
Finding|Finding|Discharge Instructions|16834,16841|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|Discharge Instructions|16834,16841|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|Discharge Instructions|16834,16841|false|false|false|C2174421|examination of balance|balance
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16834,16850|false|false|false|C4699741|Balance training|balance training
Event|Event|Discharge Instructions|16842,16850|false|false|false|||training
Finding|Intellectual Product|Discharge Instructions|16842,16850|false|false|false|C1554161|Processing ID - Training|training
Procedure|Educational Activity|Discharge Instructions|16842,16850|false|false|false|C0040607;C0220931|Training;Training Programs|training
Event|Event|Discharge Instructions|16857,16864|false|false|false|||lifting
Procedure|Laboratory Procedure|Discharge Instructions|16869,16872|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Idea or Concept|Discharge Instructions|16878,16889|true|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Discharge Instructions|16890,16897|true|false|false|C0011119|Decompression Sickness|bending
Event|Event|Discharge Instructions|16890,16897|false|false|false|||bending
Finding|Finding|Discharge Instructions|16890,16897|true|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|Discharge Instructions|16890,16897|true|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|Discharge Instructions|16898,16906|false|false|false|||twisting
Finding|Pathologic Function|Discharge Instructions|16898,16906|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Finding|Physiologic Function|Discharge Instructions|16898,16906|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Event|Event|Discharge Instructions|16909,16919|false|false|false|||Treatments
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16909,16919|false|false|false|C0087111|Therapeutic procedure|Treatments
Event|Event|Discharge Instructions|16920,16929|false|false|false|||Frequency
Finding|Intellectual Product|Discharge Instructions|16920,16929|false|false|false|C3898838;C4321352|Frequency;How Often|Frequency
Event|Event|Discharge Instructions|16938,16942|false|false|false|||keep
Anatomy|Body Location or Region|Discharge Instructions|16947,16955|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|16947,16955|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|16947,16955|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16947,16955|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|16956,16963|false|false|false|||covered
Drug|Biomedical or Dental Material|Discharge Instructions|16975,16983|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|Discharge Instructions|16975,16983|false|false|false|||dressing
Finding|Daily or Recreational Activity|Discharge Instructions|16975,16983|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Discharge Instructions|16975,16983|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Discharge Instructions|16975,16983|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16975,16983|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|Discharge Instructions|16987,16992|false|false|false|||until
Event|Event|Discharge Instructions|16999,17005|false|false|false|||follow
Finding|Functional Concept|Discharge Instructions|16999,17005|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|16999,17005|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|16999,17008|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Discharge Instructions|16999,17008|false|false|false|C1522577|follow-up|follow up
Event|Activity|Discharge Instructions|17009,17020|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|17029,17033|false|false|false|||soak
Anatomy|Body Location or Region|Discharge Instructions|17038,17046|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|17038,17046|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|17038,17046|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17038,17046|false|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|Discharge Instructions|17052,17056|false|false|false|C0150141|Bathing|bath
Attribute|Clinical Attribute|Discharge Instructions|17061,17065|false|false|false|C1509144|Sample pool|pool
Event|Event|Discharge Instructions|17061,17065|false|false|false|||pool
Finding|Functional Concept|Discharge Instructions|17061,17065|false|false|false|C2349200|Pool (action)|pool
Anatomy|Body Location or Region|Discharge Instructions|17073,17081|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|17073,17081|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|17073,17081|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17073,17081|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|17082,17088|false|false|false|||starts
Event|Event|Discharge Instructions|17089,17097|false|false|false|||draining
Event|Event|Discharge Instructions|17116,17123|false|false|false|||surgery
Finding|Finding|Discharge Instructions|17116,17123|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|17116,17123|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|17116,17123|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17116,17123|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|Discharge Instructions|17139,17147|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|17139,17147|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|17139,17147|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|17148,17151|false|false|false|||wet
Event|Event|Discharge Instructions|17152,17156|false|false|false|||Call
Event|Event|Discharge Instructions|17161,17167|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|17161,17167|false|false|false|C1549636|Address type - Office|office
Finding|Finding|Discharge Instructions|17177,17181|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|17177,17181|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|17177,17181|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Procedure|Health Care Activity|Discharge Instructions|17185,17193|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|17194,17206|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|17194,17206|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|17194,17206|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

