CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Corgard|Drug|false|false||Corgard
null|Corgard|Drug|false|false||Corgardnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Claims attachment|Finding|false|false||attach
null|HIPAA attachments|Finding|false|false||attachnull|Fix|Phenomenon|false|false||attachnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4522245;C1415181;C1420113;C5960784;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false|C2987514|Base
null|Base|Drug|false|false|C2987514|Base
null|Dental Base|Drug|false|false|C2987514|Base
null|base - RoleClass|Drug|false|false|C2987514|Basenull|Base - General Qualifier|Finding|false|false|C2987514|Base
null|BPIFA4P gene|Finding|false|false|C2987514|Base
null|Base - RX Component Type|Finding|false|false|C2987514|Basenull|Anatomical base|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C1549548;C1705938;C1843354|Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Relevance|Modifier|false|false||RELEVANTnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|Comparison|Event|true|false||comparisonnull|Lung Volumes|Finding|false|false|C4037972;C0024109|lung volumesnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0231953;C5203106;C4522223;C1550472;C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0231953;C5203106;C4522223;C1550472;C0024115;C0740941|lungnull|Volume|LabModifier|false|false||volumesnull|IPSS-R Risk Category Low|Finding|false|false|C4037972;C0024109|low
null|IPSS Risk Category Low|Finding|false|false|C4037972;C0024109|low
null|low confidentiality|Finding|false|false|C4037972;C0024109|lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Cardiomegaly|Finding|false|false||cardiomegalynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Alignment|Modifier|false|false||alignmentnull|Wiring of sternum|Procedure|false|false|C0038293|sternal wiresnull|Sternum|Anatomy|false|false|C0407260|sternalnull|Bone Wires|Device|false|false||wiresnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Bilateral|Modifier|false|false||bilateralnull|Pleural effusion (disorder)|Finding|false|false|C0032225|pleural effusionsnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0032226;C0013687;C0032227|pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false|C0032225|effusionsnull|Aspects of signs|Finding|false|false|C0024109|Signs
null|Physical findings|Finding|false|false|C0024109|Signsnull|Manufactured sign|Device|false|false||Signsnull|Moderate - Severity of Illness Code|Finding|false|false|C0024109|moderate
null|Moderate|Finding|false|false|C0024109|moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C5201148;C1547226;C0220912;C0311392;C4522268;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Atelectasis|Finding|false|false||atelectasisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Pneumonia|Disorder|true|false||pneumonianull|Plain chest X-ray|Procedure|false|false||CXRnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|null|Procedure|false|false||wedge resectionnull|Wedge|Modifier|false|false||wedgenull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of lower lobe of lung|Anatomy|false|false|C3539671;C1428707;C2003888|lower lobenull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C3539671;C1428707|lowernull|Lower (action)|Event|false|false|C1548802;C0796494;C0225758|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false|C0225758;C0796494;C1548802|lobe
null|AKT1S1 gene|Finding|false|false|C0225758;C0796494;C1548802|lobenull|lobe|Anatomy|false|false|C2003888;C3539671;C1428707|lobenull|Small|LabModifier|false|false||Smallnull|Bilateral|Modifier|false|false||bilateralnull|effusion|Finding|false|false||effusionsnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Cardiomegaly|Finding|false|false||cardiomegalynull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Mild Severity of Illness Code|Finding|false|false|C0024109|Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Pulmonary Edema|Finding|false|false|C0024109|pulmonary edemanull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C1547225;C1717255;C0013604;C0034063;C4522268|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false|C0024109|edemanull|null|Attribute|false|false|C0024109|edemanull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4522245;C0004002;C0242192;C1121182;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|Persistence|Finding|false|false||persistencenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Adrenergic beta-Antagonists|Drug|false|false||beta blockernull|Beta adrenergic receptor antagonist (disposition)|Modifier|false|false||beta blockernull|Greek letter beta|Finding|false|false||betanull|Beta <eudicots>|Entity|false|false||betanull|Beta Distribution|LabModifier|false|false||betanull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hypotension|Finding|false|false||hypotensionnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertransaminasaemia|Finding|false|false||transaminitisnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|rosuvastatin|Drug|false|false||rosuvastatin
null|rosuvastatin|Drug|false|false||rosuvastatinnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C1420113;C5960784;C4522245;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||Alk phos
null|Alkaline Phosphatase|Drug|false|false||Alk phosnull|Alkaline phosphatase measurement|Procedure|false|false||Alk phosnull|ALK protein, human|Drug|false|false||Alk
null|ALK protein, human|Drug|false|false||Alknull|ALK protein, human|Finding|false|false||Alk
null|ALK gene|Finding|false|false||Alk
null|ALK wt Allele|Finding|false|false||Alknull|Phos <Photinae>|Entity|false|false||phosnull|Neoplasms|Disorder|false|false||Oncologynull|oncology services|Procedure|false|false||Oncologynull|oncology (field)|Title|false|false||Oncologynull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Supplement|Finding|false|false||supplementalnull|Requirement|Finding|false|false||requirementnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Pneumonia|Disorder|false|false||pneumonianull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Diuretic [APC]|Drug|false|false||DIURETIC
null|Diuretics|Drug|false|false||DIURETICnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|Male population group|Subject|false|false||man
null|Homo sapiens|Subject|false|false||man
null|Males|Subject|false|false||mannull|Mandinka Language|Entity|false|false||mannull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Tricuspid regurgitation, moderate|Finding|false|false||moderate tricuspid regurgitationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Tricuspid Valve Insufficiency|Disorder|false|false||tricuspid regurgitationnull|Tricuspid|Modifier|false|false||tricuspidnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Right Ventricular Dysfunction|Finding|false|false|C0018827|right ventricular dysfunctionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Ventricular Dysfunction|Finding|false|false|C0018827|ventricular dysfunctionnull|Heart Ventricle|Anatomy|false|false|C0242707;C3887505;C0242973|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Moderate pulmonary hypertension|Finding|false|false|C0024109|moderate pulmonary hypertensionnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Pulmonary Hypertension|Finding|false|false|C0024109|pulmonary hypertensionnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C5395246;C4522268;C0020538;C0020542|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Hypertensive disease|Disorder|false|false|C0024109|hypertensionnull|Paroxysmal|Time|false|false||paroxysmalnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidney
null|examination of kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C1561643;C0022658;C4554465;C0869841;C0012634;C0812426;C0496927;C0496892|kidney
null|Both kidneys|Anatomy|false|false|C1561643;C0022658;C4554465;C0869841;C0012634;C0812426;C0496927;C0496892|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|BaseLine dental cement|Drug|false|false||Baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||Baselinenull|Baseline|LabModifier|false|false||Baselinenull|Cerebrovascular Disorders|Disorder|false|false||cerebrovascular diseasenull|Cerebrovascular|Modifier|false|false||cerebrovascularnull|Disease|Disorder|false|false||diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Melanoma of Unknown Primary|Disorder|false|false||melanoma of unknown primarynull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumabnull|On hold|Finding|false|false||on holdnull|Hold - dosing instruction fragment|Finding|false|false||hold
null|hold - Data Operation|Finding|false|false||holdnull|Hold (action)|Event|false|false||holdnull|Hypertransaminasaemia|Finding|false|false||transaminitisnull|Concern|Finding|false|false||concernnull|Cardiotoxicity|Disorder|false|false||cardiotoxicitynull|Hypervolemia (finding)|Finding|false|false||volume overloadnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exacerbation|Finding|false|false||exacerbationnull|Pneumonia|Disorder|false|false||pneumonianull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Initially|Time|false|false||initiallynull|Coronary Care Units|Device|false|false||CCUnull|Coronary Care Units|Entity|false|false||CCUnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Flow|Phenomenon|false|false||flownull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C1550622;C1546577;C4520890;C1522019;C1272939;C0721966|nasalnull|Specimen Type - Cannula|Finding|false|false|C0028429;C1550232|cannula
null|null|Finding|false|false|C0028429;C1550232|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Precaution Code - Aggressive|Finding|false|false||aggressive
null|Aggressive behavior|Finding|false|false||aggressive
null|Risk Codes - Aggressive|Finding|false|false||aggressivenull|Aggressive course|Time|false|false||aggressivenull|Entity Risk - aggressive|Modifier|false|false||aggressivenull|Diuresis|Finding|false|false||diuresisnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Pneumonia|Disorder|false|false||pneumonianull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Floor (anatomic)|Anatomy|false|false|C5575035|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Well (answer to question)|Finding|false|false|C3714591|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Euvolemia|Finding|false|false||euvolemianull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Acute on chronic systolic heart failure|Disorder|false|false|C4037974;C0018787|Acute on chronic systolic heart failurenull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic systolic heart failure|Disorder|false|false|C4037974;C0018787|chronic systolic heart failurenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Heart Failure, Systolic|Disorder|false|false|C4037974;C0018787|systolic heart failurenull|Systole|Finding|false|false||systolicnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C1135191;C0153957;C0153500;C1135194;C0018801;C0018802;C2733492;C0795691|heart
null|Heart|Anatomy|false|false|C1135191;C0153957;C0153500;C1135194;C0018801;C0018802;C2733492;C0795691|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exacerbation|Finding|false|false||exacerbationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|null|Finding|false|false|C4037974;C0018787|history of heart failurenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0018801;C0018802;C0455531;C0680095;C0231174;C5200924;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0018801;C0018802;C0455531;C0680095;C0231174;C5200924;C0795691|heartnull|Failure (biologic function)|Finding|false|false|C4037974;C0018787|failure
null|Failure|Finding|false|false|C4037974;C0018787|failure
null|Personal failure|Finding|false|false|C4037974;C0018787|failurenull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Ischemic cardiomyopathy|Disorder|false|false||ischemic cardiomyopathynull|Ischemic|Finding|false|false||ischemicnull|Cardiomyopathies|Disorder|false|false||cardiomyopathynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Fluid Overload|Finding|false|false||fluid overload
null|Hypervolemia (finding)|Finding|false|false||fluid overloadnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Pleural effusion fluid|Finding|false|false|C0032225|pleural effusion
null|Pleural effusion (disorder)|Finding|false|false|C0032225|pleural effusion
null|null|Finding|false|false|C0032225|pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C2073625;C1253943;C0032227;C2317432;C1546613;C0013687;C0032226|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false|C0032225|effusion
null|null|Finding|false|false|C0032225|effusion
null|effusion|Finding|false|false|C0032225|effusionnull|Precipitating Factors|Attribute|false|false||Triggernull|Triggered by|Modifier|false|false||Triggernull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Exacerbation|Finding|false|false||exacerbationnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Pneumonia|Disorder|false|false|C1548802;C0225758;C0796494;C1261077|pneumonianull|Structure of left lower lobe of lung|Anatomy|false|false|C3539671;C1428707;C2003888;C1552822;C0809949;C0184666;C0032285|left lower lobenull|Table Cell Horizontal Align - left|Finding|false|false|C0225758;C1261077;C1548802|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of lower lobe of lung|Anatomy|false|false|C0809949;C0184666;C1552822;C3539671;C1428707;C2003888;C0032285|lower lobenull|Body Site Modifier - Lower|Anatomy|false|false|C0032285;C2003888;C3539671;C1428707;C1552822|lowernull|Lower (action)|Event|false|false|C1261077;C0796494;C0225758;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false|C1261077;C0225758;C0796494;C1548802|lobe
null|AKT1S1 gene|Finding|false|false|C1261077;C0225758;C0796494;C1548802|lobenull|lobe|Anatomy|false|false|C2003888;C0809949;C0184666;C3539671;C1428707;C0032285|lobenull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false|C0225758;C0796494;C1261077|admission
null|Hospital admission|Procedure|false|false|C0225758;C0796494;C1261077|admissionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Diuresis|Finding|false|false||diuresisnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Diuresis|Finding|false|false||diuresisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Euvolemia|Finding|false|false||euvolemianull|Effective|Modifier|false|false||effective
null|Effectiveness|Modifier|false|false||effectivenull|Diuresis|Finding|false|false||diuresisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unable|Finding|false|false||unablenull|Blockade|Drug|false|false||blockade
null|Blockade|Drug|false|false||blockadenull|Blocking|Finding|false|false||blockadenull|Hypotension|Finding|false|false||hypotensionnull|Left lower zone pneumonia|Disorder|false|false|C1548802;C0796494|Lower left lobe pneumonianull|Body Site Modifier - Lower|Anatomy|false|false|C0032285;C0585104;C1552822;C2003888;C3539671;C1428707|Lowernull|Lower (action)|Event|false|false|C1548802|Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Table Cell Horizontal Align - left|Finding|false|false|C0796494;C1548802|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|AKT1S1 wt Allele|Finding|false|false|C0796494;C1548802|lobe
null|AKT1S1 gene|Finding|false|false|C0796494;C1548802|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C1552822;C0585104;C0032285|lobenull|Pneumonia|Disorder|false|false|C1548802;C0796494|pneumonianull|Relationship modifier - Patient|Finding|false|false|C0225758;C0796494;C1261077|Patient
null|Specimen Type - Patient|Finding|false|false|C0225758;C0796494;C1261077|Patient
null|Mail Claim Party - Patient|Finding|false|false|C0225758;C0796494;C1261077|Patient
null|Report source - Patient|Finding|false|false|C0225758;C0796494;C1261077|Patient
null|null|Finding|false|false|C0225758;C0796494;C1261077|Patient
null|Disabled Person Code - Patient|Finding|false|false|C0225758;C0796494;C1261077|Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Evidence of (contextual qualifier)|Finding|false|false|C0796494;C1261077;C0225758|evidence ofnull|Evidence|Finding|false|false|C1548802;C1261077;C0225758;C0796494|evidencenull|Pneumonia|Disorder|false|false|C0225758;C0796494;C1261077|pneumonianull|Structure of left lower lobe of lung|Anatomy|false|false|C3887511;C1552822;C2003888;C0332120;C3539671;C1428707;C0032285;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485|left lower lobenull|Table Cell Horizontal Align - left|Finding|false|false|C1261077;C0225758|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of lower lobe of lung|Anatomy|false|false|C1578483;C1550655;C1578481;C1578486;C1578484;C1578485;C0032285;C3539671;C1428707;C3887511;C1552822;C0332120;C2003888|lower lobenull|Body Site Modifier - Lower|Anatomy|false|false|C3887511;C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0796494;C1261077;C0225758|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false|C0225758;C1261077;C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0225758;C1261077;C0796494|lobenull|lobe|Anatomy|false|false|C2003888;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485;C0032285;C0332120;C3887511;C3539671;C1428707|lobenull|Zosyn|Drug|false|false||zosyn
null|Zosyn|Drug|false|false||zosynnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Zosyn|Drug|false|false||Zosyn
null|Zosyn|Drug|false|false||Zosynnull|Total|Modifier|false|false||totalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Requirement|Finding|false|false||requirementnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Slow|Modifier|false|false||slowlynull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Supplement|Finding|false|false||supplementalnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Pleural effusion (disorder)|Finding|false|false|C0032225|Pleural effusion
null|Pleural effusion fluid|Finding|false|false|C0032225|Pleural effusion
null|null|Finding|false|false|C0032225|Pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|Pleuralnull|Pleura|Anatomy|false|false|C0032226;C2073625;C1253943;C0032227;C2317432;C1546613;C0013687|Pleuralnull|Pleural|Modifier|false|false||Pleuralnull|Effusion (substance)|Finding|false|false|C0032225|effusion
null|null|Finding|false|false|C0032225|effusion
null|effusion|Finding|false|false|C0032225|effusionnull|Bilateral|Modifier|false|false||bilateralnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false|C0032225|evidencenull|Table Cell Horizontal Align - right|Finding|false|false|C0032225|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural effusion (disorder)|Finding|false|false|C0032225|pleural effusion
null|Pleural effusion fluid|Finding|false|false|C0032225|pleural effusion
null|null|Finding|false|false|C0032225|pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C2317432;C1546613;C0013687;C1552823;C0032226;C3887511;C2073625;C1253943;C0032227|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false|C0032225|effusion
null|null|Finding|false|false|C0032225|effusion
null|effusion|Finding|false|false|C0032225|effusionnull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Fluid Overload|Finding|false|false||fluid overload
null|Hypervolemia (finding)|Finding|false|false||fluid overloadnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018801;C0018802;C0795691;C0153957;C0153500;C0680095;C0231174;C5200924|heart
null|Heart|Anatomy|false|false|C0018801;C0018802;C0795691;C0153957;C0153500;C0680095;C0231174;C5200924|heartnull|Failure (biologic function)|Finding|false|false|C4037974;C0018787|failure
null|Failure|Finding|false|false|C4037974;C0018787|failure
null|Personal failure|Finding|false|false|C4037974;C0018787|failurenull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|MDFAttributeType - Fraction|Finding|false|false||fractionnull|Fraction of|LabModifier|false|false||fractionnull|Pleural effusion (disorder)|Finding|false|false|C0032225|Pleural effusion
null|Pleural effusion fluid|Finding|false|false|C0032225|Pleural effusion
null|null|Finding|false|false|C0032225|Pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|Pleuralnull|Pleura|Anatomy|false|false|C0032226;C2317432;C1546613;C0013687;C2073625;C1253943;C0032227|Pleuralnull|Pleural|Modifier|false|false||Pleuralnull|Effusion (substance)|Finding|false|false|C0032225|effusion
null|null|Finding|false|false|C0032225|effusion
null|effusion|Finding|false|false|C0032225|effusionnull|Diuresis|Finding|false|false||diuresisnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|Thoracentesis|Procedure|false|false||thoracentesisnull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0004238;C0344434;C2926591;C0232197|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|null|Finding|false|false|C0018792|history of atrial fibrillationnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0004238;C0344434;C2926591;C0232197;C0729790|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Coronary Artery Disease|Disorder|false|false|C0205042;C0226004;C0003842;C0018787|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0205042;C0226004;C0003842;C0018787|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|Coronary arterynull|Heart|Anatomy|false|false|C1956346;C0010054|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042|artery diseasenull|Arterial system|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|artery
null|Arteries|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|arterynull|Disease|Disorder|false|false|C0205042;C0226004;C0003842|diseasenull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Low dose|LabModifier|false|false||low dosenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|rosuvastatin|Drug|false|false||rosuvastatin
null|rosuvastatin|Drug|false|false||rosuvastatinnull|Daily|Time|false|false||dailynull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Has patient|Finding|true|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cell Cycle Checkpoints|Finding|true|false||checkpointnull|Inhibitor|Drug|false|false||inhibitornull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Decision|Finding|false|false||decisionnull|Restart|Modifier|false|false||restartnull|rosuvastatin|Drug|false|false||rosuvastatin
null|rosuvastatin|Drug|false|false||rosuvastatinnull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|Chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0022658;C4554465;C0869841;C0496927;C0496892;C0812426;C1561643|kidney
null|Both kidneys|Anatomy|false|false|C0022658;C4554465;C0869841;C0496927;C0496892;C0812426;C1561643|kidneynull|Disease|Disorder|false|false||diseasenull|BaseLine dental cement|Drug|false|false||Baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||Baselinenull|Baseline|LabModifier|false|false||Baselinenull|Past Year|Time|false|false||past yearnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Thrombocytopenia|Disorder|false|false||Thrombocytopenianull|Decreased platelet count|Finding|false|false||Thrombocytopenianull|Uncertainty|Finding|false|false||Uncertainnull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|Subacute|Time|false|false||subacutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Platelets Product|Drug|false|false|C0005821|plateletsnull|Platelet count (procedure)|Procedure|false|false|C0005821|plateletsnull|Blood Platelets|Anatomy|false|false|C0443116;C0032181|plateletsnull|Concern|Finding|true|false||concernnull|Hemorrhage|Finding|true|false||bleedingnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Melanoma vaccine|Drug|false|false||Melanoma
null|Melanoma vaccine|Drug|false|false||Melanomanull|melanoma|Disorder|false|false||Melanomanull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Metastatic melanoma|Disorder|false|false||metastatic melanomanull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|On Treatment|Time|false|false||On treatmentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Iso|Entity|false|false||isonull|Toxic effect|Disorder|false|false||toxicitynull|Toxicity aspects|Modifier|false|false||toxicitynull|daunorubicin|Drug|false|false||DNR
null|daunorubicin|Drug|false|false||DNRnull|Do-Not-Resuscitate Orders|Finding|false|false||DNR
null|Do not resuscitate status|Finding|false|false||DNRnull|null|Attribute|false|false||DNRnull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|Concept Relationship|Finding|false|false||Relationship
null|Object Relationship|Finding|false|false||Relationshipnull|Relationships|Modifier|false|false||Relationshipnull|SON gene|Finding|false|false||Sonnull|Son (person)|Subject|false|false||Sonnull|Songhay Languages|Entity|false|false||Sonnull|Telephone Number|Finding|false|false||Phone numbernull|Authorization Mode - Phone|Finding|false|false||Phone
null|Visit User Code - Phone|Finding|false|false||Phone
null|Telephone Number|Finding|false|false||Phone
null|MDFAttributeType - Phone|Finding|false|false||Phonenull|Telephone|Device|false|false||Phonenull|Person location type - Phone|Modifier|false|false||Phonenull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|tamsulosin|Drug|false|false||Tamsulosin
null|tamsulosin|Drug|false|false||Tamsulosinnull|Once a day, at bedtime|Time|false|false||QHSnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10null|Coenzymes|Drug|false|false||coenzyme
null|Coenzymes|Drug|false|false||coenzymenull|AGO2 wt Allele|Finding|false|false||Q10
null|AGO2 gene|Finding|false|false||Q10null|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|Align|Drug|false|false||Align
null|Align|Drug|false|false||Alignnull|herbal medicines bifidobacterium infantis|Drug|false|false||bifidobacterium infantisnull|Bifidobacterium longum subspecies infantis|Entity|false|false||bifidobacterium infantis
null|Bifidobacterium infantis|Entity|false|false||bifidobacterium infantisnull|Bifidobacterium|Entity|false|false||bifidobacteriumnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|rosuvastatin calcium|Drug|false|false||Rosuvastatin Calcium
null|rosuvastatin calcium|Drug|false|false||Rosuvastatin Calciumnull|rosuvastatin|Drug|false|false||Rosuvastatin
null|rosuvastatin|Drug|false|false||Rosuvastatinnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Align|Drug|false|false||Align
null|Align|Drug|false|false||Alignnull|herbal medicines bifidobacterium infantis|Drug|false|false||bifidobacterium infantisnull|Bifidobacterium longum subspecies infantis|Entity|false|false||bifidobacterium infantis
null|Bifidobacterium infantis|Entity|false|false||bifidobacterium infantisnull|Bifidobacterium|Entity|false|false||bifidobacteriumnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10null|Coenzymes|Drug|false|false||coenzyme
null|Coenzymes|Drug|false|false||coenzymenull|AGO2 wt Allele|Finding|false|false||Q10
null|AGO2 gene|Finding|false|false||Q10null|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|Daily|Time|false|false||DAILYnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|tamsulosin|Drug|false|false||Tamsulosin
null|tamsulosin|Drug|false|false||Tamsulosinnull|Once a day, at bedtime|Time|false|false||QHSnull|Mineralocorticoid Receptor Antagonist [EPC]|Drug|false|false||mineralocorticoid receptor antagonist
null|Mineralocorticoid Receptor Antagonists|Drug|false|false||mineralocorticoid receptor antagonistnull|Mineralocorticoid Receptor|Drug|false|false||mineralocorticoid receptor
null|NR3C2 protein, human|Drug|false|false||mineralocorticoid receptornull|Mineralocorticoid Receptor|Finding|false|false||mineralocorticoid receptor
null|NR3C2 protein, human|Finding|false|false||mineralocorticoid receptor
null|NR3C2 gene|Finding|false|false||mineralocorticoid receptornull|Mineralocorticoid (substance)|Drug|false|false||mineralocorticoid
null|Mineralocorticoids|Drug|false|false||mineralocorticoid
null|Mineralocorticoids|Drug|false|false||mineralocorticoid
null|Mineralocorticoids|Drug|false|false||mineralocorticoid
null|Mineralocorticoid (substance)|Drug|false|false||mineralocorticoidnull|Substance with receptor antagonist mechanism of action (substance)|Drug|false|false||receptor antagonist
null|Receptor Antagonist [APC]|Drug|false|false||receptor antagonistnull|Receptor antagonist (disposition)|Modifier|false|false||receptor antagonistnull|receptor|Drug|false|false||receptornull|receptor|Finding|false|false||receptornull|Substance with receptor antagonist mechanism of action (substance)|Drug|false|false||antagonistnull|Antagonist muscle action|Finding|false|false||antagonistnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Hypotension|Finding|false|false||hypotensionnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|intolerant|Finding|false|false||intolerantnull|Greek letter beta|Finding|false|false||betanull|Beta <eudicots>|Entity|false|false||betanull|Beta Distribution|LabModifier|false|false||betanull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Hypotension|Finding|false|false||hypotensionnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary diagnosisnull|Principal diagnosis|Modifier|false|false||Primary diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Acute on chronic systolic heart failure|Disorder|false|false|C4037974;C0018787|Acute on chronic systolic heart failurenull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic systolic heart failure|Disorder|false|false|C4037974;C0018787|chronic systolic heart failurenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Heart Failure, Systolic|Disorder|false|false|C4037974;C0018787|systolic heart failurenull|Systole|Finding|false|false||systolicnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C2733492;C0795691;C0153957;C0153500;C1135194;C1135191;C0018801;C0018802|heart
null|Heart|Anatomy|false|false|C2733492;C0795691;C0153957;C0153500;C1135194;C1135191;C0018801;C0018802|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exacerbation|Finding|false|false||exacerbationnull|Left lower zone pneumonia|Disorder|false|false|C0796494;C1548802|Lower left lobe pneumonianull|Body Site Modifier - Lower|Anatomy|false|false|C1552822;C2003888;C3539671;C1428707;C0585104;C0032285|Lowernull|Lower (action)|Event|false|false|C1548802|Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Table Cell Horizontal Align - left|Finding|false|false|C1548802;C0796494|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|AKT1S1 wt Allele|Finding|false|false|C1548802;C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C1548802;C0796494|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C0585104;C0032285;C1552822|lobenull|Pneumonia|Disorder|false|false|C1548802;C0796494|pneumonianull|Bilateral pleural effusion|Disorder|false|false|C0032225|Bilateral pleural effusionnull|Bilateral|Modifier|false|false||Bilateralnull|Pleural effusion (disorder)|Finding|false|false|C0032225|pleural effusion
null|Pleural effusion fluid|Finding|false|false|C0032225|pleural effusion
null|null|Finding|false|false|C0032225|pleural effusionnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0032226;C0747635;C2073625;C1253943;C0032227;C2317432;C1546613;C0013687|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false|C0032225|effusion
null|null|Finding|false|false|C0032225|effusion
null|effusion|Finding|false|false|C0032225|effusionnull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0232197;C0344434;C2926591;C0004238|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Secondary diagnosis|Finding|false|false||Secondary diagnosisnull|null|Attribute|false|false||Secondary diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C1546481;C0012634;C1956346;C0010054;C0852949;C0010055|Coronary arterynull|Heart|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0018787;C0226004;C0003842;C0205042|artery diseasenull|Arterial system|Anatomy|false|false|C0852949;C1956346;C0010054;C0010055;C1546481;C0012634|artery
null|Arteries|Anatomy|false|false|C0852949;C1956346;C0010054;C0010055;C1546481;C0012634|arterynull|Disease|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|diseasenull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false|C0205042;C0226004;C0003842|statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Coronary Artery Bypass Surgery|Procedure|false|false|C0226004;C0003842;C0205042|CABGnull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|Chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false|C0227665;C0022646|Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false|C0227665;C0022646|Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0812426;C4554465;C0869841;C1561643;C0496927;C0496892;C1555457;C1547296;C0022658;C0012634|kidney
null|Both kidneys|Anatomy|false|false|C0812426;C4554465;C0869841;C1561643;C0496927;C0496892;C1555457;C1547296;C0022658;C0012634|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Thrombocytopenia|Disorder|false|false||Thrombocytopenianull|Decreased platelet count|Finding|false|false||Thrombocytopenianull|Metastatic melanoma|Disorder|false|false||Metastatic melanomanull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Dyspnea|Finding|false|false||short of breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|Occur (action)|Event|false|false||HAPPENEDnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false|C0024109|fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Lung|Anatomy|false|false|C1546638|lungsnull|Medical Condition|Finding|false|false||medical conditionnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|heart failure
null|Heart failure|Disorder|false|false|C4037974;C0018787|heart failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018801;C0018802;C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0018801;C0018802;C0795691;C0153957;C0153500|heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|Hardness|Modifier|false|false||hardnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false|C0004600|fluidnull|Fluid behavior|Modifier|false|false||fluidnull|null|Anatomy|false|false|C1546638|backsnull|Lung|Anatomy|false|false||lungsnull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Visit User Code - Home|Finding|false|false||HOME
null|Address type - Home|Finding|false|false||HOMEnull|home health encounter|Procedure|false|false||HOMEnull|Organization unit type - Home|Entity|false|false||HOMEnull|Person location type - Home|Modifier|false|false||HOME
null|Home environment|Modifier|false|false||HOMEnull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Appointments|Event|false|false||appointmentsnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Morning|Time|false|false||in the morningnull|Morning|Time|false|false||morningnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Heartline|Drug|false|false||HeartLine
null|Heartline|Drug|false|false||HeartLinenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|NCK-Interacting Protein with SH3 Domain|Drug|false|false||wishnull|NCKIPSD wt Allele|Finding|false|false||wish
null|NCKIPSD gene|Finding|false|false||wishnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions