 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|50,59|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|50,59|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|50,64|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|84,93|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|84,93|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|84,98|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|140,143|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|151,158|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|151,158|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Body Substance|Allergies|182,189|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|182,189|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|182,189|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Allergies|190,198|true|false|false|||recorded
Attribute|Clinical Attribute|Allergies|218,227|true|false|false|C1717415||Allergies
Event|Event|Allergies|218,227|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|218,227|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|231,236|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|Allergies|231,236|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|231,236|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|Allergies|239,248|true|false|false|||Attending
Finding|Functional Concept|Allergies|239,248|true|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|274,279|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Chief Complaint|274,279|false|false|false|C0042075|Urologic Diseases|renal
Finding|Finding|Chief Complaint|274,284|false|false|false|C0262613|Renal mass|renal mass
Event|Event|Chief Complaint|280,284|false|false|false|||mass
Finding|Finding|Chief Complaint|280,284|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Chief Complaint|280,284|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Chief Complaint|280,284|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Classification|Chief Complaint|287,292|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,323|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|314,323|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|314,323|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|314,323|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|314,323|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|314,323|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|325,330|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Chemical Viewed Structurally|Chief Complaint|344,351|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|344,363|false|false|false|C0401181|Radical nephrectomy|radical nephrectomy
Event|Event|Chief Complaint|352,363|false|false|false|||nephrectomy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|352,363|false|false|false|C0027695;C0176996|Nephrectomy;Total nephrectomy|nephrectomy
Finding|Functional Concept|History of Present Illness|446,456|false|false|false|C0444507|Incidental|incidental
Finding|Finding|History of Present Illness|446,464|false|false|false|C0743997|Incidental Findings|incidental finding
Event|Event|History of Present Illness|457,464|false|false|false|||finding
Finding|Finding|History of Present Illness|457,464|false|true|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|History of Present Illness|457,464|false|true|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Functional Concept|History of Present Illness|468,473|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|468,479|false|false|false|C0227613|Right kidney|right renal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|474,479|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|History of Present Illness|474,479|false|false|false|C0042075|Urologic Diseases|renal
Event|Event|History of Present Illness|481,485|false|false|false|||mass
Finding|Finding|History of Present Illness|481,485|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|History of Present Illness|481,485|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|History of Present Illness|481,485|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|History of Present Illness|486,496|false|false|false|||suspicious
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|501,504|false|false|false|C0152322|Structure of rostrum of corpus callosum|RCC
Disorder|Neoplastic Process|History of Present Illness|501,504|false|true|false|C0007134;C0279702;C2826323|Conventional (Clear Cell) Renal Cell Carcinoma;Refractory Cytopenia of Childhood;Renal Cell Carcinoma|RCC
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|501,504|false|true|false|C0250029|XRCC1 protein, human|RCC
Drug|Biologically Active Substance|History of Present Illness|501,504|false|true|false|C0250029|XRCC1 protein, human|RCC
Event|Event|History of Present Illness|501,504|false|false|false|||RCC
Finding|Gene or Genome|History of Present Illness|501,504|false|true|false|C1366475;C1705629|XRCC1 gene;XRCC1 wt Allele|RCC
Event|Event|History of Present Illness|515,518|false|false|false|||MRI
Finding|Gene or Genome|History of Present Illness|515,518|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|History of Present Illness|515,518|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|History of Present Illness|515,518|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Past Medical History|552,555|false|false|false|||PMH
Finding|Finding|Past Medical History|552,555|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Finding|Functional Concept|Past Medical History|569,574|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|Past Medical History|569,589|false|false|false|C0232296|Right axis deviation|right axis deviation
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|575,579|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|Past Medical History|575,579|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Finding|Finding|Past Medical History|575,589|false|false|false|C0262387|axis deviation|axis deviation
Event|Event|Past Medical History|580,589|false|false|false|||deviation
Finding|Finding|Past Medical History|580,589|false|false|false|C1705236|Protocol Deviation|deviation
Event|Event|Past Medical History|593,596|false|false|false|||PSH
Procedure|Therapeutic or Preventive Procedure|Past Medical History|598,606|false|false|false|C3841297|Cesarean|cesarean
Procedure|Therapeutic or Preventive Procedure|Past Medical History|598,614|false|false|false|C0007876|Cesarean section|cesarean section
Drug|Substance|Past Medical History|607,614|false|false|false|C1522472|section sample|section
Event|Event|Past Medical History|607,614|false|false|false|||section
Finding|Intellectual Product|Past Medical History|607,614|false|false|false|C1551341;C1552858|Act Class - Section;Html Link Type - section|section
Procedure|Laboratory Procedure|Past Medical History|607,614|false|false|false|C0700320|Sectioning technique|section
Event|Event|Past Medical History|620,624|false|false|false|||NKDA
Event|Event|Family Medical History|666,673|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|666,673|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|666,673|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|666,673|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|666,676|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|677,680|true|false|false|C0152322|Structure of rostrum of corpus callosum|RCC
Disorder|Neoplastic Process|Family Medical History|677,680|true|false|false|C0007134;C0279702;C2826323|Conventional (Clear Cell) Renal Cell Carcinoma;Refractory Cytopenia of Childhood;Renal Cell Carcinoma|RCC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|677,680|true|false|false|C0250029|XRCC1 protein, human|RCC
Drug|Biologically Active Substance|Family Medical History|677,680|true|false|false|C0250029|XRCC1 protein, human|RCC
Event|Event|Family Medical History|677,680|true|false|false|||RCC
Finding|Gene or Genome|Family Medical History|677,680|true|false|false|C1366475;C1705629|XRCC1 gene;XRCC1 wt Allele|RCC
Disorder|Disease or Syndrome|Family Medical History|714,719|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|714,719|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|714,719|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|720,723|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|728,731|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|728,731|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|728,731|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|738,741|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|738,741|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|738,741|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|738,741|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|748,751|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|748,751|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|759,762|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|759,762|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|759,762|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|759,762|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|759,762|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|766,769|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|766,769|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|766,769|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|766,769|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|766,769|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|766,769|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|775,779|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|775,779|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|795,798|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|815,820|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|815,820|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|815,820|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|815,828|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|815,828|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|815,828|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|821,828|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|821,828|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|821,828|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|821,828|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|821,828|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|821,828|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|874,878|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|874,878|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|874,878|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Body Substance|Hospital Course|916,923|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|916,923|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|916,923|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|928,936|false|false|false|||admitted
Event|Event|Hospital Course|965,977|false|false|false|||laparoscopic
Procedure|Diagnostic Procedure|Hospital Course|965,977|false|false|false|C0031150|Laparoscopy|laparoscopic
Finding|Functional Concept|Hospital Course|979,984|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Chemical Viewed Structurally|Hospital Course|985,992|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|985,1004|false|false|false|C0401181|Radical nephrectomy|radical nephrectomy
Event|Event|Hospital Course|993,1004|false|false|false|||nephrectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|993,1004|false|false|false|C0027695;C0176996|Nephrectomy;Total nephrectomy|nephrectomy
Event|Event|Hospital Course|1035,1041|true|false|false|||events
Event|Event|Hospital Course|1035,1041|true|false|false|C0441471|Event|events
Event|Event|Hospital Course|1043,1051|true|false|false|||occurred
Event|Event|Hospital Course|1060,1063|false|false|false|||see
Event|Event|Hospital Course|1064,1072|false|false|false|||dictated
Attribute|Clinical Attribute|Hospital Course|1073,1087|false|false|false|C0551628||operative note
Event|Event|Hospital Course|1083,1087|false|false|false|||note
Event|Event|Hospital Course|1092,1099|false|false|false|||details
Finding|Body Substance|Hospital Course|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Antibiotic|Hospital Course|1137,1147|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1137,1159|false|false|false|C0282638|Antibiotic Prophylaxis|antibiotic prophylaxis
Event|Event|Hospital Course|1148,1159|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1148,1159|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Body Substance|Hospital Course|1166,1173|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1166,1173|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1166,1173|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1178,1189|false|false|false|||transferred
Anatomy|Anatomical Structure|Hospital Course|1197,1202|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|1212,1216|false|false|false|||PACU
Event|Event|Hospital Course|1220,1226|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|1220,1226|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|1228,1237|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|1228,1237|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|1228,1237|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|1228,1237|false|false|false|C1705253|Logical Condition|condition
Attribute|Clinical Attribute|Hospital Course|1249,1253|false|false|false|C2598155||pain
Event|Event|Hospital Course|1249,1253|false|false|false|||pain
Finding|Functional Concept|Hospital Course|1249,1253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1249,1253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|1258,1262|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|1263,1273|false|false|false|||controlled
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1277,1280|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|Hospital Course|1277,1280|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|1277,1280|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|Hospital Course|1277,1280|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|1277,1280|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|Hospital Course|1277,1280|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|Hospital Course|1277,1280|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Event|Event|Hospital Course|1277,1280|false|false|false|||PCA
Finding|Finding|Hospital Course|1277,1280|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|Hospital Course|1277,1280|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|Hospital Course|1277,1280|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|Hospital Course|1277,1280|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1277,1280|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Drug|Organic Chemical|Hospital Course|1282,1290|false|false|false|C0720930|Hyrex Brand of Dimenhydrinate|hydrated
Drug|Pharmacologic Substance|Hospital Course|1282,1290|false|false|false|C0720930|Hyrex Brand of Dimenhydrinate|hydrated
Event|Event|Hospital Course|1282,1290|false|false|false|||hydrated
Finding|Body Substance|Hospital Course|1296,1301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|1296,1301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|1296,1301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|Hospital Course|1296,1308|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1296,1308|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|Hospital Course|1302,1308|false|false|false|||output
Finding|Conceptual Entity|Hospital Course|1302,1308|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|1302,1308|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|Hospital Course|1321,1329|false|false|false|||provided
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1352,1372|false|false|false|C0454512|Incentive spirometry|incentive spirometry
Event|Event|Hospital Course|1362,1372|false|false|false|||spirometry
Procedure|Diagnostic Procedure|Hospital Course|1362,1372|false|false|false|C0037981|Spirometry|spirometry
Event|Event|Hospital Course|1377,1388|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1377,1388|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|1404,1408|false|false|false|||once
Finding|Intellectual Product|Hospital Course|1404,1408|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Gene or Genome|Hospital Course|1414,1418|true|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Event|Event|Hospital Course|1419,1424|true|false|false|||foley
Event|Event|Hospital Course|1429,1436|true|false|false|||removed
Event|Event|Hospital Course|1445,1455|true|false|false|||difficulty
Finding|Finding|Hospital Course|1445,1455|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Drug|Chemical Viewed Functionally|Hospital Course|1457,1462|true|false|false|C0178499|Base|basic
Finding|Functional Concept|Hospital Course|1457,1462|true|false|false|C1527178|Basis - conceptual entity|basic
Procedure|Laboratory Procedure|Hospital Course|1457,1478|true|false|false|C2237045|Basic metabolic panel|basic metabolic panel
Event|Event|Hospital Course|1463,1472|true|false|false|||metabolic
Finding|Cell Function|Hospital Course|1463,1472|true|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|Hospital Course|1463,1472|true|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|Hospital Course|1463,1472|true|false|false|C4263342|Multisection metabolic|metabolic
Event|Event|Hospital Course|1473,1478|true|false|false|||panel
Finding|Idea or Concept|Hospital Course|1473,1478|true|false|false|C0441833|Groups|panel
Drug|Organic Chemical|Hospital Course|1484,1492|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|1484,1492|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|1484,1492|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|1484,1492|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|1484,1492|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Procedure|Laboratory Procedure|Hospital Course|1484,1504|false|false|false|C0009555|Complete Blood Count|complete blood count
Disorder|Disease or Syndrome|Hospital Course|1493,1498|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|1493,1498|false|false|false|||blood
Finding|Body Substance|Hospital Course|1493,1498|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Hospital Course|1493,1504|false|false|false|C0005771|Blood Cell Count|blood count
Event|Event|Hospital Course|1499,1504|false|false|false|||count
Event|Event|Hospital Course|1510,1517|false|false|false|||checked
Attribute|Clinical Attribute|Hospital Course|1519,1523|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|1519,1523|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1519,1523|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|1519,1531|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1519,1531|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Hospital Course|1524,1531|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|1524,1531|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|1524,1531|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|1524,1531|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|1524,1531|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|1524,1531|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|1524,1531|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Hospital Course|1537,1549|false|false|false|||transitioned
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1555,1558|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|Hospital Course|1555,1558|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|1555,1558|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|Hospital Course|1555,1558|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|1555,1558|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|Hospital Course|1555,1558|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|Hospital Course|1555,1558|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Event|Event|Hospital Course|1555,1558|false|false|false|||PCA
Finding|Finding|Hospital Course|1555,1558|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|Hospital Course|1555,1558|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|Hospital Course|1555,1558|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|Hospital Course|1555,1558|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1555,1558|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Anatomy|Body Space or Junction|Hospital Course|1562,1566|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|1562,1566|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|1562,1566|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|1562,1566|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Hazardous or Poisonous Substance|Hospital Course|1567,1577|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Organic Chemical|Hospital Course|1567,1577|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Pharmacologic Substance|Hospital Course|1567,1577|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Event|Event|Hospital Course|1567,1577|false|false|false|||analgesics
Drug|Food|Hospital Course|1579,1583|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1579,1583|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1579,1583|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1579,1583|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|1588,1596|false|false|false|||advanced
Finding|Classification|Hospital Course|1610,1615|false|false|false|C1710306|TOAST Classification|toast
Drug|Food|Hospital Course|1620,1628|false|false|false|C0452505|Cracker|crackers
Drug|Food|Hospital Course|1629,1633|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1629,1633|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1629,1633|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1629,1633|false|false|false|C0012159|Diet therapy|diet
Drug|Food|Hospital Course|1644,1648|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1644,1648|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1644,1648|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1644,1648|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|1653,1661|false|false|false|||advanced
Event|Event|Hospital Course|1666,1675|false|false|false|||tolerated
Event|Event|Hospital Course|1681,1690|false|false|false|||remainder
Finding|Idea or Concept|Hospital Course|1698,1706|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|1698,1713|false|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|1698,1713|false|false|false|C0489547|Hospital course|hospital course
Event|Event|Hospital Course|1707,1713|false|false|false|||course
Event|Event|Hospital Course|1718,1728|false|false|false|||relatively
Event|Event|Hospital Course|1730,1742|false|false|false|||unremarkable
Finding|Body Substance|Hospital Course|1748,1755|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1748,1755|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1748,1755|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1760,1770|false|false|false|||discharged
Finding|Intellectual Product|Hospital Course|1774,1780|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|1781,1790|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|1781,1790|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|1781,1790|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|1781,1790|false|false|false|C1705253|Logical Condition|condition
Event|Event|Hospital Course|1793,1799|true|false|false|||eating
Finding|Finding|Hospital Course|1800,1804|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|1806,1816|true|false|false|||ambulating
Event|Event|Hospital Course|1832,1839|true|false|false|||voiding
Finding|Functional Concept|Hospital Course|1832,1839|true|false|false|C0042034;C4067975|Urination;Voids|voiding
Finding|Organism Function|Hospital Course|1832,1839|true|false|false|C0042034;C4067975|Urination;Voids|voiding
Event|Event|Hospital Course|1849,1859|true|false|false|||difficulty
Finding|Finding|Hospital Course|1849,1859|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Attribute|Clinical Attribute|Hospital Course|1870,1874|true|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|1870,1874|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1870,1874|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|1870,1882|true|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1870,1882|true|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Hospital Course|1875,1882|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|1875,1882|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|1875,1882|true|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|1875,1882|true|false|false|||control
Finding|Conceptual Entity|Hospital Course|1875,1882|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|1875,1882|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|1875,1882|true|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Space or Junction|Hospital Course|1886,1890|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|1886,1890|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|1886,1890|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|1886,1890|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Hazardous or Poisonous Substance|Hospital Course|1891,1901|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Organic Chemical|Hospital Course|1891,1901|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Drug|Pharmacologic Substance|Hospital Course|1891,1901|false|false|false|C0002771;C4722089|Analgesics;Analgesics [TC]|analgesics
Event|Event|Hospital Course|1891,1901|false|false|false|||analgesics
Event|Event|Hospital Course|1906,1910|false|false|false|||exam
Finding|Functional Concept|Hospital Course|1906,1910|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|1906,1910|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Location or Region|Hospital Course|1913,1921|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Hospital Course|1913,1921|false|false|false|C0332803|Surgical wound|incision
Event|Event|Hospital Course|1913,1921|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1913,1921|false|false|false|C0184898|Surgical incisions|incision
Event|Activity|Hospital Course|1926,1931|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|Hospital Course|1926,1931|false|false|false|||clean
Event|Event|Hospital Course|1942,1948|true|false|false|||intact
Finding|Finding|Hospital Course|1942,1948|true|false|false|C1554187|Gender Status - Intact|intact
Event|Event|Hospital Course|1958,1966|true|false|false|||evidence
Finding|Idea or Concept|Hospital Course|1958,1966|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|1958,1969|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Hospital Course|1971,1979|true|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|1971,1979|true|false|false|C0018944|Hematoma|hematoma
Event|Event|Hospital Course|1980,1990|true|false|false|||collection
Finding|Conceptual Entity|Hospital Course|1980,1990|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|1980,1990|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|1980,1990|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|1980,1990|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|Hospital Course|1994,2003|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|1994,2003|true|false|false|||infection
Finding|Pathologic Function|Hospital Course|1994,2003|true|false|false|C3714514|Infection|infection
Finding|Body Substance|Hospital Course|2009,2016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2009,2016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2009,2016|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2027,2035|false|false|false|||explicit
Attribute|Clinical Attribute|Hospital Course|2037,2049|false|false|false|C3263700||instructions
Event|Event|Hospital Course|2037,2049|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|2037,2049|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|2053,2059|false|false|false|||follow
Finding|Functional Concept|Hospital Course|2053,2059|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|2053,2059|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|2053,2062|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|2053,2062|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|2060,2062|false|false|false|||up
Attribute|Clinical Attribute|Hospital Course|2097,2108|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2097,2108|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|2097,2108|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|2097,2108|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|2097,2121|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|2112,2121|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|2112,2121|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Hospital Course|2130,2139|true|false|false|||Discharge
Finding|Body Substance|Hospital Course|2130,2139|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2130,2139|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2130,2139|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2130,2139|true|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|2130,2151|true|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|2140,2151|true|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2140,2151|true|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|2140,2151|true|false|false|||Medications
Finding|Intellectual Product|Hospital Course|2140,2151|true|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|2156,2167|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Pharmacologic Substance|Hospital Course|2156,2167|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Organic Chemical|Hospital Course|2168,2181|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|2168,2181|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|2168,2181|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|2168,2181|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|2189,2195|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|2205,2212|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|Hospital Course|2205,2212|false|false|false|||Tablets
Event|Event|Hospital Course|2240,2246|false|false|false|||needed
Event|Event|Hospital Course|2251,2256|false|false|false|||break
Attribute|Clinical Attribute|Hospital Course|2265,2269|false|false|false|C2598155||pain
Event|Event|Hospital Course|2265,2269|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2265,2269|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2265,2269|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|2276,2281|false|false|false|||score
Finding|Finding|Hospital Course|2276,2281|false|false|false|C0449820|Score|score
Drug|Biomedical or Dental Material|Hospital Course|2298,2304|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|2309,2316|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|2324,2332|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|2324,2332|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|2324,2332|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|2324,2339|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|2324,2339|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|2333,2339|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|2333,2339|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|2333,2339|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|2333,2339|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|2333,2339|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|2333,2339|false|false|false|C0337443|Sodium measurement|Sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2347,2354|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|2347,2354|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|2347,2354|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2368,2375|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|2368,2375|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|2368,2375|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Mental or Behavioral Dysfunction|Hospital Course|2379,2382|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2379,2382|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|2379,2382|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|2379,2382|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|2379,2382|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|2387,2392|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|2395,2398|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|2395,2398|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2410,2417|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|2410,2417|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|2410,2417|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|2422,2429|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|2437,2446|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|2437,2446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2437,2446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2437,2446|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2437,2446|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|2437,2458|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|2437,2458|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|2447,2458|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|2447,2458|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|2447,2458|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|2460,2464|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|2460,2464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|2460,2464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|2460,2464|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|2467,2476|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|2467,2476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2467,2476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2467,2476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2467,2476|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|2467,2486|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|2477,2486|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|2477,2486|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|2477,2486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|2477,2486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|2477,2486|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2488,2493|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|2488,2493|false|false|false|C0042075|Urologic Diseases|renal
Anatomy|Cell|Hospital Course|2488,2498|false|false|false|C0553257|Epithelial cell of renal tubule|renal cell
Disorder|Neoplastic Process|Hospital Course|2488,2508|false|false|false|C0007134;C0279702|Conventional (Clear Cell) Renal Cell Carcinoma;Renal Cell Carcinoma|renal cell carcinoma
Anatomy|Cell|Hospital Course|2494,2498|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|2494,2498|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Disorder|Neoplastic Process|Hospital Course|2499,2508|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|2499,2508|false|false|false|||carcinoma
Event|Event|Discharge Condition|2533,2539|false|false|false|||stable
Finding|Intellectual Product|Discharge Condition|2533,2539|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|2576,2582|false|false|false|||shower
Event|Event|Discharge Instructions|2594,2599|true|false|false|||bathe
Event|Event|Discharge Instructions|2601,2605|true|false|false|||swim
Event|Event|Discharge Instructions|2609,2616|true|false|false|||immerse
Anatomy|Body Location or Region|Discharge Instructions|2622,2630|true|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|2622,2630|true|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|2622,2630|true|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|2622,2630|true|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|2641,2644|true|false|false|||eat
Event|Event|Discharge Instructions|2645,2657|true|false|false|||constipating
Drug|Food|Discharge Instructions|2658,2663|true|false|false|C0016452|Food|foods
Event|Event|Discharge Instructions|2658,2663|true|false|false|||foods
Drug|Food|Discharge Instructions|2679,2684|false|false|false|C0452428|Drink (dietary substance)|drink
Event|Event|Discharge Instructions|2679,2684|false|false|false|||drink
Drug|Substance|Discharge Instructions|2696,2702|true|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|2696,2702|true|false|false|||fluids
Finding|Body Substance|Discharge Instructions|2696,2702|true|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|2696,2702|true|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Discharge Instructions|2712,2716|true|false|false|||lift
Finding|Idea or Concept|Discharge Instructions|2741,2746|true|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Intellectual Product|Discharge Instructions|2741,2746|true|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Event|Event|Discharge Instructions|2747,2751|true|false|false|||book
Finding|Intellectual Product|Discharge Instructions|2747,2751|true|false|false|C0006002|Books|book
Finding|Finding|Discharge Instructions|2753,2762|false|false|false|C3845310|10 pounds|10 pounds
Event|Event|Discharge Instructions|2768,2773|false|false|false|||drive
Event|Event|Discharge Instructions|2788,2792|false|false|false|||seen
Finding|Functional Concept|Discharge Instructions|2814,2820|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|2814,2820|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|2814,2823|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|2814,2823|false|false|false|C1522577|follow-up|follow-up
Drug|Organic Chemical|Discharge Instructions|2826,2833|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|2826,2833|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|2844,2848|false|false|false|||used
Drug|Biologically Active Substance|Discharge Instructions|2863,2867|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Discharge Instructions|2863,2867|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Discharge Instructions|2863,2867|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|Discharge Instructions|2863,2867|false|false|false|C1546701|line source specimen code|line
Attribute|Clinical Attribute|Discharge Instructions|2868,2872|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|2868,2872|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|2868,2872|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|2868,2872|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|2873,2883|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|2873,2883|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|2873,2883|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Attribute|Clinical Attribute|Discharge Instructions|2894,2898|true|false|false|C2598155||pain
Event|Event|Discharge Instructions|2894,2898|true|false|false|||pain
Finding|Functional Concept|Discharge Instructions|2894,2898|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|2894,2898|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|2906,2910|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|2911,2921|true|false|false|||controlled
Drug|Organic Chemical|Discharge Instructions|2925,2932|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|2925,2932|true|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|2948,2958|false|false|false|||prescribed
Drug|Hazardous or Poisonous Substance|Discharge Instructions|2961,2969|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|2961,2969|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|2970,2974|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|2970,2974|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|2970,2974|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|2970,2974|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|2975,2985|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|2975,2985|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|2975,2985|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|2987,2990|false|false|false|||Use
Finding|Functional Concept|Discharge Instructions|2987,2990|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Finding|Intellectual Product|Discharge Instructions|2987,2990|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Event|Activity|Discharge Instructions|2994,2999|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Discharge Instructions|2994,2999|false|false|false|||place
Finding|Functional Concept|Discharge Instructions|2994,2999|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Discharge Instructions|2994,2999|false|false|false|C1533810||place
Drug|Organic Chemical|Discharge Instructions|3003,3010|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|3003,3010|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|3020,3026|true|false|false|||exceed
Event|Event|Discharge Instructions|3029,3032|true|false|false|||gms
Drug|Organic Chemical|Discharge Instructions|3036,3043|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|3036,3043|true|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|3068,3073|true|false|false|||drive
Event|Event|Discharge Instructions|3077,3082|true|false|false|||drink
Drug|Organic Chemical|Discharge Instructions|3083,3090|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|3083,3090|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Discharge Instructions|3083,3090|true|false|false|||alcohol
Finding|Intellectual Product|Discharge Instructions|3083,3090|true|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Hazardous or Poisonous Substance|Discharge Instructions|3104,3113|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Discharge Instructions|3104,3113|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Discharge Instructions|3104,3113|false|false|false|||narcotics
Event|Event|Discharge Instructions|3116,3122|false|false|false|||Resume
Finding|Functional Concept|Discharge Instructions|3116,3122|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Idea or Concept|Discharge Instructions|3116,3122|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Intellectual Product|Discharge Instructions|3116,3122|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Idea or Concept|Discharge Instructions|3135,3139|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|3135,3139|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|3135,3139|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|3140,3151|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|3140,3151|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|3140,3151|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|3140,3151|false|false|false|C4284232|Medications|medications
Event|Activity|Discharge Instructions|3160,3164|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|Discharge Instructions|3160,3164|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|Discharge Instructions|3160,3164|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Drug|Pharmacologic Substance|Discharge Instructions|3165,3170|false|false|false|C0003211;C3536840|Anti-Inflammatory Agents, Non-Steroidal|NSAID
Event|Event|Discharge Instructions|3165,3170|false|false|false|||NSAID
Drug|Organic Chemical|Discharge Instructions|3173,3180|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Discharge Instructions|3173,3180|false|false|false|C0004057|aspirin|aspirin
Event|Event|Discharge Instructions|3173,3180|false|false|false|||aspirin
Drug|Organic Chemical|Discharge Instructions|3182,3187|false|false|false|C0593507|Advil|advil
Drug|Pharmacologic Substance|Discharge Instructions|3182,3187|false|false|false|C0593507|Advil|advil
Event|Event|Discharge Instructions|3182,3187|false|false|false|||advil
Finding|Gene or Genome|Discharge Instructions|3182,3187|false|false|false|C1422473|AVIL gene|advil
Drug|Organic Chemical|Discharge Instructions|3189,3195|false|false|false|C0699203|Motrin|motrin
Drug|Pharmacologic Substance|Discharge Instructions|3189,3195|false|false|false|C0699203|Motrin|motrin
Event|Event|Discharge Instructions|3189,3195|false|false|false|||motrin
Drug|Organic Chemical|Discharge Instructions|3197,3206|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|3197,3206|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|Discharge Instructions|3197,3206|false|false|false|||ibuprofen
Event|Event|Discharge Instructions|3218,3221|false|false|false|||see
Event|Event|Discharge Instructions|3227,3236|false|false|false|||urologist
Finding|Functional Concept|Discharge Instructions|3241,3247|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|3241,3247|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|3241,3250|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|3241,3250|false|false|false|C1522577|follow-up|follow-up
Event|Event|Discharge Instructions|3265,3271|false|false|false|||fevers
Finding|Sign or Symptom|Discharge Instructions|3265,3271|false|false|false|C0015967|Fever|fevers
Event|Event|Discharge Instructions|3283,3291|false|false|false|||vomiting
Finding|Sign or Symptom|Discharge Instructions|3283,3291|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|Discharge Instructions|3296,3305|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Discharge Instructions|3296,3305|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Disorder|Disease or Syndrome|Discharge Instructions|3306,3313|false|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|3306,3313|false|false|false|||redness
Finding|Finding|Discharge Instructions|3306,3313|false|false|false|C0332575|Redness|redness
Event|Event|Discharge Instructions|3316,3324|false|false|false|||swelling
Finding|Finding|Discharge Instructions|3316,3324|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|3316,3324|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Discharge Instructions|3329,3338|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|3329,3338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|3329,3338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|3329,3338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|3329,3338|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Location or Region|Discharge Instructions|3349,3357|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|3349,3357|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|3349,3357|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3349,3357|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|3359,3363|false|false|false|||call
Event|Event|Discharge Instructions|3369,3375|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|3369,3375|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|3380,3382|false|false|false|||go
Event|Event|Discharge Instructions|3403,3407|false|false|false|||Call
Finding|Functional Concept|Discharge Instructions|3403,3407|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|Discharge Instructions|3403,3407|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|Discharge Instructions|3403,3407|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|Discharge Instructions|3403,3407|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Event|Activity|Discharge Instructions|3436,3447|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|3436,3447|false|false|false|||appointment
Event|Event|Discharge Instructions|3480,3489|true|false|false|||questions
Procedure|Health Care Activity|Discharge Instructions|3498,3506|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|3507,3519|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|3507,3519|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|3507,3519|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

