 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Finding|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|156,163|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|166,175|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|166,175|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Functional Concept|SIMPLE_SEGMENT|184,193|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|202,217|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|208,217|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|208,217|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|219,233|false|false|false|C0028756|Morbid obesity|Morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|226,233|false|false|false|C0028754|Obesity|obesity
Finding|Finding|SIMPLE_SEGMENT|226,233|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Finding|Classification|SIMPLE_SEGMENT|236,241|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|242,250|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|242,250|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|254,272|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|263,272|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|263,272|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|263,272|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|263,272|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|283,295|false|false|false|C0031150|Laparoscopy|Laparoscopic
Finding|Functional Concept|SIMPLE_SEGMENT|296,302|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|296,302|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|296,302|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|296,302|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|306,327|false|false|false|C0267725|Paraesophageal hernia|paraesophageal hernia
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|321,327|false|false|false|C0019270|Hernia|hernia
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|332,344|false|false|false|C0031150|Laparoscopy|Laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|332,368|false|false|false|C1532765|Laparoscopic adjustable gastric banding|Laparoscopic adjustable gastric band
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|356,363|false|false|false|C0038351|Stomach|gastric
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|356,368|false|false|false|C1960832|Partitioning of stomach using band|gastric band
Finding|Conceptual Entity|SIMPLE_SEGMENT|373,380|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|373,380|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|373,380|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|373,383|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|373,399|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|373,399|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|384,391|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|384,391|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|384,399|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|392,399|false|false|false|C0221423|Illness (finding)|Illness
Finding|Classification|SIMPLE_SEGMENT|417,422|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Functional Concept|SIMPLE_SEGMENT|417,422|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Intellectual Product|SIMPLE_SEGMENT|417,422|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Finding|SIMPLE_SEGMENT|417,426|false|false|false|C0441887;C2698969|Canadian Cardiovascular Society Grading of Angina Pectoris CCSGA101 Standardized Character Result Grade III;Class 3|class III
Finding|Intellectual Product|SIMPLE_SEGMENT|417,426|false|false|false|C0441887;C2698969|Canadian Cardiovascular Society Grading of Angina Pectoris CCSGA101 Standardized Character Result Grade III;Class 3|class III
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|427,441|false|false|false|C0028756|Morbid obesity|morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|434,441|false|false|false|C0028754|Obesity|obesity
Finding|Finding|SIMPLE_SEGMENT|434,441|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Finding|Idea or Concept|SIMPLE_SEGMENT|483,490|false|false|false|C1555582|Initial (abbreviation)|initial
Procedure|Health Care Activity|SIMPLE_SEGMENT|483,497|false|false|false|C3844397|Initial screening|initial screen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|491,497|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|491,497|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|551,554|false|false|false|C1305855;C1542867|Body mass index|BMI
Finding|Finding|SIMPLE_SEGMENT|551,554|false|false|false|C0578022|Finding of body mass index|BMI
Finding|Finding|SIMPLE_SEGMENT|583,587|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|629,633|false|false|false|C5890125|Loss (adaptation)|Loss
Finding|Gene or Genome|SIMPLE_SEGMENT|635,639|false|false|false|C1422329;C2681633;C3810629|KLHDC10 gene;PDLIM2 gene;PDLIM2 wt Allele|Slim
Finding|Finding|SIMPLE_SEGMENT|640,644|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|Fast
Finding|Gene or Genome|SIMPLE_SEGMENT|640,644|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|Fast
Finding|Molecular Function|SIMPLE_SEGMENT|640,644|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|Fast
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|655,662|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|SIMPLE_SEGMENT|655,662|false|false|false|C0702263|Counter brand of Terbufos|counter
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|663,673|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|663,673|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|SIMPLE_SEGMENT|663,673|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|663,673|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|663,680|false|false|false|C0443469;C1872737|PNLIP protein, human;pancreatic lipase|pancreatic lipase
Drug|Enzyme|SIMPLE_SEGMENT|663,680|false|false|false|C0443469;C1872737|PNLIP protein, human;pancreatic lipase|pancreatic lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|663,680|false|false|false|C0443469;C1872737|PNLIP protein, human;pancreatic lipase|pancreatic lipase
Finding|Gene or Genome|SIMPLE_SEGMENT|663,680|false|false|false|C1418708|PNLIP gene|pancreatic lipase
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|674,680|false|false|false|C0023764|lipase|lipase
Drug|Enzyme|SIMPLE_SEGMENT|674,680|false|false|false|C0023764|lipase|lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|674,680|false|false|false|C0023764|lipase|lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|674,680|false|false|false|C0373670|Lipase measurement|lipase
Drug|Biologically Active Substance|SIMPLE_SEGMENT|682,691|false|false|false|C1999216|Inhibitor|inhibitor
Finding|Social Behavior|SIMPLE_SEGMENT|696,702|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|SIMPLE_SEGMENT|696,702|false|false|false|C1512346|Patient Visit|visits
Finding|Finding|SIMPLE_SEGMENT|724,733|false|false|false|C3845313|20 pounds|20 pounds
Finding|Finding|SIMPLE_SEGMENT|739,745|false|false|false|C1299582|Unable|unable
Finding|Idea or Concept|SIMPLE_SEGMENT|839,846|false|false|false|C1555582|Initial (abbreviation)|initial
Procedure|Health Care Activity|SIMPLE_SEGMENT|839,853|false|false|false|C3844397|Initial screening|initial screen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|847,853|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|847,853|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Finding|Gene or Genome|SIMPLE_SEGMENT|912,915|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Idea or Concept|SIMPLE_SEGMENT|936,940|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|936,940|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Gene or Genome|SIMPLE_SEGMENT|941,944|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1016,1019|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1016,1019|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|1016,1019|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Functional Concept|SIMPLE_SEGMENT|1073,1081|false|false|false|C0017399;C0314603|Genetic;genetic aspects|genetics
Procedure|Health Care Activity|SIMPLE_SEGMENT|1073,1081|false|false|false|C1948182|genetics (procedure)|genetics
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1097,1101|false|false|false|C1998602|Meal (occasion for eating)|meal
Finding|Individual Behavior|SIMPLE_SEGMENT|1097,1109|false|false|false|C0392339|Eating routine|meal pattern
Finding|Gene or Genome|SIMPLE_SEGMENT|1130,1135|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Organic Chemical|SIMPLE_SEGMENT|1156,1169|false|false|false|C0007004;C3541972|Carbohydrate nutrients;Carbohydrates|carbohydrates
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1171,1178|false|false|false|C0043242|Superficial abrasion|grazing
Finding|Finding|SIMPLE_SEGMENT|1183,1192|false|false|false|C0013987;C0849912|Emotional;Emotions|emotional
Finding|Mental Process|SIMPLE_SEGMENT|1183,1192|false|false|false|C0013987;C0849912|Emotional;Emotions|emotional
Finding|Individual Behavior|SIMPLE_SEGMENT|1183,1199|false|false|false|C5940613|Emotional Eating|emotional eating
Finding|Organism Function|SIMPLE_SEGMENT|1193,1199|false|false|false|C0013470|Eating|eating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1203,1208|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1216,1224|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1216,1224|false|false|false|C1522704|Exercise Pain Management|exercise
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1251,1256|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Intellectual Product|SIMPLE_SEGMENT|1261,1265|false|false|false|C1561540|Transaction counts and value totals - week|week
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1295,1300|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Intellectual Product|SIMPLE_SEGMENT|1305,1309|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Intellectual Product|SIMPLE_SEGMENT|1331,1339|false|false|false|C1554161|Processing ID - Training|training
Procedure|Educational Activity|SIMPLE_SEGMENT|1331,1339|false|false|false|C0040607;C0220931|Training;Training Programs|training
Finding|Conceptual Entity|SIMPLE_SEGMENT|1353,1360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1353,1360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1353,1360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1353,1363|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1371,1380|false|false|false|C0012634|Disease|disorders
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1395,1405|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Finding|Functional Concept|SIMPLE_SEGMENT|1395,1405|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|1395,1405|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Mental Process|SIMPLE_SEGMENT|1479,1485|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1479,1492|false|false|false|C5781144||mental health
Finding|Mental Process|SIMPLE_SEGMENT|1479,1492|false|false|false|C0025353|mental health|mental health
Finding|Idea or Concept|SIMPLE_SEGMENT|1486,1492|false|false|false|C0018684|Health|health
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1522,1534|true|false|false|C0033978|Psychotropic Drugs|psychotropic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1536,1547|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1536,1547|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|1536,1547|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|1556,1560|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1556,1560|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1556,1560|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|1565,1585|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1570,1577|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1570,1577|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1570,1577|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1570,1577|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1570,1585|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1578,1585|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1578,1585|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1578,1585|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1593,1607|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|1593,1607|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1626,1638|false|false|false|C0041004|Triglycerides|triglyceride
Drug|Organic Chemical|SIMPLE_SEGMENT|1626,1638|false|false|false|C0041004|Triglycerides|triglyceride
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1640,1644|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1640,1644|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1640,1644|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1640,1644|false|false|false|C0337439|Iron measurement|iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1645,1655|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|1645,1655|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1645,1662|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1656,1662|false|false|false|C0002871|Anemia|anemia
Finding|Finding|SIMPLE_SEGMENT|1664,1673|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Finding|Mental Process|SIMPLE_SEGMENT|1664,1673|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1664,1679|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1664,1688|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1674,1679|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1680,1688|false|false|false|C0039082|Syndrome|syndrome
Finding|Functional Concept|SIMPLE_SEGMENT|1690,1698|false|false|false|C0700624|Allergic|allergic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1690,1707|false|false|false|C2607914|Allergic rhinitis (disorder)|allergic rhinitis
Finding|Gene or Genome|SIMPLE_SEGMENT|1690,1707|false|false|false|C1334103|IL13 gene|allergic rhinitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1699,1707|false|false|false|C0035455|Rhinitis|rhinitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1709,1721|false|false|false|C0013390|Dysmenorrhea|dysmenorrhea
Drug|Organic Chemical|SIMPLE_SEGMENT|1723,1730|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1723,1730|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|1723,1730|false|false|false|C0042890|Vitamins|vitamin
Drug|Hormone|SIMPLE_SEGMENT|1723,1732|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|1723,1732|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1723,1732|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|1723,1732|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1723,1732|false|false|false|C0919758|Vitamin D measurement|vitamin D
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1723,1743|false|false|false|C0042870|Vitamin D Deficiency|vitamin D deficiency
Finding|Finding|SIMPLE_SEGMENT|1723,1743|false|false|false|C5886864|Decreased circulating vitamin D concentration|vitamin D deficiency
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1733,1743|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|1733,1743|false|false|false|C0011155|Deficiency|deficiency
Finding|Intellectual Product|SIMPLE_SEGMENT|1745,1753|false|false|false|C1522634|Question (inquiry)|question
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1757,1771|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Finding|Finding|SIMPLE_SEGMENT|1777,1789|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1786,1789|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1786,1789|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|1786,1789|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1786,1789|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1786,1789|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1786,1795|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH level
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1797,1808|false|false|false|C0039730|Thalassemia|thalassemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1797,1814|false|false|false|C0702157|Thalassemia trait|thalassemia trait
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1816,1827|false|false|false|C0015695;C2711227|Fatty Liver;Steatohepatitis|fatty liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|1822,1827|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|1822,1827|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|1822,1827|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1832,1846|false|false|false|C0008350|Cholelithiasis|cholelithiasis
Finding|Functional Concept|SIMPLE_SEGMENT|1850,1860|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1850,1860|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1850,1860|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Intellectual Product|SIMPLE_SEGMENT|1861,1866|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|1861,1866|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Conceptual Entity|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1870,1880|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1889,1896|false|false|false|C0040421;C0836921|Palatine Tonsil;Tonsil|tonsils
Procedure|Health Care Activity|SIMPLE_SEGMENT|1889,1896|false|false|false|C2239123|examination of tonsils|tonsils
Finding|Functional Concept|SIMPLE_SEGMENT|1922,1933|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1922,1945|false|false|false|C0520679|Sleep Apnea, Obstructive|obstructive sleep apnea
Drug|Organic Chemical|SIMPLE_SEGMENT|1934,1939|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1934,1939|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|1934,1939|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1934,1945|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1940,1945|false|false|false|C0003578|Apnea|apnea
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1950,1966|false|false|false|C0744316|gastroesophageal|gastroesophageal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1950,1973|false|false|false|C0017168|Gastroesophageal reflux disease|gastroesophageal reflux
Finding|Finding|SIMPLE_SEGMENT|1950,1973|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|gastroesophageal reflux
Finding|Pathologic Function|SIMPLE_SEGMENT|1967,1973|false|false|false|C0232483|Reflux|reflux
Finding|Conceptual Entity|SIMPLE_SEGMENT|1986,1994|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|SIMPLE_SEGMENT|1986,1994|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Finding|SIMPLE_SEGMENT|1986,2005|false|false|false|C5419890|Completely Resolved|resolved completely
Finding|Intellectual Product|SIMPLE_SEGMENT|1995,2005|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2017,2030|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Finding|Conceptual Entity|SIMPLE_SEGMENT|2039,2046|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2039,2046|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2039,2046|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2039,2049|false|false|false|C0262926|Medical History|History of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2050,2066|false|false|false|C0032460|Polycystic Ovary Syndrome|polycystic ovary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2061,2066|false|false|false|C0029939;C0227898;C4266530|Both ovaries;Ovary;Pelvis>Ovary|ovary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2061,2066|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2061,2066|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2067,2075|false|false|false|C0039082|Syndrome|syndrome
Finding|Classification|SIMPLE_SEGMENT|2078,2084|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2078,2084|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2078,2084|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2078,2084|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2078,2092|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2085,2092|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2085,2092|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2085,2092|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2094,2101|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2094,2101|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2094,2101|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2094,2104|false|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2111,2119|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2121,2127|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2121,2127|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|SIMPLE_SEGMENT|2121,2127|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2121,2127|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2128,2137|false|false|false|C0027651;C1882062|Neoplasms;Neoplastic disease|neoplasia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2139,2144|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2139,2144|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2139,2144|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|2139,2144|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2139,2147|false|false|false|C0007102|Malignant tumor of colon|colon CA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2149,2156|false|false|false|C0205065|Ovarian|ovarian
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2165,2172|false|false|false|C1261473;C4551686|Malignant neoplasm of soft tissue;Sarcoma|sarcoma
Finding|Finding|SIMPLE_SEGMENT|2175,2183|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2175,2183|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2175,2183|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2175,2188|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2175,2188|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2184,2188|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2184,2188|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|2194,2208|false|false|false|C0740738;C1511487|CONSTITUTIONAL PROBLEM;Constitutional|Constitutional
Finding|Idea or Concept|SIMPLE_SEGMENT|2194,2208|false|false|false|C0740738;C1511487|CONSTITUTIONAL PROBLEM;Constitutional|Constitutional
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2210,2213|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2210,2213|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2210,2213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2210,2213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2210,2213|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|2210,2213|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2221,2226|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2221,2226|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2221,2226|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|2221,2226|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2221,2226|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2221,2226|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Finding|SIMPLE_SEGMENT|2231,2239|false|false|false|C1961028|Oriented to place|oriented
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2244,2251|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2244,2251|false|false|false|C1314974|Cardiac attachment|Cardiac
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2267,2272|false|false|false|C0024109|Lung|Lungs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2274,2277|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2274,2277|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2274,2277|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2280,2283|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2280,2283|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2285,2290|false|false|false|C0028754|Obesity|Obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2292,2296|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Mental Process|SIMPLE_SEGMENT|2329,2339|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2329,2339|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2344,2362|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2352,2362|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2352,2362|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Finding|SIMPLE_SEGMENT|2363,2371|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2372,2378|false|false|false|C0043250|Traumatic Wound|Wounds
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2380,2383|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2380,2383|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2384,2387|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2384,2387|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|2384,2387|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|SIMPLE_SEGMENT|2384,2387|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|2384,2387|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2384,2387|false|false|false|C0031150|Laparoscopy|lap
Drug|Organic Chemical|SIMPLE_SEGMENT|2407,2410|false|false|false|C0284559|gusperimus|dsg
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2407,2410|false|false|false|C0284559|gusperimus|dsg
Finding|Gene or Genome|SIMPLE_SEGMENT|2407,2410|false|false|false|C1414168;C5443972|DSG1 gene;DSG1 wt Allele|dsg
Finding|Finding|SIMPLE_SEGMENT|2412,2418|false|false|false|C5202796|Intensity and Distress 1|slight
Finding|Finding|SIMPLE_SEGMENT|2435,2443|false|false|false|C1704680|Staining (finding)|staining
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2435,2443|false|false|false|C0487602|Staining method|staining
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2452,2461|false|false|false|C3534099|Periwound|periwound
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2462,2470|true|false|false|C0041834|Erythema|erythema
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2471,2474|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2471,2474|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2479,2484|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2479,2484|true|false|false|C0013604|Edema|edema
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2506,2510|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2524,2529|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2524,2529|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2530,2533|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2538,2541|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2538,2541|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2538,2541|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2547,2550|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2547,2550|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2547,2550|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2547,2550|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2556,2559|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2556,2559|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2566,2569|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2566,2569|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2566,2569|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2566,2569|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2574,2577|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2574,2577|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2574,2577|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2574,2577|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2574,2577|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2583,2587|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2602,2605|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2622,2627|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2622,2627|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2628,2631|false|false|false|C0201617|Primed lymphocyte test|Plt
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|2649,2657|false|false|false|C0009924|Contrast Media|CONTRAST
Finding|Intellectual Product|SIMPLE_SEGMENT|2666,2676|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|2666,2676|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2711,2714|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2711,2714|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|2711,2714|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|SIMPLE_SEGMENT|2711,2714|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|2711,2714|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2711,2714|false|false|false|C0031150|Laparoscopy|lap
Finding|Intellectual Product|SIMPLE_SEGMENT|2728,2734|false|false|false|C0030650|Legal patent|patent
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2735,2740|false|false|false|C1955856|Surgical Stoma|stoma
Finding|Idea or Concept|SIMPLE_SEGMENT|2748,2756|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|2748,2759|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|2760,2764|true|false|false|C0332234|Leaking|leak
Finding|Intellectual Product|SIMPLE_SEGMENT|2770,2775|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|2776,2784|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2776,2791|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|2776,2791|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Sign or Symptom|SIMPLE_SEGMENT|2847,2858|false|false|false|C0278134|Absence of sensation|anaesthesia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2847,2858|false|false|false|C0002903|Anesthesia procedures|anaesthesia
Finding|Finding|SIMPLE_SEGMENT|2876,2885|false|false|false|C4738506|Operating|operating
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2914,2926|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2914,2950|false|false|false|C1532765|Laparoscopic adjustable gastric banding|laparoscopic adjustable gastric band
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2938,2945|false|false|false|C0038351|Stomach|gastric
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2938,2950|false|false|false|C1960832|Partitioning of stomach using band|gastric band
Procedure|Health Care Activity|SIMPLE_SEGMENT|2951,2960|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2951,2960|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|2966,2972|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|2966,2972|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|2966,2972|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2966,2972|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2976,2997|false|false|false|C0267725|Paraesophageal hernia|paraesophageal hernia
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2991,2997|false|false|false|C0019270|Hernia|hernia
Event|Event|SIMPLE_SEGMENT|3022,3028|false|false|false|C0441471|Event|events
Finding|Finding|SIMPLE_SEGMENT|3036,3045|false|false|false|C4738506|Operating|operating
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3067,3081|false|false|false|C0551628||operative note
Finding|Intellectual Product|SIMPLE_SEGMENT|3138,3144|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|SIMPLE_SEGMENT|3146,3150|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|SIMPLE_SEGMENT|3180,3191|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Finding|Idea or Concept|SIMPLE_SEGMENT|3180,3191|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3180,3191|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3180,3191|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Research Activity|SIMPLE_SEGMENT|3180,3191|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Finding|Body Substance|SIMPLE_SEGMENT|3217,3224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3217,3224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3217,3224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|3234,3242|false|false|false|C0277797|Apyrexial|afebrile
Finding|Intellectual Product|SIMPLE_SEGMENT|3248,3254|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|SIMPLE_SEGMENT|3256,3261|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3256,3267|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|3256,3267|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|3262,3267|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|3262,3267|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Body Substance|SIMPLE_SEGMENT|3274,3281|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3274,3281|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3274,3281|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3284,3288|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3284,3288|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3284,3288|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|3293,3297|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3314,3318|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3314,3318|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|3314,3318|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|3314,3318|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|3320,3327|false|false|false|C0723148|Roxicet|Roxicet
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3320,3327|false|false|false|C0723148|Roxicet|Roxicet
Finding|Gene or Genome|SIMPLE_SEGMENT|3328,3331|false|false|false|C1422467|CIAO3 gene|prn
Finding|Body Substance|SIMPLE_SEGMENT|3338,3345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3338,3345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3338,3345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3355,3361|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body System|SIMPLE_SEGMENT|3375,3389|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|cardiovascular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3394,3403|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3394,3403|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3394,3403|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Gene or Genome|SIMPLE_SEGMENT|3439,3443|false|false|false|C1424863|CENPJ gene|CPAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3439,3443|false|false|false|C0199451|Continuous Positive Airway Pressure|CPAP
Drug|Organic Chemical|SIMPLE_SEGMENT|3464,3469|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3464,3469|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|3464,3469|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3464,3475|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3470,3475|false|false|false|C0003578|Apnea|apnea
Finding|Body Substance|SIMPLE_SEGMENT|3482,3489|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3482,3489|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3482,3489|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3520,3525|false|false|false|C1300072|Tumor stage|stage
Finding|Classification|SIMPLE_SEGMENT|3520,3527|false|false|false|C0441766;C3840271|Stage 1;Stage level 1|stage 1
Finding|Finding|SIMPLE_SEGMENT|3520,3527|false|false|false|C0441766;C3840271|Stage 1;Stage level 1|stage 1
Drug|Food|SIMPLE_SEGMENT|3528,3532|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|3528,3532|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|3528,3532|false|false|false|C0012159|Diet therapy|diet
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3547,3550|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Finding|Gene or Genome|SIMPLE_SEGMENT|3558,3562|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Finding|Classification|SIMPLE_SEGMENT|3596,3604|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|3596,3604|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3596,3604|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|3596,3608|false|false|false|C0205160|Negative|negative for
Finding|Functional Concept|SIMPLE_SEGMENT|3609,3613|true|false|false|C0332234|Leaking|leak
Finding|Finding|SIMPLE_SEGMENT|3617,3628|true|false|false|C0028778|Obstruction|obstruction
Finding|Body Substance|SIMPLE_SEGMENT|3646,3653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3646,3653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3646,3653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Food|SIMPLE_SEGMENT|3656,3660|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|3656,3660|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|3656,3660|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3697,3702|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|3697,3704|false|false|false|C0441771|Stage level 3|stage 3
Finding|Finding|SIMPLE_SEGMENT|3709,3713|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|SIMPLE_SEGMENT|3730,3736|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|3730,3736|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|3730,3747|false|false|false|C0204708|Measuring intake and output|intake and output
Finding|Conceptual Entity|SIMPLE_SEGMENT|3741,3747|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|3741,3747|false|false|false|C3251815|Measurement of fluid output|output
Finding|Body Substance|SIMPLE_SEGMENT|3774,3779|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|3774,3779|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3774,3779|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3774,3786|false|false|false|C0232856;C0489132||Urine output
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3774,3786|false|false|false|C2094175|monitoring of urine output for fluid balance|Urine output
Finding|Conceptual Entity|SIMPLE_SEGMENT|3780,3786|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|3780,3786|false|false|false|C3251815|Measurement of fluid output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|3821,3836|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Functional Concept|SIMPLE_SEGMENT|3852,3864|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|SIMPLE_SEGMENT|3852,3872|false|false|false|C0353681|subcutaneous heparin|subcutaneous heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3852,3872|false|false|false|C0353681|subcutaneous heparin|subcutaneous heparin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3865,3872|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|3865,3872|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3865,3872|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Procedure|Health Care Activity|SIMPLE_SEGMENT|3910,3919|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3940,3950|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|3940,3950|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Body Substance|SIMPLE_SEGMENT|3983,3990|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3983,3990|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3983,3990|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4022,4026|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4022,4026|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4022,4026|false|false|false|C1553498|home health encounter|home
Finding|Gene or Genome|SIMPLE_SEGMENT|4030,4034|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Finding|Body Substance|SIMPLE_SEGMENT|4042,4049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4042,4049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4042,4049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|SIMPLE_SEGMENT|4059,4068|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4059,4068|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4059,4068|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4059,4068|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4069,4077|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|SIMPLE_SEGMENT|4069,4077|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4092,4104|false|false|false|C3263700||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4092,4104|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Mental Process|SIMPLE_SEGMENT|4111,4124|false|false|false|C0162340|Comprehension|understanding
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4140,4149|false|false|false|C4255433||agreement
Finding|Intellectual Product|SIMPLE_SEGMENT|4140,4149|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Social Behavior|SIMPLE_SEGMENT|4140,4149|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Body Substance|SIMPLE_SEGMENT|4159,4168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4159,4168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4159,4168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4159,4168|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4170,4174|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|SIMPLE_SEGMENT|4170,4174|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|4170,4174|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|4170,4174|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4258,4269|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4258,4269|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4258,4269|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|4258,4282|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4273,4282|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4301,4311|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|4301,4311|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|4301,4316|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|4312,4316|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Finding|Intellectual Product|SIMPLE_SEGMENT|4356,4369|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4356,4369|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|SIMPLE_SEGMENT|4374,4387|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4374,4387|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|4374,4387|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4390,4398|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4401,4404|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|4418,4431|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4418,4431|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Vitamin|SIMPLE_SEGMENT|4418,4431|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4418,4431|false|false|false|C0201898|Ascorbic acid measurement|Ascorbic Acid
Drug|Organic Chemical|SIMPLE_SEGMENT|4452,4467|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4452,4467|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Vitamin|SIMPLE_SEGMENT|4452,4467|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Organic Chemical|SIMPLE_SEGMENT|4452,4480|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4452,4480|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Vitamin|SIMPLE_SEGMENT|4452,4480|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Organic Chemical|SIMPLE_SEGMENT|4469,4476|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4469,4476|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|4469,4476|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|4469,4479|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4469,4479|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|4469,4479|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4497,4501|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4497,4501|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|4497,4501|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|4497,4501|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|SIMPLE_SEGMENT|4512,4527|false|false|false|C0056732|cyclobenzaprine|Cyclobenzaprine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4512,4527|false|false|false|C0056732|cyclobenzaprine|Cyclobenzaprine
Finding|Gene or Genome|SIMPLE_SEGMENT|4542,4545|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4546,4552|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|4546,4552|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|SIMPLE_SEGMENT|4546,4559|false|false|false|C0037763|Spasm|muscle spasms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4553,4559|false|false|false|C0037763|Spasm|spasms
Finding|Body Substance|SIMPLE_SEGMENT|4564,4573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4564,4573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4564,4573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4564,4573|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|4564,4585|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4574,4585|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4574,4585|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4574,4585|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|4590,4599|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4590,4599|false|false|false|C0030049|oxycodone|OxycoDONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4590,4599|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4590,4613|false|false|false|C0717368|acetaminophen / oxycodone|OxycoDONE-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|4600,4613|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4600,4613|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4600,4613|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4614,4620|false|false|false|C0678430|Elixir|Elixir
Finding|Gene or Genome|SIMPLE_SEGMENT|4635,4638|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4639,4643|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|4639,4643|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4639,4643|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|4649,4658|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4649,4658|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4649,4658|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4649,4672|false|false|false|C0717368|acetaminophen / oxycodone|oxycodone-acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|4659,4672|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4659,4672|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4659,4672|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|4674,4681|false|false|false|C0723148|Roxicet|Roxicet
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4674,4681|false|false|false|C0723148|Roxicet|Roxicet
Finding|Functional Concept|SIMPLE_SEGMENT|4708,4716|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4711,4716|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4711,4716|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|4760,4767|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|4774,4782|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4774,4782|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|4774,4789|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4774,4789|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4783,4789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4783,4789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4783,4789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|4783,4789|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4783,4789|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4791,4797|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|SIMPLE_SEGMENT|4791,4797|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Finding|Finding|SIMPLE_SEGMENT|4791,4797|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4791,4797|false|false|false|C0301571|Liquid diet|Liquid
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4809,4812|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4809,4812|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4809,4812|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4809,4812|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4813,4816|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|4817,4829|false|false|false|C0009806|Constipation|Constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|4835,4843|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4835,4843|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|4835,4850|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4835,4850|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4844,4850|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4844,4850|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4844,4850|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|4844,4850|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4844,4850|false|false|false|C0337443|Sodium measurement|sodium
Finding|Functional Concept|SIMPLE_SEGMENT|4869,4877|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4872,4877|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4872,4877|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|4886,4889|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|4886,4889|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|4890,4894|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|4890,4894|false|false|false|C2828567|PRSS30P gene|Disp
Finding|Idea or Concept|SIMPLE_SEGMENT|4913,4920|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|4927,4940|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4927,4940|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Vitamin|SIMPLE_SEGMENT|4927,4940|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4927,4940|false|false|false|C0201898|Ascorbic acid measurement|Ascorbic Acid
Drug|Organic Chemical|SIMPLE_SEGMENT|4961,4976|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4961,4976|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Vitamin|SIMPLE_SEGMENT|4961,4976|false|false|false|C0008318|cholecalciferol|cholecalciferol
Drug|Organic Chemical|SIMPLE_SEGMENT|4961,4989|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4961,4989|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Vitamin|SIMPLE_SEGMENT|4961,4989|false|false|false|C0008318|cholecalciferol|cholecalciferol (vitamin D3)
Drug|Organic Chemical|SIMPLE_SEGMENT|4978,4985|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4978,4985|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|4978,4985|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|4978,4988|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4978,4988|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|4978,4988|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5006,5010|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5006,5010|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|5006,5010|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5006,5010|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|SIMPLE_SEGMENT|5021,5034|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5021,5034|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|5021,5034|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5037,5045|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5048,5051|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Body Substance|SIMPLE_SEGMENT|5065,5074|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5065,5074|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5065,5074|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5065,5074|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5065,5086|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|5065,5086|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5075,5086|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|5075,5086|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|5088,5092|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|5088,5092|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5088,5092|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|SIMPLE_SEGMENT|5095,5104|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5095,5104|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5095,5104|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5095,5104|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5095,5114|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5105,5114|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|5105,5114|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|5105,5114|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5105,5114|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5116,5130|false|false|false|C0028756|Morbid obesity|Morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5123,5130|false|false|false|C0028754|Obesity|obesity
Finding|Finding|SIMPLE_SEGMENT|5123,5130|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Finding|Functional Concept|SIMPLE_SEGMENT|5131,5142|false|false|false|C0549186|Obstructed|Obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5131,5154|false|false|false|C0520679|Sleep Apnea, Obstructive|Obstructive sleep apnea
Drug|Organic Chemical|SIMPLE_SEGMENT|5143,5148|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5143,5148|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|5143,5148|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5143,5154|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5149,5154|false|false|false|C0003578|Apnea|apnea
Finding|Body Substance|SIMPLE_SEGMENT|5158,5167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5158,5167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5158,5167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5158,5167|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5168,5177|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5168,5177|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|5168,5177|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|5179,5185|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5179,5192|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|5179,5192|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5186,5192|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|5186,5192|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|5194,5199|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|5204,5212|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5214,5236|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|5214,5236|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|5223,5236|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|5223,5236|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5238,5243|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|5238,5243|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5238,5243|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|5238,5243|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|5238,5243|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|5238,5243|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|5248,5259|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|5261,5269|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5261,5269|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|5261,5269|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5270,5276|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|5270,5276|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|5278,5288|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|5278,5288|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|5278,5288|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|5278,5288|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|5291,5302|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|5291,5302|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|5307,5316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5307,5316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5307,5316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5307,5316|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5307,5329|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5307,5329|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|5307,5329|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5317,5329|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5317,5329|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Body Substance|SIMPLE_SEGMENT|5331,5340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5331,5340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5331,5340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5331,5340|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5331,5353|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5331,5353|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|5331,5353|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5341,5353|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5341,5353|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5372,5379|false|false|false|C5444295||surgeon
Finding|Finding|SIMPLE_SEGMENT|5398,5407|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|5398,5407|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|5398,5407|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|5398,5407|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5398,5407|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|5398,5407|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|5408,5418|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Finding|Finding|SIMPLE_SEGMENT|5436,5441|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|5436,5441|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5463,5468|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|5463,5468|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5463,5473|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5463,5473|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5469,5473|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5469,5473|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5469,5473|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5475,5494|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|5475,5494|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|5488,5494|false|false|false|C0225386|Breath|breath
Finding|Finding|SIMPLE_SEGMENT|5496,5502|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5496,5502|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5503,5512|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|5503,5517|false|true|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5513,5517|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5513,5517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5513,5517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5520,5524|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5520,5524|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5520,5524|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5544,5548|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5544,5548|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5544,5548|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5549,5559|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5549,5559|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|SIMPLE_SEGMENT|5561,5567|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5561,5567|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|SIMPLE_SEGMENT|5561,5574|false|false|false|C5936462|Severe nausea|severe nausea
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5568,5574|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5568,5574|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5579,5587|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|SIMPLE_SEGMENT|5589,5595|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5589,5595|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5596,5605|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|5596,5614|false|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|abdominal bloating
Finding|Sign or Symptom|SIMPLE_SEGMENT|5596,5614|false|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|abdominal bloating
Finding|Finding|SIMPLE_SEGMENT|5606,5614|false|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|bloating
Finding|Sign or Symptom|SIMPLE_SEGMENT|5606,5614|false|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|bloating
Finding|Organism Function|SIMPLE_SEGMENT|5649,5657|false|false|false|C0037361|Smell Perception|smelling
Finding|Body Substance|SIMPLE_SEGMENT|5670,5678|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|5670,5678|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5670,5678|false|false|false|C0013103|Drainage procedure|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5689,5698|false|false|false|C0184898|Surgical incisions|incisions
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5700,5707|false|false|false|C0041834|Erythema|redness
Finding|Finding|SIMPLE_SEGMENT|5700,5707|false|false|false|C0332575|Redness|redness
Finding|Finding|SIMPLE_SEGMENT|5712,5720|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|5712,5720|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5733,5742|false|false|false|C0184898|Surgical incisions|incisions
Finding|Functional Concept|SIMPLE_SEGMENT|5757,5765|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|5757,5765|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Food|SIMPLE_SEGMENT|5797,5801|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Finding|Functional Concept|SIMPLE_SEGMENT|5797,5801|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5797,5801|false|false|false|C0012159|Diet therapy|Diet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5811,5816|false|false|false|C1300072|Tumor stage|Stage
Drug|Food|SIMPLE_SEGMENT|5821,5825|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|5821,5825|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5821,5825|false|false|false|C0012159|Diet therapy|diet
Finding|Functional Concept|SIMPLE_SEGMENT|5837,5843|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5837,5843|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5837,5846|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5837,5846|false|false|false|C1522577|follow-up|follow up
Event|Activity|SIMPLE_SEGMENT|5847,5858|false|false|false|C0003629|Appointments|appointment
Drug|Food|SIMPLE_SEGMENT|5881,5885|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|5881,5885|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5881,5885|false|false|false|C0012159|Diet therapy|diet
Drug|Organic Chemical|SIMPLE_SEGMENT|5909,5914|false|true|false|C4047917|Cereal plant straw|straw
Finding|Finding|SIMPLE_SEGMENT|5918,5922|false|false|false|C0024888;C0699816;C1549534|Chew (administration method);Chewing;Does chew (finding)|chew
Finding|Functional Concept|SIMPLE_SEGMENT|5918,5922|false|false|false|C0024888;C0699816;C1549534|Chew (administration method);Chewing;Does chew (finding)|chew
Finding|Organism Function|SIMPLE_SEGMENT|5918,5922|false|false|false|C0024888;C0699816;C1549534|Chew (administration method);Chewing;Does chew (finding)|chew
Anatomy|Tissue|SIMPLE_SEGMENT|5924,5927|false|false|false|C0017562|Gingiva|gum
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5924,5927|false|false|false|C0812395;C1378701|Gum Dose Form;Gum as an ingredient|gum
Finding|Gene or Genome|SIMPLE_SEGMENT|5924,5927|false|false|false|C1825233;C5444202|OTULIN gene;OTULIN wt Allele|gum
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5930,5940|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5930,5940|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5941,5953|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5941,5953|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Idea or Concept|SIMPLE_SEGMENT|5967,5971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5967,5971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5967,5971|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6016,6031|false|false|false|C0056732|cyclobenzaprine|cyclobenzaprine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6016,6031|false|false|false|C0056732|cyclobenzaprine|cyclobenzaprine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6045,6049|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6045,6049|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6045,6049|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6063,6068|false|false|false|C0185060|Crushing (procedure)|CRUSH
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6073,6078|false|false|false|C0994475|Pills|PILLS
Finding|Finding|SIMPLE_SEGMENT|6106,6109|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6106,6109|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6106,6121|false|false|false|C1718097|New medications|new medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6110,6121|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6110,6121|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6110,6121|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6155,6166|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6155,6166|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6155,6166|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6180,6184|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6180,6184|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6180,6184|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Activity|SIMPLE_SEGMENT|6196,6205|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|6196,6205|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6196,6205|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6213,6224|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6213,6224|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6213,6224|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|6239,6245|false|false|false|C0013144|Drowsiness|drowsy
Finding|Functional Concept|SIMPLE_SEGMENT|6263,6270|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|SIMPLE_SEGMENT|6263,6273|false|false|false|C5420000|Ability Question|ability to
Finding|Functional Concept|SIMPLE_SEGMENT|6282,6287|false|false|false|C1513492|motor movement|motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6288,6295|false|false|false|C0042444|Drug vehicle|vehicle
Finding|Functional Concept|SIMPLE_SEGMENT|6299,6306|false|false|false|C3242339|operate|operate
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6308,6317|false|false|false|C0337246|Contact with machinery|machinery
Event|Activity|SIMPLE_SEGMENT|6353,6363|false|false|false|C0441655|Activities|activities
Finding|Finding|SIMPLE_SEGMENT|6353,6363|false|false|false|C2239122|activities (history)|activities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6384,6395|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6384,6395|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6384,6395|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|6435,6443|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6435,6443|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|6444,6456|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6444,6456|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|SIMPLE_SEGMENT|6444,6456|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6463,6471|false|false|false|C0026162|Minerals|minerals
Drug|Organic Chemical|SIMPLE_SEGMENT|6482,6490|true|false|false|C0042890;C3540032;C3714649|VITAMINS [VA Class];Vitamin IV solution additives;Vitamins|vitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6482,6490|true|false|false|C0042890;C3540032;C3714649|VITAMINS [VA Class];Vitamin IV solution additives;Vitamins|vitamins
Drug|Vitamin|SIMPLE_SEGMENT|6482,6490|true|false|false|C0042890;C3540032;C3714649|VITAMINS [VA Class];Vitamin IV solution additives;Vitamins|vitamins
Finding|Body Substance|SIMPLE_SEGMENT|6513,6518|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|6513,6527|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6513,6527|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Organic Chemical|SIMPLE_SEGMENT|6529,6535|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6529,6535|false|false|false|C0282139|Colace|Colace
Finding|Sign or Symptom|SIMPLE_SEGMENT|6554,6566|false|false|false|C0009806|Constipation|constipation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6607,6612|false|false|false|C0021853|Intestines|bowel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6643,6649|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6665,6682|false|true|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6684,6689|false|false|false|C0013227|Pharmaceutical Preparations|drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6684,6689|false|false|false|C3687832|Drugs - dental services|drugs
Drug|Organic Chemical|SIMPLE_SEGMENT|6704,6713|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6704,6713|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Organic Chemical|SIMPLE_SEGMENT|6715,6721|false|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6715,6721|false|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|SIMPLE_SEGMENT|6723,6728|false|false|false|C0718343|Aleve|Aleve
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6723,6728|false|false|false|C0718343|Aleve|Aleve
Drug|Organic Chemical|SIMPLE_SEGMENT|6730,6736|false|false|false|C0699205|Nuprin|Nuprin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6730,6736|false|false|false|C0699205|Nuprin|Nuprin
Drug|Organic Chemical|SIMPLE_SEGMENT|6742,6750|false|false|false|C0027396|naproxen|Naproxen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6742,6750|false|false|false|C0027396|naproxen|Naproxen
Finding|Pathologic Function|SIMPLE_SEGMENT|6776,6784|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|6789,6795|false|false|false|C0041582|Ulcer|ulcers
Anatomy|Body System|SIMPLE_SEGMENT|6805,6814|false|false|false|C0012240|Gastrointestinal system|digestive
Finding|Organism Function|SIMPLE_SEGMENT|6805,6814|false|false|false|C0012238|Digestion|digestive
Anatomy|Body System|SIMPLE_SEGMENT|6805,6821|false|false|false|C0012240|Gastrointestinal system|digestive system
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6815,6821|false|false|false|C5671121|System (basic dose form)|system
Finding|Functional Concept|SIMPLE_SEGMENT|6815,6821|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Activity|SIMPLE_SEGMENT|6824,6832|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6824,6832|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|6824,6832|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Activity|SIMPLE_SEGMENT|6843,6850|true|false|false|C0206244|Lifting|lifting
Finding|Finding|SIMPLE_SEGMENT|6900,6908|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6900,6908|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6900,6917|false|false|false|C1513375|Moderate Exercise|moderate exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6909,6917|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6909,6917|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Functional Concept|SIMPLE_SEGMENT|6926,6936|false|false|false|C5556474|Discretion|discretion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6941,6950|false|false|false|C0000726|Abdomen|abdominal
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6952,6961|false|false|false|C0015259|Exercise|exercises
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6952,6961|false|false|false|C0452240|Physical therapy exercises|exercises
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6964,6969|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Finding|Body Substance|SIMPLE_SEGMENT|6964,6969|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|6964,6969|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|6964,6969|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6964,6974|false|false|false|C0886052;C1272654|Wound care management;wound care|Wound Care
Event|Activity|SIMPLE_SEGMENT|6970,6974|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|6970,6974|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|6970,6974|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Gene or Genome|SIMPLE_SEGMENT|6995,6998|true|false|false|C1421225|TUB gene|tub
Procedure|Health Care Activity|SIMPLE_SEGMENT|6999,7004|true|false|false|C0150141|Bathing|baths
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7008,7016|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|SIMPLE_SEGMENT|7008,7016|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Idea or Concept|SIMPLE_SEGMENT|7031,7036|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Body Substance|SIMPLE_SEGMENT|7037,7045|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|7037,7045|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7037,7045|false|false|false|C0013103|Drainage procedure|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7056,7065|false|false|false|C0184898|Surgical incisions|incisions
Finding|Functional Concept|SIMPLE_SEGMENT|7067,7072|false|false|false|C1999244||cover
Event|Activity|SIMPLE_SEGMENT|7079,7084|false|false|false|C1947930|Cleaning (activity)|clean
Finding|Finding|SIMPLE_SEGMENT|7139,7142|false|false|false|C5939094|Own|own
Finding|Finding|SIMPLE_SEGMENT|7189,7202|false|false|false|C0241311|post operative (finding)|after surgery
Finding|Finding|SIMPLE_SEGMENT|7195,7202|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|7195,7202|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|7195,7202|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7195,7202|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Intellectual Product|SIMPLE_SEGMENT|7220,7226|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7249,7253|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7249,7253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7249,7253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|7255,7263|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|7255,7263|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7266,7273|false|false|false|C0041834|Erythema|redness
Finding|Finding|SIMPLE_SEGMENT|7266,7273|false|false|false|C0332575|Redness|redness
Finding|Body Substance|SIMPLE_SEGMENT|7278,7286|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|7278,7286|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7278,7286|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7296,7304|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7296,7304|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7296,7304|false|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|SIMPLE_SEGMENT|7316,7324|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7325,7337|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7325,7337|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

