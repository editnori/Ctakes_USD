 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|176,183|false|false|false|C0591292|Corgard|Corgard
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|176,183|false|false|false|C0591292|Corgard|Corgard
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Classification|SIMPLE_SEGMENT|210,215|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|216,224|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|216,224|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|228,246|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|237,246|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|237,246|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|237,246|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|237,246|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|237,246|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|254,260|false|false|false|||attach
Finding|Intellectual Product|SIMPLE_SEGMENT|254,260|false|false|false|C1314972;C2598091|Claims attachment;HIPAA attachments|attach
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|254,260|false|false|false|C3714578|Fix|attach
Procedure|Health Care Activity|SIMPLE_SEGMENT|282,291|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|292,296|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|292,296|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|326,331|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|326,331|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|326,331|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|332,335|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|342,345|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|342,345|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|342,345|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|352,355|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|352,355|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|352,355|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|352,355|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|362,365|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|362,365|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|373,376|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|373,376|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|373,376|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|373,376|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|373,376|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|381,384|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|381,384|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|381,384|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|381,384|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|381,384|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|381,384|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|390,394|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|390,394|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|423,426|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|443,448|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|443,448|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|443,448|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|453,456|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|453,456|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|453,456|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|479,484|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|479,484|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|479,484|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|479,492|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|479,492|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|479,492|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|485,492|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|485,492|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|485,492|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|485,492|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|485,492|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|485,492|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|540,544|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|540,544|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|540,544|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|569,574|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|569,574|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|569,574|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|575,578|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|575,578|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|575,578|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|575,578|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|575,578|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|575,578|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|575,578|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|575,578|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|583,586|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|583,586|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|583,586|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|583,586|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|583,586|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|583,586|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|583,586|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|591,598|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|591,598|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|628,633|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|628,633|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|628,633|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|650,655|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|650,655|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|650,655|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|650,663|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|656,663|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|656,663|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|656,663|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|656,663|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|656,663|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|656,663|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|656,663|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|656,663|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|696,701|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|696,701|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|696,701|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|706,709|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|706,709|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|706,709|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|706,709|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|714,718|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|714,718|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|743,747|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|743,747|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|743,747|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|743,747|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|743,747|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|743,747|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Event|Event|SIMPLE_SEGMENT|764,768|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|764,768|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|797,802|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|797,802|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|797,802|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|808,815|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|808,815|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|808,815|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|826,829|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|826,829|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Activity|SIMPLE_SEGMENT|838,848|true|false|false|C1707455|Comparison|comparison
Event|Event|SIMPLE_SEGMENT|838,848|false|false|false|||comparison
Anatomy|Body Location or Region|SIMPLE_SEGMENT|855,859|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|855,859|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|855,859|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|855,859|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|855,867|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|SIMPLE_SEGMENT|860,867|false|false|false|||volumes
Event|Event|SIMPLE_SEGMENT|872,875|false|false|false|||low
Finding|Finding|SIMPLE_SEGMENT|872,875|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|872,875|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|878,886|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|878,886|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|887,899|false|false|false|||cardiomegaly
Finding|Finding|SIMPLE_SEGMENT|887,899|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|SIMPLE_SEGMENT|904,911|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|904,911|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|904,911|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|921,930|false|false|false|||alignment
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|938,945|false|false|false|C0038293|Sternum|sternal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|938,951|false|false|false|C0407260|Wiring of sternum|sternal wires
Event|Event|SIMPLE_SEGMENT|946,951|false|false|false|||wires
Event|Event|SIMPLE_SEGMENT|958,962|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|958,962|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Intellectual Product|SIMPLE_SEGMENT|966,970|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Tissue|SIMPLE_SEGMENT|981,988|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|981,988|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|981,998|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|989,998|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|989,998|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|1001,1006|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|1001,1006|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|1001,1006|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Finding|SIMPLE_SEGMENT|1010,1018|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|1010,1018|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1019,1028|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1019,1028|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1019,1028|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1030,1035|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1030,1035|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1030,1035|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1051,1062|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|1051,1062|false|false|false|C0004144|Atelectasis|atelectasis
Event|Event|SIMPLE_SEGMENT|1067,1075|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|1067,1075|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1067,1078|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1079,1088|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1079,1088|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|1092,1095|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1092,1095|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1111,1117|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1111,1117|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|1131,1138|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1131,1138|false|false|false|C0392747|Changing|changes
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1149,1164|false|false|false|C0184909||wedge resection
Event|Event|SIMPLE_SEGMENT|1155,1164|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1155,1164|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Finding|Functional Concept|SIMPLE_SEGMENT|1170,1175|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1177,1182|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1177,1182|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1177,1187|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1183,1187|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|1183,1187|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|1206,1215|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|1206,1215|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|1216,1221|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|1216,1221|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|1235,1239|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|1235,1239|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|1245,1254|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|1245,1254|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|1274,1284|false|false|false|||silhouette
Event|Event|SIMPLE_SEGMENT|1288,1294|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1288,1294|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|1307,1315|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|1307,1315|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|1316,1328|false|false|false|||cardiomegaly
Finding|Finding|SIMPLE_SEGMENT|1316,1328|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1334,1346|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|1334,1346|false|false|false|||pneumothorax
Finding|Intellectual Product|SIMPLE_SEGMENT|1349,1353|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1354,1363|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1354,1363|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1354,1363|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|1354,1369|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1364,1369|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1364,1369|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1364,1369|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1374,1383|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|1374,1383|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|1397,1401|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1397,1401|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1435,1440|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1435,1440|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1435,1440|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|1441,1444|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1449,1452|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1449,1452|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1449,1452|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1459,1462|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1459,1462|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1459,1462|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1459,1462|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1469,1472|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1469,1472|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|1480,1483|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|1480,1483|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1480,1483|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1480,1483|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1480,1483|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|1487,1490|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1487,1490|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|1487,1490|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|1487,1490|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|1487,1490|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1487,1490|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|1496,1500|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1496,1500|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1529,1532|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1549,1554|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1549,1554|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1549,1554|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|1549,1562|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1549,1562|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1549,1562|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1555,1562|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|1555,1562|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1555,1562|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|1555,1562|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1555,1562|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1555,1562|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1607,1611|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1607,1611|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1607,1611|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1636,1641|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1636,1641|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1636,1641|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1642,1645|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1642,1645|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|1642,1645|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|1642,1645|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|1642,1645|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|1642,1645|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|1642,1645|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1642,1645|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1649,1652|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1649,1652|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1649,1652|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1649,1652|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|1649,1652|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|1649,1652|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|1649,1652|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1660,1663|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|1660,1663|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|1660,1663|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|1660,1663|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1660,1663|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1669,1676|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|1669,1676|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1706,1711|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1706,1711|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1706,1711|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1706,1719|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1712,1719|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1712,1719|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1712,1719|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1712,1719|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|1712,1719|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|1712,1719|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|1712,1719|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1712,1719|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Intellectual Product|SIMPLE_SEGMENT|1742,1747|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|1748,1756|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1748,1763|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|1748,1763|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|1765,1777|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|1778,1784|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|1810,1818|false|false|false|||Consider
Drug|Organic Chemical|SIMPLE_SEGMENT|1833,1843|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1833,1843|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|1833,1843|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1833,1843|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|1850,1861|false|false|false|||persistence
Finding|Mental Process|SIMPLE_SEGMENT|1850,1861|false|false|false|C0546816|Persistence|persistence
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1882,1892|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|1882,1892|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|1882,1892|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|1896,1904|false|false|false|||Consider
Event|Event|SIMPLE_SEGMENT|1905,1913|false|false|false|||starting
Finding|Intellectual Product|SIMPLE_SEGMENT|1914,1918|false|false|false|C0439096|Greek letter beta|beta
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1914,1926|false|false|false|C0001645|Adrenergic beta-Antagonists|beta blocker
Event|Event|SIMPLE_SEGMENT|1919,1926|false|false|false|||blocker
Event|Event|SIMPLE_SEGMENT|1937,1941|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1937,1941|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|1945,1953|false|false|false|||tolerate
Finding|Body Substance|SIMPLE_SEGMENT|1956,1963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1956,1963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1956,1963|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1983,1991|false|false|false|||tolerate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1997,2007|false|true|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|1997,2007|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|1997,2007|false|true|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2018,2031|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|SIMPLE_SEGMENT|2018,2031|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2018,2031|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|SIMPLE_SEGMENT|2018,2031|false|false|false|||pembrolizumab
Event|Event|SIMPLE_SEGMENT|2033,2042|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2033,2042|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|2056,2063|false|false|false|||patient
Finding|Body Substance|SIMPLE_SEGMENT|2056,2063|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2056,2063|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2056,2063|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|2056,2067|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|2073,2076|false|false|false|||off
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2081,2094|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|SIMPLE_SEGMENT|2081,2094|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2081,2094|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|SIMPLE_SEGMENT|2081,2094|false|false|false|||pembrolizumab
Event|Event|SIMPLE_SEGMENT|2108,2116|false|false|false|||Consider
Event|Event|SIMPLE_SEGMENT|2117,2125|false|false|false|||starting
Drug|Organic Chemical|SIMPLE_SEGMENT|2126,2140|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2126,2140|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|SIMPLE_SEGMENT|2126,2140|false|false|false|||spironolactone
Finding|Idea or Concept|SIMPLE_SEGMENT|2149,2156|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2157,2162|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|2157,2162|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|2157,2162|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|2164,2173|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|2164,2173|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2164,2173|false|false|false|C0033095||pressures
Event|Event|SIMPLE_SEGMENT|2175,2182|false|false|false|||trialed
Drug|Organic Chemical|SIMPLE_SEGMENT|2183,2191|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2183,2191|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|2183,2191|false|false|false|||losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|2196,2210|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2196,2210|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|SIMPLE_SEGMENT|2196,2210|false|false|false|||spironolactone
Event|Event|SIMPLE_SEGMENT|2224,2233|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2224,2233|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|2250,2254|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|2262,2273|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|2262,2273|false|false|false|C0020649|Hypotension|hypotension
Event|Event|SIMPLE_SEGMENT|2283,2287|false|false|false|||LFTs
Event|Event|SIMPLE_SEGMENT|2298,2307|false|false|false|||rechecked
Event|Event|SIMPLE_SEGMENT|2323,2332|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|2323,2332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2323,2332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2323,2332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2323,2332|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|2350,2357|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2350,2360|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|2361,2374|false|false|false|||transaminitis
Finding|Finding|SIMPLE_SEGMENT|2361,2374|false|false|false|C2242708|Hypertransaminasaemia|transaminitis
Event|Event|SIMPLE_SEGMENT|2375,2385|false|false|false|||attributed
Finding|Idea or Concept|SIMPLE_SEGMENT|2389,2393|false|false|false|C1552020|Role Class - part|part
Drug|Organic Chemical|SIMPLE_SEGMENT|2398,2404|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2398,2404|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|SIMPLE_SEGMENT|2398,2404|false|false|false|C1414273|EEF1A2 gene|statin
Event|Event|SIMPLE_SEGMENT|2405,2408|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2405,2408|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2405,2408|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|SIMPLE_SEGMENT|2429,2438|false|false|false|||restarted
Drug|Organic Chemical|SIMPLE_SEGMENT|2442,2454|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2442,2454|false|false|false|C0965129|rosuvastatin|rosuvastatin
Event|Event|SIMPLE_SEGMENT|2442,2454|false|false|false|||rosuvastatin
Event|Event|SIMPLE_SEGMENT|2461,2470|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2461,2470|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|2478,2485|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2478,2485|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2478,2485|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2478,2485|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2478,2488|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2489,2492|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2489,2492|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2489,2492|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2489,2492|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2489,2492|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2489,2492|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2489,2492|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2489,2492|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|2497,2501|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2497,2501|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|2508,2512|false|false|false|||LFTs
Finding|Idea or Concept|SIMPLE_SEGMENT|2516,2519|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|2516,2519|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|2524,2533|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2524,2533|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2539,2542|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2539,2542|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|2539,2542|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|2539,2542|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|2539,2542|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|2539,2542|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|2539,2542|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2539,2542|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2547,2550|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2547,2550|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2547,2550|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2547,2550|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|2547,2550|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|2547,2550|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|2547,2550|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2555,2558|false|false|false|C1663627|ALK protein, human|Alk
Drug|Enzyme|SIMPLE_SEGMENT|2555,2558|false|false|false|C1663627|ALK protein, human|Alk
Finding|Gene or Genome|SIMPLE_SEGMENT|2555,2558|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|Alk
Finding|Receptor|SIMPLE_SEGMENT|2555,2558|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|Alk
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2555,2563|false|false|false|C0002059|Alkaline Phosphatase|Alk phos
Drug|Enzyme|SIMPLE_SEGMENT|2555,2563|false|false|false|C0002059|Alkaline Phosphatase|Alk phos
Event|Event|SIMPLE_SEGMENT|2555,2563|false|false|false|||Alk phos
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2555,2563|false|false|false|C0201850|Alkaline phosphatase measurement|Alk phos
Event|Event|SIMPLE_SEGMENT|2583,2589|false|false|false|||Follow
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2598,2606|false|false|false|C0027651|Neoplasms|Oncology
Event|Event|SIMPLE_SEGMENT|2598,2606|false|false|false|||Oncology
Procedure|Health Care Activity|SIMPLE_SEGMENT|2598,2606|false|false|false|C1555459|oncology services|Oncology
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2617,2625|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|SIMPLE_SEGMENT|2617,2625|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2617,2625|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|SIMPLE_SEGMENT|2617,2625|false|false|false|||melanoma
Event|Event|SIMPLE_SEGMENT|2630,2637|false|false|false|||Monitor
Event|Event|SIMPLE_SEGMENT|2642,2652|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|2642,2652|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|2642,2652|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Functional Concept|SIMPLE_SEGMENT|2656,2668|false|false|false|C2348609|Supplement|supplemental
Event|Event|SIMPLE_SEGMENT|2672,2683|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|2672,2683|false|false|false|C1514873|Requirement|requirement
Event|Event|SIMPLE_SEGMENT|2691,2700|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|2691,2700|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2691,2700|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2691,2700|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2691,2700|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|2709,2718|false|false|false|||requiring
Finding|Finding|SIMPLE_SEGMENT|2738,2742|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|2738,2742|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|2738,2742|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|2747,2756|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2747,2756|false|false|false|C0030685|Patient Discharge|discharge
Finding|Mental Process|SIMPLE_SEGMENT|2765,2772|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|2776,2786|false|false|false|||recovering
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2792,2801|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|2792,2801|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|2804,2813|false|false|false|||DISCHARGE
Finding|Body Substance|SIMPLE_SEGMENT|2804,2813|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2804,2813|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2804,2813|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2804,2813|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2825,2828|false|false|false|||lbs
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2825,2828|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Body Substance|SIMPLE_SEGMENT|2847,2856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2847,2856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2847,2856|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2847,2856|false|false|false|C0030685|Patient Discharge|DISCHARGE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2857,2865|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|DIURETIC
Event|Event|SIMPLE_SEGMENT|2857,2865|false|false|false|||DIURETIC
Drug|Organic Chemical|SIMPLE_SEGMENT|2867,2876|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2867,2876|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|2867,2876|false|false|false|||torsemide
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2886,2889|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2886,2889|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2886,2889|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|2886,2889|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|2886,2889|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|2891,2898|false|false|false|||SUMMARY
Finding|Intellectual Product|SIMPLE_SEGMENT|2891,2898|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Event|Event|SIMPLE_SEGMENT|2942,2945|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|2942,2945|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2966,2969|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2966,2969|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2966,2969|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2966,2969|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2966,2969|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2966,2969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2966,2969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2966,2969|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|2977,2981|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2977,2981|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3003,3006|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3003,3006|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|3003,3006|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|3003,3006|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|3003,3006|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3003,3006|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3014,3017|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3014,3017|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3014,3017|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3014,3017|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|3025,3033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|3025,3033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|SIMPLE_SEGMENT|3025,3057|false|false|false|C3276922|Tricuspid regurgitation, moderate|moderate tricuspid regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3034,3057|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|SIMPLE_SEGMENT|3044,3057|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|3044,3057|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3044,3057|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3044,3057|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Functional Concept|SIMPLE_SEGMENT|3059,3064|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Pathologic Function|SIMPLE_SEGMENT|3059,3088|false|false|false|C0242707|Right Ventricular Dysfunction|right ventricular dysfunction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3065,3076|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|SIMPLE_SEGMENT|3065,3088|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3077,3088|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|3077,3088|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|3077,3088|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|3077,3088|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|3077,3088|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|SIMPLE_SEGMENT|3090,3098|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|3090,3098|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Pathologic Function|SIMPLE_SEGMENT|3090,3121|false|false|false|C5395246|Moderate pulmonary hypertension|moderate pulmonary hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3099,3108|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3099,3108|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3099,3108|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|3099,3121|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3109,3121|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|3109,3121|false|false|false|||hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3138,3144|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3146,3158|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|3146,3158|false|false|false|||fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|3162,3170|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3162,3170|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|3162,3170|false|false|false|||apixaban
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3172,3177|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|3182,3189|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|3182,3189|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3182,3204|false|false|false|C1561643|Chronic Kidney Diseases|chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3190,3196|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3190,3196|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|3190,3196|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3190,3196|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3190,3196|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3190,3204|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3197,3204|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|3197,3204|false|false|false|||disease
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3207,3215|false|false|false|C0168634|BaseLine dental cement|Baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|3207,3215|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3229,3252|false|false|false|C0007820|Cerebrovascular Disorders|cerebrovascular disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3245,3252|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|3245,3252|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|3258,3268|false|false|false|||metastatic
Finding|Functional Concept|SIMPLE_SEGMENT|3258,3268|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3270,3278|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|SIMPLE_SEGMENT|3270,3278|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3270,3278|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|SIMPLE_SEGMENT|3270,3278|false|false|false|||melanoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3270,3297|false|false|false|C4745280|Melanoma of Unknown Primary|melanoma of unknown primary
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3282,3289|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|3282,3289|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3282,3289|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|3282,3289|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|3282,3289|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|3282,3289|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|3282,3289|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|3282,3289|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3301,3314|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Immunologic Factor|SIMPLE_SEGMENT|3301,3314|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3301,3314|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Finding|Functional Concept|SIMPLE_SEGMENT|3316,3323|false|false|false|C4520523|On hold|on hold
Event|Activity|SIMPLE_SEGMENT|3319,3323|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|SIMPLE_SEGMENT|3319,3323|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|SIMPLE_SEGMENT|3319,3323|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Event|Event|SIMPLE_SEGMENT|3324,3329|false|false|false|||since
Event|Event|SIMPLE_SEGMENT|3349,3362|false|false|false|||transaminitis
Finding|Finding|SIMPLE_SEGMENT|3349,3362|false|false|false|C2242708|Hypertransaminasaemia|transaminitis
Event|Event|SIMPLE_SEGMENT|3367,3374|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|3367,3374|false|false|false|C2699424|Concern|concern
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3380,3394|false|false|false|C0876994|Cardiotoxicity|cardiotoxicity
Event|Event|SIMPLE_SEGMENT|3380,3394|false|false|false|||cardiotoxicity
Event|Event|SIMPLE_SEGMENT|3404,3412|false|false|false|||admitted
Finding|Intellectual Product|SIMPLE_SEGMENT|3418,3424|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|3418,3433|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|3425,3433|false|false|false|||overload
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3439,3444|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3439,3444|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3439,3444|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Functional Concept|SIMPLE_SEGMENT|3446,3453|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|3446,3453|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|3446,3453|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|3454,3466|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|3454,3466|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3471,3480|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|3471,3480|false|false|false|||pneumonia
Finding|Finding|SIMPLE_SEGMENT|3486,3490|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|3486,3490|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|3486,3490|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3491,3497|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3491,3497|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3491,3497|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|3491,3497|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3491,3497|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|3499,3511|false|false|false|||requirements
Event|Event|SIMPLE_SEGMENT|3539,3548|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3539,3548|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|3553,3557|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|3553,3557|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|3553,3557|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|3558,3562|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3558,3562|false|false|false|C0806140|Flow|flow
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3564,3570|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3564,3570|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3564,3570|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|3564,3570|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3564,3570|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|3572,3578|false|false|false|||weaned
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3582,3587|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3582,3587|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|3582,3587|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3582,3587|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|3582,3587|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|3582,3587|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3588,3595|false|false|false|C1550232|Body Parts - Cannula|cannula
Event|Event|SIMPLE_SEGMENT|3588,3595|false|false|false|||cannula
Finding|Body Substance|SIMPLE_SEGMENT|3588,3595|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|3588,3595|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Individual Behavior|SIMPLE_SEGMENT|3602,3612|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|3602,3612|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Event|Event|SIMPLE_SEGMENT|3616,3624|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3616,3624|false|false|false|C0012797|Diuresis|diuresis
Event|Event|SIMPLE_SEGMENT|3630,3639|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|3630,3639|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|3630,3639|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|3630,3639|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3630,3639|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3643,3652|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|3643,3652|false|false|false|||pneumonia
Finding|Idea or Concept|SIMPLE_SEGMENT|3660,3663|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|3660,3663|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|3664,3670|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|3674,3679|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|3674,3679|false|false|false|C0250482|Zosyn|Zosyn
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3697,3707|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|3697,3707|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|3697,3707|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3697,3707|false|false|false|C0489941|Vancomycin measurement|vancomycin
Event|Event|SIMPLE_SEGMENT|3723,3734|false|false|false|||transferred
Anatomy|Body System|SIMPLE_SEGMENT|3738,3748|false|false|false|C0007226|Cardiovascular system|cardiology
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3750,3755|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|3765,3774|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|3778,3785|false|false|false|||diurese
Finding|Finding|SIMPLE_SEGMENT|3786,3790|false|false|false|C5575035|Well (answer to question)|well
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3799,3805|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3799,3805|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3799,3805|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|3799,3805|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3799,3805|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|3807,3818|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|3807,3818|false|false|false|C1514873|Requirement|requirement
Event|Event|SIMPLE_SEGMENT|3823,3829|false|false|false|||weaned
Event|Event|SIMPLE_SEGMENT|3845,3857|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|3868,3877|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3868,3877|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|3868,3877|false|false|false|||torsemide
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3881,3884|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3881,3884|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3881,3884|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|3881,3884|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|3881,3884|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|3902,3912|false|false|false|||maintained
Event|Event|SIMPLE_SEGMENT|3913,3922|false|false|false|||euvolemia
Finding|Finding|SIMPLE_SEGMENT|3913,3922|false|false|false|C1845208|Euvolemia|euvolemia
Finding|Intellectual Product|SIMPLE_SEGMENT|3926,3931|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|3932,3938|false|false|false|||ISSUES
Finding|Intellectual Product|SIMPLE_SEGMENT|3958,3963|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3958,3997|false|false|false|C2733492|Acute on chronic systolic heart failure|Acute on chronic systolic heart failure
Finding|Intellectual Product|SIMPLE_SEGMENT|3967,3974|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|3967,3974|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3967,3997|false|false|false|C1135194|Chronic systolic heart failure|chronic systolic heart failure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3975,3983|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3975,3997|false|false|false|C1135191|Heart Failure, Systolic|systolic heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3984,3989|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3984,3989|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3984,3989|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3984,3997|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|3990,3997|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|3990,3997|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|3990,3997|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|3990,3997|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|3998,4010|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|3998,4010|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Body Substance|SIMPLE_SEGMENT|4011,4018|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4011,4018|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4011,4018|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|4024,4031|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4024,4031|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4024,4031|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4024,4031|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4024,4034|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|4024,4048|false|false|false|C0455531||history of heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4035,4040|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4035,4040|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4035,4040|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4035,4048|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|4041,4048|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|4041,4048|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|4041,4048|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|4041,4048|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|4054,4062|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|4054,4062|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|4054,4062|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Finding|SIMPLE_SEGMENT|4063,4069|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4063,4069|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Functional Concept|SIMPLE_SEGMENT|4071,4079|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4071,4094|false|false|false|C0349782|Ischemic cardiomyopathy|ischemic cardiomyopathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4080,4094|false|false|false|C0878544|Cardiomyopathies|cardiomyopathy
Event|Event|SIMPLE_SEGMENT|4080,4094|false|false|false|||cardiomyopathy
Event|Event|SIMPLE_SEGMENT|4101,4108|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4101,4108|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4101,4108|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4101,4108|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4101,4111|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4112,4115|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4112,4115|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|4112,4115|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|4112,4115|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|4112,4115|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4112,4115|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|4112,4115|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4112,4115|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|4120,4124|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4120,4124|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4129,4132|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4129,4132|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|4129,4132|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|4129,4132|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|4129,4132|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4129,4132|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Event|SIMPLE_SEGMENT|4135,4143|false|false|false|||Admitted
Drug|Substance|SIMPLE_SEGMENT|4149,4154|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4149,4154|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4149,4154|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|SIMPLE_SEGMENT|4149,4163|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Finding|Pathologic Function|SIMPLE_SEGMENT|4149,4163|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Event|Event|SIMPLE_SEGMENT|4155,4163|false|false|false|||overload
Anatomy|Tissue|SIMPLE_SEGMENT|4168,4175|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4168,4175|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|4168,4184|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|4168,4184|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4168,4184|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|4176,4184|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|4176,4184|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|4176,4184|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4176,4184|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4186,4193|false|false|false|C0032930|Precipitating Factors|Trigger
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4199,4206|false|false|false|C1705970|Electrical Current|current
Event|Event|SIMPLE_SEGMENT|4207,4219|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|4207,4219|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4229,4239|false|false|false|C0009450|Communicable Diseases|infectious
Event|Event|SIMPLE_SEGMENT|4229,4239|false|false|false|||infectious
Event|Event|SIMPLE_SEGMENT|4246,4254|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4246,4254|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4246,4257|false|true|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4259,4268|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|4259,4268|false|false|false|||pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|4272,4276|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4272,4287|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4277,4282|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4277,4282|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4277,4287|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4283,4287|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4283,4287|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|4291,4300|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4291,4300|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|4302,4309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4302,4309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4302,4309|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|4315,4319|false|false|false|||high
Finding|Finding|SIMPLE_SEGMENT|4315,4319|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|4315,4319|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|4315,4319|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4321,4327|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4321,4327|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4321,4327|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4321,4327|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|4328,4340|false|false|false|||requirements
Event|Event|SIMPLE_SEGMENT|4350,4359|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4350,4359|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|4364,4373|false|false|false|||responded
Event|Event|SIMPLE_SEGMENT|4392,4400|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4392,4400|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|SIMPLE_SEGMENT|4406,4411|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4406,4411|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|4422,4430|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4422,4430|false|false|false|C0012797|Diuresis|diuresis
Finding|Body Substance|SIMPLE_SEGMENT|4432,4439|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4432,4439|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4432,4439|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|4445,4457|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|4461,4470|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4461,4470|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|4461,4470|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|4475,4485|false|false|false|||maintained
Event|Event|SIMPLE_SEGMENT|4489,4498|false|false|false|||euvolemia
Finding|Finding|SIMPLE_SEGMENT|4489,4498|false|false|false|C1845208|Euvolemia|euvolemia
Event|Event|SIMPLE_SEGMENT|4516,4524|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4516,4524|false|false|false|C0012797|Diuresis|diuresis
Finding|Body Substance|SIMPLE_SEGMENT|4530,4537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4530,4537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4530,4537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4540,4546|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4540,4546|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4540,4546|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4540,4546|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|4547,4558|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|4547,4558|false|false|false|C1514873|Requirement|requirement
Event|Event|SIMPLE_SEGMENT|4570,4577|false|false|false|||lowered
Event|Event|SIMPLE_SEGMENT|4607,4617|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|4621,4630|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4621,4630|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|4621,4630|false|false|false|||torsemide
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4641,4644|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4641,4644|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4641,4644|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|4641,4644|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4641,4644|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|4653,4659|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|4653,4659|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|4663,4671|false|false|false|||tolerate
Event|Event|SIMPLE_SEGMENT|4691,4697|false|false|false|||agents
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4716,4724|false|false|false|C3540676|Blockade|blockade
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4716,4724|false|false|false|C3540676|Blockade|blockade
Event|Event|SIMPLE_SEGMENT|4716,4724|false|false|false|||blockade
Finding|Functional Concept|SIMPLE_SEGMENT|4716,4724|false|false|false|C0332206|Blocking|blockade
Event|Event|SIMPLE_SEGMENT|4725,4731|false|false|false|||agents
Event|Event|SIMPLE_SEGMENT|4739,4750|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|4739,4750|false|false|false|C0020649|Hypotension|hypotension
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4756,4761|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|SIMPLE_SEGMENT|4756,4761|false|false|false|C2003888|Lower (action)|Lower
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4756,4781|false|false|false|C0585104|Left lower zone pneumonia|Lower left lobe pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|4762,4766|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4767,4771|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4767,4771|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4772,4781|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|4772,4781|false|false|false|||pneumonia
Finding|Body Substance|SIMPLE_SEGMENT|4782,4789|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4782,4789|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4782,4789|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|4795,4803|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4795,4803|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4795,4806|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4807,4816|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|4807,4816|false|false|false|||pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|4824,4828|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4824,4839|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4829,4834|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4829,4834|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4829,4839|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4835,4839|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4835,4839|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Drug|Antibiotic|SIMPLE_SEGMENT|4856,4861|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|4856,4861|false|false|false|C0250482|Zosyn|zosyn
Event|Event|SIMPLE_SEGMENT|4856,4861|false|false|false|||zosyn
Event|Event|SIMPLE_SEGMENT|4873,4881|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|4873,4881|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|4886,4895|false|false|false|||continued
Drug|Antibiotic|SIMPLE_SEGMENT|4899,4904|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|4899,4904|false|false|false|C0250482|Zosyn|Zosyn
Finding|Idea or Concept|SIMPLE_SEGMENT|4928,4931|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|4928,4931|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|4944,4954|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|4944,4954|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|4944,4954|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Event|Event|SIMPLE_SEGMENT|4958,4966|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|4958,4966|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4958,4966|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|4972,4979|false|false|false|||suspect
Event|Event|SIMPLE_SEGMENT|5002,5013|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|5002,5013|false|false|false|C1514873|Requirement|requirement
Finding|Idea or Concept|SIMPLE_SEGMENT|5029,5033|false|false|false|C1552020|Role Class - part|part
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5059,5072|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|5059,5072|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|5073,5077|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|5073,5077|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5093,5102|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5093,5102|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5093,5102|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|5111,5120|false|false|false|||requiring
Finding|Functional Concept|SIMPLE_SEGMENT|5128,5140|false|false|false|C2348609|Supplement|supplemental
Finding|Finding|SIMPLE_SEGMENT|5154,5158|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|5154,5158|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|5154,5158|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|5162,5171|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|5162,5171|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5162,5171|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5162,5171|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5162,5171|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Tissue|SIMPLE_SEGMENT|5176,5183|false|false|false|C0032225|Pleura|Pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5176,5183|false|false|false|C0032226|Pleural Diseases|Pleural
Finding|Body Substance|SIMPLE_SEGMENT|5176,5192|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5176,5192|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5176,5192|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Event|Event|SIMPLE_SEGMENT|5184,5192|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5184,5192|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5184,5192|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5184,5192|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Body Substance|SIMPLE_SEGMENT|5204,5211|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5204,5211|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5204,5211|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|5217,5225|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5217,5225|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5217,5228|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|5229,5234|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|SIMPLE_SEGMENT|5235,5242|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5235,5242|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|5235,5251|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5235,5251|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5235,5251|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|5243,5251|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5243,5251|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5243,5251|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5243,5251|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Conceptual Entity|SIMPLE_SEGMENT|5253,5261|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|SIMPLE_SEGMENT|5253,5261|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Finding|SIMPLE_SEGMENT|5262,5268|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5262,5268|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Substance|SIMPLE_SEGMENT|5270,5275|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5270,5275|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|SIMPLE_SEGMENT|5270,5284|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Finding|Pathologic Function|SIMPLE_SEGMENT|5270,5284|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Event|Event|SIMPLE_SEGMENT|5276,5284|false|false|false|||overload
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5291,5296|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5291,5296|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5291,5296|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5291,5304|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|5297,5304|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|5297,5304|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|5297,5304|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|5297,5304|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5318,5326|false|false|false|C0812388|Ejection time|ejection
Event|Event|SIMPLE_SEGMENT|5318,5326|false|false|false|||ejection
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5318,5326|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5318,5326|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Event|Event|SIMPLE_SEGMENT|5328,5336|false|false|false|||fraction
Finding|Intellectual Product|SIMPLE_SEGMENT|5328,5336|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Anatomy|Tissue|SIMPLE_SEGMENT|5338,5345|false|false|false|C0032225|Pleura|Pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5338,5345|false|false|false|C0032226|Pleural Diseases|Pleural
Finding|Body Substance|SIMPLE_SEGMENT|5338,5354|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5338,5354|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5338,5354|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|Pleural effusion
Event|Event|SIMPLE_SEGMENT|5346,5354|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5346,5354|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5346,5354|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5346,5354|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5355,5363|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|5364,5372|false|false|false|||improved
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5378,5386|false|false|false|C0012797|Diuresis|diuresis
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5396,5402|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5396,5402|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5396,5402|false|false|false|C0030054|oxygen|oxygen
Event|Event|SIMPLE_SEGMENT|5396,5402|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5396,5402|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|5403,5414|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|5403,5414|false|false|false|C1514873|Requirement|requirement
Event|Event|SIMPLE_SEGMENT|5415,5422|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|5452,5465|false|false|false|||thoracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5452,5465|false|false|false|C0189477|Thoracentesis|thoracentesis
Event|Event|SIMPLE_SEGMENT|5470,5478|false|false|false|||deferred
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5484,5490|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5484,5503|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5484,5503|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5484,5503|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5491,5503|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|5491,5503|false|false|false|||fibrillation
Finding|Body Substance|SIMPLE_SEGMENT|5504,5511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5504,5511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5504,5511|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5517,5524|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5517,5524|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|SIMPLE_SEGMENT|5525,5532|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5525,5532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5525,5532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5525,5532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5525,5535|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|5525,5555|false|false|false|C0729790||history of atrial fibrillation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5536,5542|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5536,5555|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5536,5555|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5536,5555|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5543,5555|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|5543,5555|false|false|false|||fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5560,5564|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5560,5564|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|5582,5591|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5582,5591|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|5593,5602|false|false|false|||Continued
Drug|Organic Chemical|SIMPLE_SEGMENT|5603,5613|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5603,5613|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|5603,5613|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5603,5613|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|5618,5626|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5618,5626|false|false|false|C1831808|apixaban|apixaban
Event|Event|SIMPLE_SEGMENT|5618,5626|false|false|false|||apixaban
Event|Event|SIMPLE_SEGMENT|5649,5659|false|false|false|||controlled
Finding|Intellectual Product|SIMPLE_SEGMENT|5662,5669|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|5662,5669|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5696,5704|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5696,5711|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5696,5719|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5705,5711|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5705,5711|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5705,5719|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5712,5719|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|5712,5719|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|5724,5728|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5724,5728|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Body Substance|SIMPLE_SEGMENT|5729,5736|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5729,5736|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5729,5736|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|5742,5749|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5742,5749|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5742,5749|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5742,5749|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5742,5752|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5755,5761|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5755,5761|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|SIMPLE_SEGMENT|5762,5766|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5762,5766|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5795,5798|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5795,5798|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|5795,5798|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|5795,5798|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|5795,5798|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5795,5798|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5802,5805|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5802,5805|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5802,5805|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|5813,5822|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|5823,5827|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5823,5827|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5823,5827|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|5828,5835|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5828,5835|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|5828,5835|false|false|false|||aspirin
Finding|Body Substance|SIMPLE_SEGMENT|5837,5844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5837,5844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5837,5844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|5850,5857|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|5861,5864|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5861,5864|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Organic Chemical|SIMPLE_SEGMENT|5870,5882|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5870,5882|false|false|false|C0965129|rosuvastatin|rosuvastatin
Event|Event|SIMPLE_SEGMENT|5870,5882|false|false|false|||rosuvastatin
Event|Event|SIMPLE_SEGMENT|5898,5904|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|5898,5904|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|5898,5904|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5938,5948|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|5938,5948|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5938,5948|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|5957,5961|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|5986,5998|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|6006,6018|false|false|false|||transamnitis
Finding|Finding|SIMPLE_SEGMENT|6037,6041|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|6037,6041|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|6037,6041|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|6049,6056|false|false|false|||unclear
Event|Event|SIMPLE_SEGMENT|6077,6083|false|false|false|||effect
Drug|Organic Chemical|SIMPLE_SEGMENT|6091,6097|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6091,6097|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|SIMPLE_SEGMENT|6091,6097|false|false|false|||statin
Finding|Gene or Genome|SIMPLE_SEGMENT|6091,6097|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6102,6115|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|SIMPLE_SEGMENT|6102,6115|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6102,6115|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|SIMPLE_SEGMENT|6102,6115|false|false|false|||pembrolizumab
Finding|Body Substance|SIMPLE_SEGMENT|6132,6139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6132,6139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6132,6139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|6132,6143|true|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|6156,6166|false|false|false|||checkpoint
Finding|Cell Function|SIMPLE_SEGMENT|6156,6166|true|false|false|C1155874|Cell Cycle Checkpoints|checkpoint
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6168,6177|false|false|false|C1999216|Inhibitor|inhibitor
Event|Event|SIMPLE_SEGMENT|6178,6185|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|6178,6185|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|6178,6185|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6178,6185|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|6201,6209|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|6201,6209|false|false|false|C0679006|Decision|decision
Drug|Organic Chemical|SIMPLE_SEGMENT|6226,6238|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6226,6238|false|false|false|C0965129|rosuvastatin|rosuvastatin
Event|Event|SIMPLE_SEGMENT|6226,6238|false|false|false|||rosuvastatin
Event|Event|SIMPLE_SEGMENT|6244,6251|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|6244,6251|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6244,6251|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6244,6266|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6252,6258|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6252,6258|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6252,6258|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6252,6258|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6252,6258|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6252,6266|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6259,6266|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6259,6266|false|false|false|||disease
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6267,6275|false|false|false|C0168634|BaseLine dental cement|Baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6267,6275|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6311,6315|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|6311,6315|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|6320,6328|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|6357,6366|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6357,6366|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6372,6378|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|6372,6378|false|false|false|||Anemia
Event|Event|SIMPLE_SEGMENT|6379,6386|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|6379,6386|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6379,6386|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Event|Event|SIMPLE_SEGMENT|6397,6406|false|false|false|||worsening
Event|Event|SIMPLE_SEGMENT|6421,6430|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6421,6430|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6432,6442|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6432,6442|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|6432,6442|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6432,6442|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|SIMPLE_SEGMENT|6432,6442|false|false|false|||hemoglobin
Finding|Finding|SIMPLE_SEGMENT|6432,6442|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6432,6442|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|SIMPLE_SEGMENT|6452,6460|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|6461,6467|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6461,6467|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6473,6489|false|false|false|C0040034|Thrombocytopenia|Thrombocytopenia
Event|Event|SIMPLE_SEGMENT|6473,6489|false|false|false|||Thrombocytopenia
Finding|Finding|SIMPLE_SEGMENT|6473,6489|false|false|false|C0392386|Decreased platelet count|Thrombocytopenia
Finding|Finding|SIMPLE_SEGMENT|6490,6499|false|false|false|C0087130|Uncertainty|Uncertain
Event|Event|SIMPLE_SEGMENT|6500,6508|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|6500,6508|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|6500,6508|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Event|Event|SIMPLE_SEGMENT|6527,6534|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|6527,6534|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6527,6534|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|SIMPLE_SEGMENT|6539,6548|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6539,6548|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Cell|SIMPLE_SEGMENT|6549,6558|false|false|false|C0005821|Blood Platelets|platelets
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6549,6558|false|false|false|C0443116|Platelets Product|platelets
Event|Event|SIMPLE_SEGMENT|6549,6558|false|false|false|||platelets
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6549,6558|false|false|false|C0032181|Platelet count (procedure)|platelets
Event|Event|SIMPLE_SEGMENT|6568,6575|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|6588,6595|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|6588,6595|true|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|6600,6608|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|6600,6608|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|6621,6630|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6621,6630|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6636,6644|false|false|false|C0025202|melanoma|Melanoma
Drug|Immunologic Factor|SIMPLE_SEGMENT|6636,6644|false|false|false|C0796561|Melanoma vaccine|Melanoma
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6636,6644|false|false|false|C0796561|Melanoma vaccine|Melanoma
Event|Event|SIMPLE_SEGMENT|6636,6644|false|false|false|||Melanoma
Finding|Body Substance|SIMPLE_SEGMENT|6645,6652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6645,6652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6645,6652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6658,6665|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6658,6665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6658,6665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6658,6665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6658,6668|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|SIMPLE_SEGMENT|6669,6679|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6669,6688|false|false|false|C0278883|Metastatic melanoma|metastatic melanoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6680,6688|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|SIMPLE_SEGMENT|6680,6688|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6680,6688|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|SIMPLE_SEGMENT|6680,6688|false|false|false|||melanoma
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6694,6701|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|6694,6701|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6694,6701|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|6694,6701|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|6694,6701|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|6694,6701|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|6694,6701|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|6694,6701|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|6715,6724|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|6715,6724|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|6715,6724|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|6715,6724|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6715,6724|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6730,6743|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|SIMPLE_SEGMENT|6730,6743|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6730,6743|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|SIMPLE_SEGMENT|6730,6743|false|false|false|||pembrolizumab
Event|Event|SIMPLE_SEGMENT|6749,6753|false|false|false|||held
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6768,6776|false|false|false|C0600688|Toxic effect|toxicity
Event|Event|SIMPLE_SEGMENT|6768,6776|false|false|false|||toxicity
Event|Event|SIMPLE_SEGMENT|6780,6784|false|false|false|||CODE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6786,6789|false|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|6786,6789|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|6786,6789|false|false|false|C0011015|daunorubicin|DNR
Event|Event|SIMPLE_SEGMENT|6786,6789|false|false|false|||DNR
Finding|Finding|SIMPLE_SEGMENT|6786,6789|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|6786,6789|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Activity|SIMPLE_SEGMENT|6794,6801|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|6794,6801|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|6794,6801|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|6794,6801|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|6794,6801|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6794,6801|false|false|false|C0392367|Physical contact|CONTACT
Event|Event|SIMPLE_SEGMENT|6813,6825|false|false|false|||Relationship
Finding|Idea or Concept|SIMPLE_SEGMENT|6813,6825|false|false|false|C1705630;C1706279|Concept Relationship;Object Relationship|Relationship
Finding|Gene or Genome|SIMPLE_SEGMENT|6827,6830|false|false|false|C1420310|SON gene|Son
Finding|Idea or Concept|SIMPLE_SEGMENT|6832,6837|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|Phone
Finding|Intellectual Product|SIMPLE_SEGMENT|6832,6837|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|Phone
Finding|Intellectual Product|SIMPLE_SEGMENT|6832,6844|false|false|false|C1515258|Telephone Number|Phone number
Event|Event|SIMPLE_SEGMENT|6838,6844|false|false|false|||number
Finding|Idea or Concept|SIMPLE_SEGMENT|6838,6844|false|false|false|C1554106|MDF AttributeType - Number|number
Procedure|Health Care Activity|SIMPLE_SEGMENT|6859,6868|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6887,6897|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6887,6897|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6887,6902|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|6898,6902|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|6898,6902|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|6906,6914|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|6919,6927|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6919,6927|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6919,6927|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|6919,6927|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|6919,6927|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6919,6927|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|6932,6942|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6932,6942|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|6932,6942|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6932,6942|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|6963,6971|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6963,6971|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6982,6985|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6982,6985|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6982,6985|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6982,6985|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6982,6985|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6990,6997|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6990,6997|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|7017,7025|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7017,7025|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|7017,7025|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|7017,7032|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7017,7032|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7026,7032|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7026,7032|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7026,7032|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7026,7032|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7026,7032|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7026,7032|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7043,7046|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7043,7046|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7043,7046|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7043,7046|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7043,7046|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7051,7058|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7051,7066|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7051,7066|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7059,7066|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7059,7066|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7059,7066|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|7059,7066|false|false|false|||Sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|7087,7092|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7087,7092|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|SIMPLE_SEGMENT|7111,7121|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7111,7121|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|7141,7151|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7141,7151|false|false|false|C0257343|tamsulosin|Tamsulosin
Event|Event|SIMPLE_SEGMENT|7162,7165|false|false|false|||QHS
Drug|Organic Chemical|SIMPLE_SEGMENT|7170,7179|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7170,7179|false|false|false|C0076840|torsemide|Torsemide
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7200,7208|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|SIMPLE_SEGMENT|7200,7208|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|SIMPLE_SEGMENT|7200,7208|false|false|false|||coenzyme
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7200,7212|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|SIMPLE_SEGMENT|7200,7212|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7200,7212|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|SIMPLE_SEGMENT|7209,7212|false|false|false|||Q10
Finding|Gene or Genome|SIMPLE_SEGMENT|7209,7212|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7220,7224|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7220,7224|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|7220,7224|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|7220,7224|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|7225,7230|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|7236,7241|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7236,7241|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7243,7267|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|SIMPLE_SEGMENT|7259,7267|false|false|false|||infantis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7274,7278|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7274,7278|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|7274,7278|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|7274,7278|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|7279,7284|false|false|false|||DAILY
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7290,7299|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7290,7299|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|7290,7299|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7290,7299|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7290,7299|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|7290,7299|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|7290,7299|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7290,7299|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7290,7308|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7290,7308|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7300,7308|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|SIMPLE_SEGMENT|7300,7308|false|false|false|||Chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|7300,7308|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7300,7308|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|SIMPLE_SEGMENT|7312,7315|false|false|false|||mEq
Event|Event|SIMPLE_SEGMENT|7329,7338|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7329,7338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7329,7338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7329,7338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7329,7338|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7329,7350|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7339,7350|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7339,7350|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7339,7350|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7339,7350|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|7356,7368|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7356,7368|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Event|Event|SIMPLE_SEGMENT|7356,7368|false|false|false|||Rosuvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|7356,7376|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7356,7376|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7369,7376|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7369,7376|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7369,7376|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7369,7376|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|7369,7376|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|7369,7376|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|7369,7376|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7369,7376|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|7385,7388|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|7395,7402|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7395,7402|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|7395,7402|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|7395,7404|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|7395,7404|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7395,7404|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|7395,7404|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7395,7404|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|7403,7404|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|7410,7414|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|7430,7439|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7430,7439|false|false|false|C0076840|torsemide|Torsemide
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7449,7452|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7449,7452|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7449,7452|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7449,7452|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7449,7452|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|7459,7464|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7459,7464|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7466,7490|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|SIMPLE_SEGMENT|7482,7490|false|false|false|||infantis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7497,7501|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7497,7501|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|7497,7501|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|7497,7501|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|7502,7507|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|7514,7524|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7514,7524|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|7514,7524|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7514,7524|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|7547,7555|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7547,7555|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7566,7569|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7566,7569|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7566,7569|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7566,7569|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7566,7569|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|7576,7583|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7576,7583|false|false|false|C0004057|aspirin|Aspirin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7605,7613|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|SIMPLE_SEGMENT|7605,7613|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|SIMPLE_SEGMENT|7605,7613|false|false|false|||coenzyme
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7605,7617|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|SIMPLE_SEGMENT|7605,7617|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7605,7617|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|SIMPLE_SEGMENT|7614,7617|false|false|false|||Q10
Finding|Gene or Genome|SIMPLE_SEGMENT|7614,7617|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7625,7629|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7625,7629|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|7625,7629|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|7625,7629|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|7630,7635|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|7642,7650|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7642,7650|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|7642,7650|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|7642,7657|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7642,7657|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7651,7657|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7651,7657|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7651,7657|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7651,7657|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7651,7657|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7651,7657|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7668,7671|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7668,7671|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7668,7671|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7668,7671|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7668,7671|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7679,7686|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7679,7694|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7679,7694|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7687,7694|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7687,7694|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7687,7694|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|7687,7694|false|false|false|||Sulfate
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7718,7727|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7718,7727|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|7718,7727|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7718,7727|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7718,7727|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|7718,7727|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|7718,7727|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7718,7727|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7718,7736|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7718,7736|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7728,7736|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|SIMPLE_SEGMENT|7728,7736|false|false|false|||Chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|7728,7736|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7728,7736|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|SIMPLE_SEGMENT|7740,7743|false|false|false|||mEq
Drug|Organic Chemical|SIMPLE_SEGMENT|7760,7765|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7760,7765|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|SIMPLE_SEGMENT|7787,7797|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7787,7797|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|7820,7830|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7820,7830|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Hormone|SIMPLE_SEGMENT|7856,7873|false|false|false|C0026160;C1641843|Mineralocorticoid (substance);Mineralocorticoids|mineralocorticoid
Drug|Organic Chemical|SIMPLE_SEGMENT|7856,7873|false|false|false|C0026160;C1641843|Mineralocorticoid (substance);Mineralocorticoids|mineralocorticoid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7856,7873|false|false|false|C0026160;C1641843|Mineralocorticoid (substance);Mineralocorticoids|mineralocorticoid
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7856,7882|false|false|false|C0066563;C3254418|Mineralocorticoid Receptor;NR3C2 protein, human|mineralocorticoid receptor
Finding|Gene or Genome|SIMPLE_SEGMENT|7856,7882|false|false|false|C0066563;C1417835;C3254418|Mineralocorticoid Receptor;NR3C2 gene;NR3C2 protein, human|mineralocorticoid receptor
Finding|Receptor|SIMPLE_SEGMENT|7856,7882|false|false|false|C0066563;C1417835;C3254418|Mineralocorticoid Receptor;NR3C2 gene;NR3C2 protein, human|mineralocorticoid receptor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7856,7893|false|false|false|C1579268;C5552626|Mineralocorticoid Receptor Antagonist [EPC];Mineralocorticoid Receptor Antagonists|mineralocorticoid receptor antagonist
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7874,7882|false|false|false|C0597357|receptor|receptor
Event|Event|SIMPLE_SEGMENT|7874,7882|false|false|false|||receptor
Finding|Receptor|SIMPLE_SEGMENT|7874,7882|false|false|false|C0597357|receptor|receptor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7874,7893|false|false|false|C4721408;C5399721|Receptor Antagonist [APC];Substance with receptor antagonist mechanism of action (substance)|receptor antagonist
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7883,7893|false|false|false|C4721408|Substance with receptor antagonist mechanism of action (substance)|antagonist
Event|Event|SIMPLE_SEGMENT|7883,7893|false|false|false|||antagonist
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7883,7893|false|false|false|C0231491|Antagonist muscle action|antagonist
Event|Event|SIMPLE_SEGMENT|7894,7898|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|7907,7914|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|7907,7914|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|7918,7929|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|7918,7929|false|false|false|C0020649|Hypotension|hypotension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7934,7937|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|7934,7937|false|false|false|||CKD
Finding|Body Substance|SIMPLE_SEGMENT|7939,7946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7939,7946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7939,7946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7950,7960|false|false|false|||intolerant
Finding|Functional Concept|SIMPLE_SEGMENT|7950,7960|false|false|false|C0231200|intolerant|intolerant
Event|Event|SIMPLE_SEGMENT|7964,7968|false|false|false|||beta
Finding|Intellectual Product|SIMPLE_SEGMENT|7964,7968|false|false|false|C0439096|Greek letter beta|beta
Event|Event|SIMPLE_SEGMENT|7970,7978|false|false|false|||blockers
Event|Event|SIMPLE_SEGMENT|7986,7995|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7986,7995|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|7996,8007|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|7996,8007|false|false|false|C0020649|Hypotension|hypotension
Event|Event|SIMPLE_SEGMENT|8022,8031|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8022,8031|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8022,8031|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8022,8031|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8022,8031|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8022,8043|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8022,8043|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8032,8043|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8032,8043|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8032,8043|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|8045,8053|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8045,8053|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|8045,8058|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|8054,8058|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|8054,8058|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|8054,8058|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|8054,8058|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|8061,8069|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|8061,8069|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|8077,8086|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8077,8086|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8077,8086|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8077,8086|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8077,8086|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8077,8096|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8087,8096|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8087,8096|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8087,8096|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8087,8096|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8087,8096|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8098,8115|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8106,8115|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|8106,8115|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|8106,8115|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8106,8115|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8106,8115|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|8139,8144|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8139,8178|false|false|false|C2733492|Acute on chronic systolic heart failure|Acute on chronic systolic heart failure
Finding|Intellectual Product|SIMPLE_SEGMENT|8148,8155|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|8148,8155|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8148,8178|false|false|false|C1135194|Chronic systolic heart failure|chronic systolic heart failure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8156,8164|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8156,8178|false|false|false|C1135191|Heart Failure, Systolic|systolic heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8165,8170|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8165,8170|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|8165,8170|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8165,8178|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|8171,8178|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|8171,8178|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|8171,8178|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|8171,8178|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|8179,8191|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|8179,8191|false|false|false|C4086268|Exacerbation|exacerbation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8192,8197|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|SIMPLE_SEGMENT|8192,8197|false|false|false|C2003888|Lower (action)|Lower
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8192,8217|false|false|false|C0585104|Left lower zone pneumonia|Lower left lobe pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|8198,8202|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8203,8207|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|8203,8207|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8208,8217|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|8208,8217|false|false|false|||pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8218,8244|false|false|false|C0747635|Bilateral pleural effusion|Bilateral pleural effusion
Anatomy|Tissue|SIMPLE_SEGMENT|8228,8235|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8228,8235|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|8228,8244|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|8228,8244|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|8228,8244|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|8236,8244|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|8236,8244|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|8236,8244|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|8236,8244|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8245,8251|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8245,8264|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8245,8264|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8245,8264|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8252,8264|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|8252,8264|false|false|false|||fibrillation
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8266,8275|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|8266,8275|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|8266,8275|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8266,8285|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|SIMPLE_SEGMENT|8266,8285|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8276,8285|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|8276,8285|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|8276,8285|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8276,8285|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8276,8285|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8309,8317|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8309,8324|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8309,8332|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8318,8324|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|8318,8324|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8318,8332|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8325,8332|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8325,8332|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8333,8339|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|8333,8339|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|8333,8339|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|8345,8349|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8345,8349|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|8350,8357|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|8350,8357|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|8350,8357|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8350,8372|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8358,8364|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8358,8364|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|8358,8364|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8358,8364|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8358,8364|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8358,8372|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8365,8372|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8365,8372|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8373,8379|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|8373,8379|false|false|false|||Anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8380,8396|false|false|false|C0040034|Thrombocytopenia|Thrombocytopenia
Event|Event|SIMPLE_SEGMENT|8380,8396|false|false|false|||Thrombocytopenia
Finding|Finding|SIMPLE_SEGMENT|8380,8396|false|false|false|C0392386|Decreased platelet count|Thrombocytopenia
Finding|Functional Concept|SIMPLE_SEGMENT|8397,8407|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8397,8416|false|false|false|C0278883|Metastatic melanoma|Metastatic melanoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8408,8416|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|SIMPLE_SEGMENT|8408,8416|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8408,8416|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|SIMPLE_SEGMENT|8408,8416|false|false|false|||melanoma
Event|Event|SIMPLE_SEGMENT|8420,8429|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8420,8429|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8420,8429|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8420,8429|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8420,8429|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8430,8439|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8430,8439|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|8430,8439|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8430,8439|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|8441,8447|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8441,8454|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8441,8454|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8448,8454|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8448,8454|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|8456,8461|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|8456,8461|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|8466,8474|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|8466,8474|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|8476,8481|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8476,8498|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8476,8498|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|8485,8498|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|8485,8498|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8485,8498|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8500,8505|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8500,8505|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8500,8505|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|8500,8505|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|8500,8505|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8500,8505|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8500,8505|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|8510,8521|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|8510,8521|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|8523,8531|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8523,8531|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8523,8531|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8532,8538|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|8532,8538|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8532,8538|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|8540,8550|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|8540,8550|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|8540,8550|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|8540,8550|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|8553,8561|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|8562,8572|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|8562,8572|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8576,8579|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|8576,8579|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|SIMPLE_SEGMENT|8576,8579|false|false|false|||aid
Finding|Gene or Genome|SIMPLE_SEGMENT|8576,8579|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8576,8579|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|SIMPLE_SEGMENT|8581,8587|false|false|false|||walker
Event|Event|SIMPLE_SEGMENT|8602,8611|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8602,8611|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8602,8611|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8602,8611|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8602,8611|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8602,8624|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8602,8624|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8602,8624|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8612,8624|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8612,8624|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8612,8624|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|8626,8630|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|8650,8658|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|8650,8658|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|8650,8658|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|8666,8670|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8666,8670|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8666,8670|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8666,8670|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8666,8673|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|8701,8704|false|false|false|||WAS
Event|Event|SIMPLE_SEGMENT|8714,8722|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|8714,8722|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|8767,8775|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|8796,8801|false|false|false|||short
Finding|Sign or Symptom|SIMPLE_SEGMENT|8796,8811|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|8805,8811|false|false|false|C0225386|Breath|breath
Event|Activity|SIMPLE_SEGMENT|8819,8827|false|false|false|C1709305|Occur (action)|HAPPENED
Event|Event|SIMPLE_SEGMENT|8819,8827|false|false|false|||HAPPENED
Finding|Idea or Concept|SIMPLE_SEGMENT|8835,8843|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|8891,8896|false|false|false|||found
Drug|Substance|SIMPLE_SEGMENT|8905,8910|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8905,8910|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8905,8910|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8919,8924|false|false|false|C0024109|Lung|lungs
Finding|Functional Concept|SIMPLE_SEGMENT|8955,8962|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|8955,8962|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|8955,8962|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|8955,8962|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|8955,8972|false|false|false|C4745084|Medical Condition|medical condition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8963,8972|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8963,8972|false|false|false|C0012634|Disease|condition
Event|Event|SIMPLE_SEGMENT|8963,8972|false|false|false|||condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8963,8972|false|false|false|C1705253|Logical Condition|condition
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8980,8985|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8980,8985|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|8980,8985|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8980,8993|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|8986,8993|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|8986,8993|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|8986,8993|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|8986,8993|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9007,9012|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9007,9012|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|9007,9012|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9007,9012|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|9022,9026|false|false|false|||pump
Event|Event|SIMPLE_SEGMENT|9032,9038|false|false|false|||enough
Drug|Substance|SIMPLE_SEGMENT|9043,9048|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9043,9048|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9043,9048|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9049,9054|false|false|false|C0004600||backs
Event|Event|SIMPLE_SEGMENT|9055,9057|false|false|false|||up
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9069,9074|false|false|false|C0024109|Lung|lungs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9096,9104|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9105,9115|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9105,9115|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9105,9115|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9119,9123|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|9124,9127|false|false|false|||get
Drug|Substance|SIMPLE_SEGMENT|9132,9137|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9132,9137|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9132,9137|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|9148,9156|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|9178,9183|false|false|false|||ready
Event|Event|SIMPLE_SEGMENT|9187,9192|false|false|false|||leave
Event|Event|SIMPLE_SEGMENT|9198,9206|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|9198,9206|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|9228,9232|false|false|false|||WHEN
Event|Event|SIMPLE_SEGMENT|9238,9242|false|false|false|||HOME
Finding|Idea or Concept|SIMPLE_SEGMENT|9238,9242|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|HOME
Finding|Intellectual Product|SIMPLE_SEGMENT|9238,9242|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|HOME
Procedure|Health Care Activity|SIMPLE_SEGMENT|9238,9242|false|false|false|C1553498|home health encounter|HOME
Event|Event|SIMPLE_SEGMENT|9283,9285|false|false|false|||Be
Event|Event|SIMPLE_SEGMENT|9286,9290|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|9286,9290|false|false|false|C4724437|SURE Test|sure
Event|Event|SIMPLE_SEGMENT|9294,9298|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9308,9319|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9308,9319|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9308,9319|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9308,9319|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9324,9330|false|false|false|||attend
Event|Activity|SIMPLE_SEGMENT|9344,9356|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|9344,9356|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|9357,9363|false|false|false|||listed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9379,9385|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|9379,9385|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|9379,9385|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|9379,9385|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|9379,9385|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|9389,9398|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9389,9398|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9389,9398|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9389,9398|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9389,9398|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9409,9412|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|SIMPLE_SEGMENT|9421,9426|false|false|false|||weigh
Finding|Finding|SIMPLE_SEGMENT|9443,9450|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|9446,9450|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|9446,9450|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|9446,9450|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9446,9450|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|9455,9458|false|false|false|||use
Finding|Finding|SIMPLE_SEGMENT|9472,9475|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|9472,9475|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9476,9484|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|9476,9484|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|9476,9484|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|9496,9501|false|false|false|||weigh
Finding|Idea or Concept|SIMPLE_SEGMENT|9517,9520|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9517,9520|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|9537,9541|false|false|false|||Call
Event|Event|SIMPLE_SEGMENT|9548,9554|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|9548,9554|false|false|false|C2348314|Doctor - Title|doctor
Drug|Organic Chemical|SIMPLE_SEGMENT|9562,9571|false|false|false|C1306677|Heartline|HeartLine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9562,9571|false|false|false|C1306677|Heartline|HeartLine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9587,9593|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|9587,9593|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|9587,9593|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|9587,9593|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|9587,9593|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|9594,9598|false|false|false|||goes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9618,9621|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Idea or Concept|SIMPLE_SEGMENT|9640,9651|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9652,9657|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9652,9657|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9652,9662|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9652,9662|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9658,9662|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9658,9662|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9658,9662|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9658,9662|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9668,9677|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9668,9687|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|9668,9687|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|9681,9687|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|9706,9714|false|false|false|||allowing
Event|Event|SIMPLE_SEGMENT|9724,9732|false|false|false|||involved
Event|Activity|SIMPLE_SEGMENT|9741,9745|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|9741,9745|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|9741,9745|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9741,9745|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9750,9754|false|false|false|C3273412|NCK-Interacting Protein with SH3 Domain|wish
Event|Event|SIMPLE_SEGMENT|9750,9754|false|false|false|||wish
Finding|Gene or Genome|SIMPLE_SEGMENT|9750,9754|false|false|false|C1423524;C3273411|NCKIPSD gene;NCKIPSD wt Allele|wish
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9768,9772|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|9768,9772|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|9768,9772|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|9806,9814|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9815,9827|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9815,9827|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9815,9827|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

