 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
MEDICINE|158,166
<EOL>|166,167
<EOL>|168,169
Sulfa|181,186
(|187,188
Sulfonamide|188,199
Antibiotics|200,211
)|211,212
/|213,214
Codeine|215,222
/|223,224
Bactrim|225,232
<EOL>|232,233
<EOL>|234,235
Attending|235,244
:|244,245
_|246,247
_|247,248
_|248,249
.|249,250
<EOL>|250,251
<EOL>|252,253
Shortness|270,279
of|280,282
breath|283,289
<EOL>|289,290
<EOL>|291,292
Major|292,297
Surgical|298,306
or|307,309
Invasive|310,318
Procedure|319,328
:|328,329
<EOL>|329,330
Percutaneous|330,342
liver|343,348
biopsy|349,355
<EOL>|355,356
<EOL>|357,358
Ms.|386,389
_|390,391
_|391,392
_|392,393
is|394,396
a|397,398
_|399,400
_|400,401
_|401,402
with|403,407
metastatic|408,418
cancer|419,425
of|426,428
unknown|429,436
primary|437,444
<EOL>|445,446
(|446,447
known|447,452
lesions|453,460
in|461,463
lungs|464,469
and|470,473
liver|474,479
)|479,480
presenting|481,491
with|492,496
shortness|497,506
of|507,509
<EOL>|510,511
breath|511,517
.|517,518
She|519,522
initially|523,532
presented|533,542
to|543,545
_|546,547
_|547,548
_|548,549
in|550,552
_|553,554
_|554,555
_|555,556
with|557,561
abdominal|562,571
<EOL>|572,573
pain|573,577
and|578,581
failure|582,589
to|590,592
thrive|593,599
.|599,600
Evaluation|601,611
at|612,614
that|615,619
time|620,624
included|625,633
an|634,636
<EOL>|637,638
abdominal|638,647
CT|648,650
scan|651,655
that|656,660
showed|661,667
multiple|668,676
lung|677,681
and|682,685
liver|686,691
<EOL>|692,693
metastases|693,703
.|703,704
She|705,708
has|709,712
yet|713,716
to|717,719
undergo|720,727
definite|728,736
diagnosis|737,746
with|747,751
<EOL>|752,753
biopsy|753,759
,|759,760
and|761,764
per|765,768
recent|769,775
oncology|776,784
documentation|785,798
seems|799,804
disengaged|805,815
<EOL>|816,817
with|817,821
care|822,826
.|826,827
<EOL>|829,830
She|830,833
was|834,837
reportedly|838,848
in|849,851
her|852,855
usual|856,861
state|862,867
of|868,870
health|871,877
until|878,883
the|884,887
<EOL>|888,889
evening|889,896
prior|897,902
to|903,905
admission|906,915
,|915,916
when|917,921
she|922,925
developed|926,935
acute|936,941
on|942,944
chronic|945,952
<EOL>|953,954
shortness|954,963
of|964,966
breath|967,973
while|974,979
at|980,982
rest|983,987
.|987,988
She|989,992
reported|993,1001
midsternal|1002,1012
chest|1013,1018
<EOL>|1019,1020
ache|1020,1024
associated|1025,1035
with|1036,1040
this|1041,1045
shortness|1046,1055
of|1056,1058
breath|1059,1065
.|1065,1066
Pain|1067,1071
is|1072,1074
<EOL>|1075,1076
exacerbated|1076,1087
by|1088,1090
direct|1091,1097
pressure|1098,1106
;|1106,1107
nothing|1108,1115
seems|1116,1121
to|1122,1124
alleviate|1125,1134
pain|1135,1139
.|1139,1140
<EOL>|1141,1142
She|1142,1145
denied|1146,1152
any|1153,1156
pleuritic|1157,1166
or|1167,1169
exertional|1170,1180
component|1181,1190
to|1191,1193
the|1194,1197
chest|1198,1203
<EOL>|1204,1205
pain|1205,1209
or|1210,1212
shortness|1213,1222
of|1223,1225
breath|1226,1232
.|1232,1233
She|1234,1237
feels|1238,1243
that|1244,1248
symptoms|1249,1257
are|1258,1261
<EOL>|1262,1263
secondary|1263,1272
to|1273,1275
her|1276,1279
"|1280,1281
cancer|1281,1287
"|1287,1288
and|1289,1292
"|1293,1294
feels|1294,1299
as|1300,1302
if|1303,1305
the|1306,1309
cancer|1310,1316
has|1317,1320
<EOL>|1321,1322
spread|1322,1328
"|1328,1329
.|1329,1330
She|1331,1334
reports|1335,1342
stable|1343,1349
,|1349,1350
chronic|1351,1358
nonproductive|1359,1372
cough|1373,1378
,|1378,1379
which|1380,1385
<EOL>|1386,1387
has|1387,1390
been|1391,1395
present|1396,1403
over|1404,1408
the|1409,1412
preceding|1413,1422
months|1423,1429
.|1429,1430
<EOL>|1432,1433
She|1433,1436
was|1437,1440
seen|1441,1445
recently|1446,1454
in|1455,1457
the|1458,1461
ED|1462,1464
for|1465,1468
evaluation|1469,1479
of|1480,1482
left|1483,1487
greater|1488,1495
<EOL>|1496,1497
than|1497,1501
right|1502,1507
lower|1508,1513
extremity|1514,1523
edema|1524,1529
with|1530,1534
lower|1535,1540
extremity|1541,1550
venous|1551,1557
<EOL>|1558,1559
ultrasounds|1559,1570
negative|1571,1579
,|1579,1580
without|1581,1588
change|1589,1595
in|1596,1598
edema|1599,1604
since|1605,1610
since|1611,1616
that|1617,1621
<EOL>|1622,1623
visit|1623,1628
.|1628,1629
She|1630,1633
denies|1634,1640
associated|1641,1651
fever|1652,1657
,|1657,1658
chills|1659,1665
,|1665,1666
sweats|1667,1673
,|1673,1674
PND|1675,1678
,|1678,1679
<EOL>|1680,1681
orthopnea|1681,1690
,|1690,1691
or|1692,1694
positional|1695,1705
component|1706,1715
to|1716,1718
pain|1719,1723
.|1723,1724
<EOL>|1725,1726
In|1726,1728
the|1729,1732
ED|1733,1735
,|1735,1736
initial|1737,1744
vital|1745,1750
signs|1751,1756
were|1757,1761
:|1761,1762
98.0|1763,1767
116|1768,1771
100|1772,1775
/|1775,1776
49|1776,1778
24|1779,1781
99|1782,1784
%|1784,1785
RA|1786,1788
.|1788,1789
<EOL>|1790,1791
Labs|1791,1795
notable|1796,1803
for|1804,1807
leukocytosis|1808,1820
to|1821,1823
17.9|1824,1828
,|1828,1829
hematocrit|1830,1840
of|1841,1843
32|1844,1846
,|1846,1847
and|1848,1851
<EOL>|1852,1853
lactate|1853,1860
of|1861,1863
2.8|1864,1867
.|1867,1868
Urinalysis|1869,1879
was|1880,1883
positive|1884,1892
,|1892,1893
but|1894,1897
with|1898,1902
19|1903,1905
epithelial|1906,1916
<EOL>|1917,1918
cells|1918,1923
.|1923,1924
CTA|1925,1928
was|1929,1932
negative|1933,1941
for|1942,1945
central|1946,1953
pulmonary|1954,1963
embolus|1964,1971
,|1971,1972
focal|1973,1978
<EOL>|1979,1980
consolidation|1980,1993
,|1993,1994
or|1995,1997
pleural|1998,2005
effusion|2006,2014
,|2014,2015
though|2016,2022
did|2023,2026
reveal|2027,2033
<EOL>|2034,2035
innumerable|2035,2046
pulmonary|2047,2056
nodules|2057,2064
,|2064,2065
as|2066,2068
well|2069,2073
as|2074,2076
enlarged|2077,2085
liver|2086,2091
with|2092,2096
<EOL>|2097,2098
stable|2098,2104
metastases|2105,2115
.|2115,2116
EKG|2117,2120
was|2121,2124
interpreted|2125,2136
as|2137,2139
sinus|2140,2145
tachycardia|2146,2157
and|2158,2161
<EOL>|2162,2163
was|2163,2166
overall|2167,2174
consistent|2175,2185
with|2186,2190
prior|2191,2196
.|2196,2197
Ceftriaxone|2198,2209
/|2209,2210
azithromycin|2210,2222
were|2223,2227
<EOL>|2228,2229
initiated|2229,2238
for|2239,2242
possible|2243,2251
pneumonia|2252,2261
.|2261,2262
Vital|2263,2268
signs|2269,2274
on|2275,2277
transfer|2279,2287
were|2288,2292
<EOL>|2293,2294
as|2294,2296
follows|2297,2304
:|2304,2305
97.9|2306,2310
107|2311,2314
100|2315,2318
/|2318,2319
60|2319,2321
22|2322,2324
100|2325,2328
%|2328,2329
RA|2330,2332
.|2332,2333
On|2334,2336
arrival|2337,2344
to|2345,2347
the|2348,2351
floor|2352,2357
,|2357,2358
<EOL>|2359,2360
she|2360,2363
reports|2364,2371
that|2372,2376
shortness|2377,2386
of|2387,2389
breath|2390,2396
has|2397,2400
improved|2401,2409
and|2410,2413
that|2414,2418
she|2419,2422
<EOL>|2423,2424
is|2424,2426
chest|2427,2432
pain|2433,2437
free|2438,2442
.|2442,2443
<EOL>|2443,2444
<EOL>|2445,2446
Per|2468,2471
OMR|2472,2475
:|2475,2476
<EOL>|2476,2477
#|2477,2478
metastatic|2479,2489
cancer|2490,2496
of|2497,2499
unknown|2500,2507
primary|2508,2515
<EOL>|2515,2516
#|2516,2517
high|2518,2522
grade|2523,2528
SBO|2529,2532
_|2533,2534
_|2534,2535
_|2535,2536
s|2537,2538
/|2538,2539
p|2539,2540
exploratory|2541,2552
laparotomy|2553,2563
,|2563,2564
lysis|2565,2570
of|2571,2573
<EOL>|2574,2575
adhesions|2575,2584
,|2584,2585
and|2586,2589
small|2590,2595
bowel|2596,2601
resection|2602,2611
with|2612,2616
enteroenterostomy|2617,2634
<EOL>|2635,2636
#|2636,2637
carcinoid|2638,2647
<EOL>|2647,2648
#|2648,2649
hyperlipidemia|2650,2664
<EOL>|2664,2665
#|2665,2666
vitamin|2667,2674
B12|2675,2678
deficiency|2679,2689
<EOL>|2689,2690
#|2690,2691
cervical|2692,2700
DJD|2701,2704
<EOL>|2704,2705
#|2705,2706
osteoarthritis|2707,2721
<EOL>|2722,2723
<EOL>|2723,2724
s|2724,2725
/|2725,2726
p|2726,2727
R|2728,2729
lung|2730,2734
resection|2735,2744
in|2745,2747
_|2748,2749
_|2749,2750
_|2750,2751
at|2752,2754
_|2755,2756
_|2756,2757
_|2757,2758
<EOL>|2758,2759
s|2759,2760
/|2760,2761
p|2761,2762
hysterectomy|2763,2775
in|2776,2778
_|2779,2780
_|2780,2781
_|2781,2782
<EOL>|2782,2783
s|2783,2784
/|2784,2785
p|2785,2786
R|2787,2788
arm|2789,2792
surgery|2793,2800
<EOL>|2800,2801
<EOL>|2801,2802
<EOL>|2803,2804
:|2818,2819
<EOL>|2819,2820
_|2820,2821
_|2821,2822
_|2822,2823
<EOL>|2823,2824
:|2838,2839
<EOL>|2839,2840
Per|2840,2843
OMR|2844,2847
:|2847,2848
<EOL>|2848,2849
Mother|2849,2855
-|2856,2857
Died|2858,2862
of|2863,2865
pancreatic|2866,2876
cancer|2877,2883
at|2884,2886
age|2887,2890
_|2891,2892
_|2892,2893
_|2893,2894
.|2894,2895
<EOL>|2897,2898
Father|2898,2904
-|2905,2906
Died|2907,2911
of|2912,2914
_|2915,2916
_|2916,2917
_|2917,2918
disease|2919,2926
at|2927,2929
age|2930,2933
_|2934,2935
_|2935,2936
_|2936,2937
.|2937,2938
<EOL>|2939,2940
<EOL>|2941,2942
On|2957,2959
admission|2960,2969
:|2969,2970
<EOL>|2970,2971
VS|2971,2973
:|2973,2974
97.9|2975,2979
114|2980,2983
/|2983,2984
71|2984,2986
105|2987,2990
sinus|2991,2996
18|2997,2999
95|3000,3002
%|3002,3003
2L|3003,3005
<EOL>|3007,3008
GENERAL|3008,3015
:|3015,3016
non-toxic|3017,3026
appearing|3027,3036
,|3036,3037
speaking|3038,3046
in|3047,3049
full|3050,3054
sentences|3055,3064
<EOL>|3066,3067
HEENT|3067,3072
:|3072,3073
NC|3074,3076
/|3076,3077
AT|3077,3079
,|3079,3080
PERRLA|3081,3087
,|3087,3088
EOMI|3089,3093
,|3093,3094
sclerae|3095,3102
anicteric|3103,3112
,|3112,3113
MMM|3114,3117
<EOL>|3119,3120
NECK|3120,3124
:|3124,3125
supple|3126,3132
,|3132,3133
no|3134,3136
LAD|3137,3140
,|3140,3141
no|3142,3144
JVD|3145,3148
<EOL>|3150,3151
CHEST|3151,3156
:|3156,3157
mild|3158,3162
reproducible|3163,3175
pain|3176,3180
on|3181,3183
palp|3184,3188
of|3189,3191
midsternum|3192,3202
;|3202,3203
no|3204,3206
palpable|3207,3215
<EOL>|3216,3217
mass|3217,3221
<EOL>|3223,3224
LUNGS|3224,3229
:|3229,3230
poor|3231,3235
aeration|3236,3244
but|3245,3248
relatively|3249,3259
CTA|3260,3263
bilat|3264,3269
,|3269,3270
no|3271,3273
r|3274,3275
/|3275,3276
rh|3276,3278
/|3278,3279
wh|3279,3281
,|3281,3282
resp|3283,3287
<EOL>|3288,3289
unlabored|3289,3298
,|3298,3299
no|3300,3302
accessory|3303,3312
muscle|3313,3319
use|3320,3323
<EOL>|3325,3326
HEART|3326,3331
:|3331,3332
clear|3333,3338
and|3339,3342
audible|3343,3350
heart|3351,3356
sounds|3357,3363
,|3363,3364
tachycardiac|3365,3377
but|3378,3381
regular|3382,3389
<EOL>|3390,3391
rhythm|3391,3397
,|3397,3398
sofy|3399,3403
SEM|3404,3407
,|3407,3408
nl|3409,3411
S1|3412,3414
-|3414,3415
S2|3415,3417
<EOL>|3419,3420
ABDOMEN|3420,3427
:|3427,3428
normal|3429,3435
bowel|3436,3441
sounds|3442,3448
,|3448,3449
soft|3450,3454
,|3454,3455
mild|3456,3460
tenderness|3461,3471
to|3472,3474
palp|3475,3479
<EOL>|3480,3481
throughout|3481,3491
and|3492,3495
more|3496,3500
pronounced|3501,3511
in|3512,3514
the|3515,3518
RUQ|3519,3522
,|3522,3523
non-distended|3524,3537
,|3537,3538
no|3539,3541
<EOL>|3542,3543
rebound|3543,3550
or|3551,3553
guarding|3554,3562
,|3562,3563
palpable|3564,3572
liver|3573,3578
edge|3579,3583
<EOL>|3585,3586
EXTREMITIES|3586,3597
:|3597,3598
left|3599,3603
>|3604,3605
right|3606,3611
1|3612,3613
+|3613,3614
pitting|3615,3622
edema|3623,3628
to|3629,3631
mid|3632,3635
shin|3636,3640
,|3640,3641
2|3642,3643
+|3643,3644
<EOL>|3645,3646
pulses|3646,3652
radial|3653,3659
and|3660,3663
dp|3664,3666
<EOL>|3668,3669
NEURO|3669,3674
:|3674,3675
awake|3676,3681
,|3681,3682
A|3683,3684
&|3684,3685
Ox3|3685,3688
,|3688,3689
CNs|3690,3693
II|3694,3696
-|3696,3697
XII|3697,3700
grossly|3701,3708
intact|3709,3715
,|3715,3716
muscle|3717,3723
strength|3724,3732
<EOL>|3733,3734
_|3734,3735
_|3735,3736
_|3736,3737
throughout|3738,3748
,|3748,3749
sensation|3750,3759
grossly|3760,3767
intact|3768,3774
<EOL>|3774,3775
<EOL>|3775,3776
At|3776,3778
discharge|3779,3788
:|3788,3789
<EOL>|3789,3790
VS|3790,3792
-|3793,3794
Tc|3795,3797
99.7|3798,3802
,|3802,3803
116|3804,3807
/|3807,3808
59|3808,3810
,|3810,3811
131|3812,3815
,|3815,3816
18|3817,3819
,|3819,3820
99|3821,3823
%|3823,3824
RA|3825,3827
<EOL>|3827,3828
GENERAL|3828,3835
:|3835,3836
obese|3837,3842
,|3842,3843
NAD|3844,3847
,|3847,3848
lying|3849,3854
in|3855,3857
bed|3858,3861
comfortably|3862,3873
,|3873,3874
flat|3875,3879
affect|3880,3886
and|3887,3890
<EOL>|3891,3892
poor|3892,3896
eye|3897,3900
contact|3901,3908
<EOL>|3908,3909
HEENT|3909,3914
:|3914,3915
NCAT|3916,3920
,|3920,3921
EOMI|3922,3926
,|3926,3927
mild|3928,3932
scleral|3933,3940
icterus|3941,3948
,|3948,3949
pink|3950,3954
conjunctiva|3955,3966
,|3966,3967
MMM|3968,3971
,|3971,3972
<EOL>|3973,3974
poor|3974,3978
dentition|3979,3988
,|3988,3989
mild|3990,3994
palor|3995,4000
of|4001,4003
conjunctiva|4004,4015
<EOL>|4016,4017
NECK|4017,4021
:|4021,4022
supple|4023,4029
,|4029,4030
no|4031,4033
LAD|4034,4037
<EOL>|4039,4040
CARDIAC|4040,4047
:|4047,4048
tachycardic|4049,4060
but|4061,4064
regular|4065,4072
,|4072,4073
S1|4074,4076
/|4076,4077
S2|4077,4079
,|4079,4080
no|4081,4083
m|4084,4085
/|4085,4086
r|4086,4087
/|4087,4088
g|4088,4089
<EOL>|4089,4090
LUNG|4090,4094
:|4094,4095
CTAB|4096,4100
in|4101,4103
anterior|4104,4112
fields|4113,4119
,|4119,4120
decreased|4121,4130
breath|4131,4137
sounds|4138,4144
at|4145,4147
right|4148,4153
<EOL>|4154,4155
base|4155,4159
,|4159,4160
exam|4161,4165
limited|4166,4173
secondary|4174,4183
to|4184,4186
body|4187,4191
habitus|4192,4199
and|4200,4203
mobility|4204,4212
,|4212,4213
no|4214,4216
<EOL>|4217,4218
w|4218,4219
/|4219,4220
r|4220,4221
/|4221,4222
r|4222,4223
,|4223,4224
no|4225,4227
accessory|4228,4237
muscle|4238,4244
use|4245,4248
<EOL>|4248,4249
ABDOMEN|4249,4256
:|4256,4257
obese|4258,4263
,|4263,4264
ND|4265,4267
,|4267,4268
+|4269,4270
BS|4270,4272
,|4272,4273
no|4274,4276
rebound|4277,4284
/|4284,4285
guarding|4285,4293
,|4293,4294
localized|4295,4304
area|4305,4309
of|4310,4312
<EOL>|4313,4314
firmness|4314,4322
in|4323,4325
mid-upper|4326,4335
abdomen|4336,4343
and|4344,4347
tender|4348,4354
to|4355,4357
palpation|4358,4367
over|4368,4372
this|4373,4377
<EOL>|4378,4379
area|4379,4383
<EOL>|4384,4385
EXTREMITIES|4385,4396
:|4396,4397
WWP|4398,4401
,|4401,4402
2|4403,4404
+|4404,4405
DP|4406,4408
pulses|4409,4415
bilaterally|4416,4427
,|4427,4428
1|4429,4430
+|4430,4431
pitting|4432,4439
edema|4440,4445
to|4446,4448
<EOL>|4449,4450
torso|4450,4455
bilateraly|4456,4466
<EOL>|4467,4468
NEURO|4468,4473
:|4473,4474
no|4475,4477
asterixis|4478,4487
,|4487,4488
moving|4489,4495
all|4496,4499
four|4500,4504
extremities|4505,4516
,|4516,4517
minimal|4518,4525
<EOL>|4526,4527
movement|4527,4535
_|4536,4537
_|4537,4538
_|4538,4539
to|4540,4542
gravity|4543,4550
but|4551,4554
distal|4555,4561
muscles|4562,4569
4|4570,4571
+|4571,4572
/|4572,4573
5|4573,4574
,|4574,4575
good|4576,4580
hand|4581,4585
<EOL>|4586,4587
grip|4587,4591
strength|4592,4600
today|4601,4606
<EOL>|4606,4607
<EOL>|4608,4609
Pertinent|4609,4618
Results|4619,4626
:|4626,4627
<EOL>|4627,4628
On|4628,4630
admission|4631,4640
:|4640,4641
<EOL>|4641,4642
_|4642,4643
_|4643,4644
_|4644,4645
12|4646,4648
:|4648,4649
50PM|4649,4653
BLOOD|4654,4659
WBC|4660,4663
-|4663,4664
17|4664,4666
.|4666,4667
9|4667,4668
*|4668,4669
RBC|4670,4673
-|4673,4674
3|4674,4675
.|4675,4676
69|4676,4678
*|4678,4679
Hgb|4680,4683
-|4683,4684
9|4684,4685
.|4685,4686
5|4686,4687
*|4687,4688
Hct|4689,4692
-|4692,4693
32|4693,4695
.|4695,4696
1|4696,4697
*|4697,4698
<EOL>|4699,4700
MCV|4700,4703
-|4703,4704
87|4704,4706
MCH|4707,4710
-|4710,4711
25|4711,4713
.|4713,4714
8|4714,4715
*|4715,4716
MCHC|4717,4721
-|4721,4722
29|4722,4724
.|4724,4725
7|4725,4726
*|4726,4727
RDW|4728,4731
-|4731,4732
19|4732,4734
.|4734,4735
1|4735,4736
*|4736,4737
Plt|4738,4741
_|4742,4743
_|4743,4744
_|4744,4745
<EOL>|4745,4746
_|4746,4747
_|4747,4748
_|4748,4749
12|4750,4752
:|4752,4753
50PM|4753,4757
BLOOD|4758,4763
Neuts|4764,4769
-|4769,4770
82|4770,4772
.|4772,4773
8|4773,4774
*|4774,4775
Lymphs|4776,4782
-|4782,4783
11|4783,4785
.|4785,4786
7|4786,4787
*|4787,4788
Monos|4789,4794
-|4794,4795
4.4|4795,4798
<EOL>|4799,4800
Eos|4800,4803
-|4803,4804
0.7|4804,4807
Baso|4808,4812
-|4812,4813
0.3|4813,4816
<EOL>|4816,4817
_|4817,4818
_|4818,4819
_|4819,4820
12|4821,4823
:|4823,4824
50PM|4824,4828
BLOOD|4829,4834
_|4835,4836
_|4836,4837
_|4837,4838
PTT|4839,4842
-|4842,4843
31.2|4843,4847
_|4848,4849
_|4849,4850
_|4850,4851
<EOL>|4851,4852
_|4852,4853
_|4853,4854
_|4854,4855
12|4856,4858
:|4858,4859
50PM|4859,4863
BLOOD|4864,4869
Glucose|4870,4877
-|4877,4878
97|4878,4880
UreaN|4881,4886
-|4886,4887
12|4887,4889
Creat|4890,4895
-|4895,4896
0.6|4896,4899
Na|4900,4902
-|4902,4903
140|4903,4906
<EOL>|4907,4908
K|4908,4909
-|4909,4910
2|4910,4911
.|4911,4912
7|4912,4913
*|4913,4914
Cl|4915,4917
-|4917,4918
92|4918,4920
*|4920,4921
HCO3|4922,4926
-|4926,4927
31|4927,4929
AnGap|4930,4935
-|4935,4936
20|4936,4938
<EOL>|4938,4939
_|4939,4940
_|4940,4941
_|4941,4942
12|4943,4945
:|4945,4946
50PM|4946,4950
BLOOD|4951,4956
ALT|4957,4960
-|4960,4961
17|4961,4963
AST|4964,4967
-|4967,4968
73|4968,4970
*|4970,4971
LD|4972,4974
(|4974,4975
_|4975,4976
_|4976,4977
_|4977,4978
)|4978,4979
-|4979,4980
586|4980,4983
*|4983,4984
CK|4985,4987
(|4987,4988
CPK|4988,4991
)|4991,4992
-|4992,4993
218|4993,4996
*|4996,4997
<EOL>|4998,4999
AlkPhos|4999,5006
-|5006,5007
340|5007,5010
*|5010,5011
TotBili|5012,5019
-|5019,5020
2|5020,5021
.|5021,5022
6|5022,5023
*|5023,5024
DirBili|5025,5032
-|5032,5033
1|5033,5034
.|5034,5035
8|5035,5036
*|5036,5037
IndBili|5038,5045
-|5045,5046
0.8|5046,5049
<EOL>|5049,5050
_|5050,5051
_|5051,5052
_|5052,5053
12|5054,5056
:|5056,5057
50PM|5057,5061
BLOOD|5062,5067
CK|5068,5070
-|5070,5071
MB|5071,5073
-|5073,5074
1|5074,5075
cTropnT|5076,5083
-|5083,5084
<|5084,5085
0|5085,5086
.|5086,5087
01|5087,5089
<EOL>|5089,5090
_|5090,5091
_|5091,5092
_|5092,5093
12|5094,5096
:|5096,5097
50PM|5097,5101
BLOOD|5102,5107
Albumin|5108,5115
-|5115,5116
2|5116,5117
.|5117,5118
5|5118,5119
*|5119,5120
Mg|5121,5123
-|5123,5124
2.2|5124,5127
<EOL>|5127,5128
_|5128,5129
_|5129,5130
_|5130,5131
12|5132,5134
:|5134,5135
50PM|5135,5139
BLOOD|5140,5145
Hapto|5146,5151
-|5151,5152
307|5152,5155
*|5155,5156
<EOL>|5156,5157
_|5157,5158
_|5158,5159
_|5159,5160
05|5161,5163
:|5163,5164
12PM|5164,5168
BLOOD|5169,5174
Lactate|5175,5182
-|5182,5183
2|5183,5184
.|5184,5185
8|5185,5186
*|5186,5187
<EOL>|5187,5188
<EOL>|5188,5189
_|5189,5190
_|5190,5191
_|5191,5192
06|5193,5195
:|5195,5196
00PM|5196,5200
URINE|5201,5206
Color|5207,5212
-|5212,5213
YELLOW|5213,5219
Appear|5220,5226
-|5226,5227
Cloudy|5227,5233
Sp|5234,5236
_|5237,5238
_|5238,5239
_|5239,5240
<EOL>|5240,5241
_|5241,5242
_|5242,5243
_|5243,5244
06|5245,5247
:|5247,5248
00PM|5248,5252
URINE|5253,5258
Blood|5259,5264
-|5264,5265
NEG|5265,5268
Nitrite|5269,5276
-|5276,5277
NEG|5277,5280
Protein|5281,5288
-|5288,5289
30|5289,5291
<EOL>|5292,5293
Glucose|5293,5300
-|5300,5301
NEG|5301,5304
Ketone|5305,5311
-|5311,5312
10|5312,5314
Bilirub|5315,5322
-|5322,5323
SM|5323,5325
Urobiln|5327,5334
-|5334,5335
8|5335,5336
*|5336,5337
pH|5338,5340
-|5340,5341
6.0|5341,5344
Leuks|5345,5350
-|5350,5351
MOD|5351,5354
<EOL>|5354,5355
_|5355,5356
_|5356,5357
_|5357,5358
06|5359,5361
:|5361,5362
00PM|5362,5366
URINE|5367,5372
RBC|5373,5376
-|5376,5377
0|5377,5378
WBC|5379,5382
-|5382,5383
66|5383,5385
*|5385,5386
Bacteri|5387,5394
-|5394,5395
FEW|5395,5398
Yeast|5399,5404
-|5404,5405
NONE|5405,5409
<EOL>|5410,5411
Epi|5411,5414
-|5414,5415
14|5415,5417
<EOL>|5417,5418
_|5418,5419
_|5419,5420
_|5420,5421
06|5422,5424
:|5424,5425
00PM|5425,5429
URINE|5430,5435
CastHy|5436,5442
-|5442,5443
6|5443,5444
*|5444,5445
<EOL>|5445,5446
<EOL>|5446,5447
At|5447,5449
discharge|5450,5459
:|5459,5460
<EOL>|5460,5461
_|5461,5462
_|5462,5463
_|5463,5464
08|5465,5467
:|5467,5468
30AM|5468,5472
BLOOD|5473,5478
WBC|5479,5482
-|5482,5483
16|5483,5485
.|5485,5486
1|5486,5487
*|5487,5488
RBC|5489,5492
-|5492,5493
3|5493,5494
.|5494,5495
06|5495,5497
*|5497,5498
Hgb|5499,5502
-|5502,5503
8|5503,5504
.|5504,5505
3|5505,5506
*|5506,5507
Hct|5508,5511
-|5511,5512
29|5512,5514
.|5514,5515
2|5515,5516
*|5516,5517
<EOL>|5518,5519
MCV|5519,5522
-|5522,5523
95|5523,5525
MCH|5526,5529
-|5529,5530
27.1|5530,5534
MCHC|5535,5539
-|5539,5540
28|5540,5542
.|5542,5543
5|5543,5544
*|5544,5545
RDW|5546,5549
-|5549,5550
22|5550,5552
.|5552,5553
5|5553,5554
*|5554,5555
Plt|5556,5559
_|5560,5561
_|5561,5562
_|5562,5563
<EOL>|5563,5564
_|5564,5565
_|5565,5566
_|5566,5567
08|5568,5570
:|5570,5571
30AM|5571,5575
BLOOD|5576,5581
Glucose|5582,5589
-|5589,5590
95|5590,5592
UreaN|5593,5598
-|5598,5599
7|5599,5600
Creat|5601,5606
-|5606,5607
0|5607,5608
.|5608,5609
3|5609,5610
*|5610,5611
Na|5612,5614
-|5614,5615
143|5615,5618
<EOL>|5619,5620
K|5620,5621
-|5621,5622
3.5|5622,5625
Cl|5626,5628
-|5628,5629
110|5629,5632
*|5632,5633
HCO3|5634,5638
-|5638,5639
20|5639,5641
*|5641,5642
AnGap|5643,5648
-|5648,5649
17|5649,5651
<EOL>|5651,5652
_|5652,5653
_|5653,5654
_|5654,5655
08|5656,5658
:|5658,5659
30AM|5659,5663
BLOOD|5664,5669
Calcium|5670,5677
-|5677,5678
8|5678,5679
.|5679,5680
3|5680,5681
*|5681,5682
Phos|5683,5687
-|5687,5688
2|5688,5689
.|5689,5690
4|5690,5691
*|5691,5692
Mg|5693,5695
-|5695,5696
1.9|5696,5699
<EOL>|5699,5700
<EOL>|5700,5701
Microbiology|5701,5713
:|5713,5714
<EOL>|5714,5715
Blood|5715,5720
x2|5721,5723
(|5724,5725
_|5725,5726
_|5726,5727
_|5727,5728
)|5728,5729
:|5729,5730
No|5731,5733
growth|5734,5740
<EOL>|5740,5741
Urine|5741,5746
(|5747,5748
_|5748,5749
_|5749,5750
_|5750,5751
)|5751,5752
:|5752,5753
No|5754,5756
growth|5757,5763
<EOL>|5763,5764
Blood|5764,5769
x2|5770,5772
(|5773,5774
_|5774,5775
_|5775,5776
_|5776,5777
)|5777,5778
:|5778,5779
No|5780,5782
growth|5783,5789
<EOL>|5789,5790
<EOL>|5790,5791
Pathology|5791,5800
:|5800,5801
<EOL>|5801,5802
Liver|5802,5807
biopsy|5808,5814
(|5815,5816
_|5816,5817
_|5817,5818
_|5818,5819
)|5819,5820
:|5820,5821
<EOL>|5821,5822
Liver|5822,5827
,|5827,5828
core|5829,5833
needle|5834,5840
biopsy|5841,5847
(|5848,5849
A|5849,5850
)|5850,5851
:|5851,5852
<EOL>|5852,5853
Adenocarcinoma|5853,5867
,|5867,5868
involving|5869,5878
the|5879,5882
liver|5883,5888
(|5889,5890
see|5890,5893
note|5894,5898
)|5898,5899
.|5899,5900
<EOL>|5900,5901
Note|5901,5905
:|5905,5906
Immunohistochemical|5907,5926
stains|5927,5933
are|5934,5937
performed|5938,5947
.|5947,5948
The|5950,5953
tumor|5954,5959
cells|5960,5965
<EOL>|5966,5967
are|5967,5970
positive|5971,5979
for|5980,5983
CK20|5984,5988
and|5989,5992
CDX|5993,5996
-|5996,5997
2|5997,5998
,|5998,5999
and|6000,6003
negative|6004,6012
for|6013,6016
CK7|6017,6020
and|6021,6024
TTF|6025,6028
-|6028,6029
1|6029,6030
.|6030,6031
<EOL>|6032,6033
These|6034,6039
results|6040,6047
are|6048,6051
consistent|6052,6062
with|6063,6067
metastasis|6068,6078
from|6079,6083
a|6084,6085
colorectal|6086,6096
<EOL>|6097,6098
primary|6098,6105
.|6105,6106
<EOL>|6106,6107
<EOL>|6107,6108
Imaging|6108,6115
:|6115,6116
<EOL>|6116,6117
EKG|6117,6120
(|6121,6122
_|6122,6123
_|6123,6124
_|6124,6125
)|6125,6126
:|6126,6127
<EOL>|6127,6128
Sinus|6128,6133
tachycardia|6134,6145
.|6145,6146
Low|6147,6150
voltage|6151,6158
.|6158,6159
Diffuse|6160,6167
non-specific|6168,6180
<EOL>|6181,6182
repolarization|6182,6196
<EOL>|6196,6197
abnormalities|6197,6210
.|6210,6211
Compared|6212,6220
to|6221,6223
the|6224,6227
previous|6228,6236
tracing|6237,6244
of|6245,6247
_|6248,6249
_|6249,6250
_|6250,6251
<EOL>|6252,6253
repolarization|6253,6267
<EOL>|6267,6268
abnormalities|6268,6281
are|6282,6285
slightly|6286,6294
more|6295,6299
prominent|6300,6309
.|6309,6310
<EOL>|6310,6311
_|6311,6312
_|6312,6313
_|6313,6314
<EOL>|6314,6315
_|6315,6316
_|6316,6317
_|6317,6318
<EOL>|6318,6319
<EOL>|6319,6320
Portable|6320,6328
CXR|6329,6332
(|6333,6334
_|6334,6335
_|6335,6336
_|6336,6337
)|6337,6338
:|6338,6339
<EOL>|6339,6340
Innumerable|6340,6351
pulmonary|6352,6361
metastases|6362,6372
.|6372,6373
Possible|6375,6383
mild|6384,6388
pulmonary|6389,6398
<EOL>|6399,6400
vascular|6400,6408
<EOL>|6408,6409
congestion|6409,6419
.|6419,6420
Low|6422,6425
lung|6426,6430
volumes|6431,6438
.|6438,6439
<EOL>|6439,6440
<EOL>|6440,6441
CTA|6441,6444
(|6445,6446
_|6446,6447
_|6447,6448
_|6448,6449
)|6449,6450
:|6450,6451
<EOL>|6451,6452
1|6452,6453
.|6453,6454
No|6456,6458
central|6459,6466
or|6467,6469
segmental|6470,6479
filling|6480,6487
defect|6488,6494
in|6495,6497
the|6498,6501
pulmonary|6502,6511
<EOL>|6512,6513
arteries|6513,6521
.|6521,6522
<EOL>|6522,6523
Evaluation|6523,6533
is|6534,6536
slightly|6537,6545
limited|6546,6553
due|6554,6557
to|6558,6560
suboptimal|6561,6571
IV|6572,6574
bolus|6575,6580
.|6580,6581
<EOL>|6582,6583
2.|6583,6585
Innumerable|6587,6598
bilateral|6599,6608
pulmonary|6609,6618
nodules|6619,6626
,|6626,6627
simas|6628,6633
seen|6634,6638
on|6639,6641
the|6642,6645
<EOL>|6646,6647
prior|6647,6652
CT|6653,6655
study|6656,6661
on|6662,6664
_|6665,6666
_|6666,6667
_|6667,6668
,|6668,6669
slightly|6670,6678
increased|6679,6688
.|6688,6689
No|6691,6693
focal|6694,6699
<EOL>|6700,6701
consolidation|6701,6714
or|6715,6717
pleural|6718,6725
effusion|6726,6734
.|6734,6735
<EOL>|6737,6738
3.|6738,6740
Enlarged|6742,6750
liver|6751,6756
with|6757,6761
multiple|6762,6770
hypodense|6771,6780
lesions|6781,6788
,|6788,6789
with|6790,6794
<EOL>|6795,6796
suggestion|6796,6806
of|6807,6809
<EOL>|6809,6810
increased|6810,6819
burden|6820,6826
of|6827,6829
disease|6830,6837
.|6837,6838
<EOL>|6838,6839
<EOL>|6839,6840
Right|6840,6845
upper|6846,6851
quadrant|6852,6860
ultrasound|6861,6871
(|6872,6873
_|6873,6874
_|6874,6875
_|6875,6876
)|6876,6877
:|6877,6878
<EOL>|6878,6879
Extensive|6879,6888
diffuse|6889,6896
hepatic|6897,6904
metastatic|6905,6915
disease|6916,6923
.|6923,6924
No|6926,6928
evidence|6929,6937
of|6938,6940
<EOL>|6941,6942
biliary|6942,6949
duct|6950,6954
<EOL>|6954,6955
obstruction|6955,6966
.|6966,6967
<EOL>|6967,6968
<EOL>|6968,6969
Portable|6969,6977
CXR|6978,6981
(|6982,6983
_|6983,6984
_|6984,6985
_|6985,6986
)|6986,6987
:|6987,6988
<EOL>|6988,6989
1.|6989,6991
Low|6992,6995
lung|6996,7000
volumes|7001,7008
and|7009,7012
mild|7013,7017
pulmonary|7018,7027
vascular|7028,7036
congestion|7037,7047
is|7048,7050
<EOL>|7051,7052
unchanged|7052,7061
.|7061,7062
<EOL>|7063,7064
2.|7064,7066
New|7067,7070
small|7071,7076
right|7077,7082
fissural|7083,7091
pleural|7092,7099
effusion|7100,7108
.|7108,7109
<EOL>|7109,7110
3.|7110,7112
No|7113,7115
new|7116,7119
focal|7120,7125
opacities|7126,7135
to|7136,7138
suggest|7139,7146
pneumonia|7147,7156
.|7156,7157
<EOL>|7159,7160
<EOL>|7160,7161
Noncontrast|7161,7172
head|7173,7177
CT|7178,7180
(|7181,7182
_|7182,7183
_|7183,7184
_|7184,7185
)|7185,7186
:|7186,7187
<EOL>|7187,7188
No|7188,7190
acute|7191,7196
intracranial|7197,7209
process|7210,7217
.|7217,7218
No|7220,7222
mass|7223,7227
is|7228,7230
identified|7231,7241
.|7241,7242
MRI|7244,7247
is|7248,7250
<EOL>|7251,7252
more|7252,7256
sensitive|7257,7266
for|7267,7270
evaluation|7271,7281
of|7282,7284
metastases|7285,7295
.|7295,7296
<EOL>|7296,7297
<EOL>|7297,7298
Left|7298,7302
hip|7303,7306
XR|7307,7309
(|7310,7311
_|7311,7312
_|7312,7313
_|7313,7314
)|7314,7315
:|7315,7316
<EOL>|7316,7317
No|7317,7319
definite|7320,7328
lytic|7329,7334
lesion|7335,7341
;|7341,7342
however|7343,7350
,|7350,7351
an|7352,7354
MRI|7355,7358
can|7359,7362
be|7363,7365
performed|7366,7375
to|7376,7378
<EOL>|7379,7380
evaluate|7380,7388
for|7389,7392
an|7393,7395
osseous|7396,7403
lesion|7404,7410
if|7411,7413
indicated|7414,7423
.|7423,7424
<EOL>|7424,7425
<EOL>|7425,7426
Portable|7426,7434
abdomen|7435,7442
(|7443,7444
_|7444,7445
_|7445,7446
_|7446,7447
)|7447,7448
:|7448,7449
<EOL>|7449,7450
Radiographs|7450,7461
of|7462,7464
the|7465,7468
abdomen|7469,7476
and|7477,7480
pelvis|7481,7487
demonstrate|7488,7499
a|7500,7501
<EOL>|7502,7503
nonobstructed|7503,7516
<EOL>|7516,7517
bowel|7517,7522
gas|7523,7526
pattern|7527,7534
.|7534,7535
A|7537,7538
relative|7539,7547
paucity|7548,7555
of|7556,7558
bowel|7559,7564
gas|7565,7568
is|7569,7571
present|7572,7579
<EOL>|7580,7581
in|7581,7583
the|7584,7587
upper|7588,7593
and|7594,7597
mid|7598,7601
abdomen|7602,7609
,|7609,7610
likely|7611,7617
due|7618,7621
to|7622,7624
marked|7625,7631
enlargement|7632,7643
<EOL>|7644,7645
of|7645,7647
the|7648,7651
liver|7652,7657
,|7657,7658
displacing|7659,7669
bowel|7670,7675
loops|7676,7681
.|7681,7682
Note|7684,7688
that|7689,7693
the|7694,7697
upright|7698,7705
<EOL>|7706,7707
view|7707,7711
is|7712,7714
technically|7715,7726
suboptimal|7727,7737
,|7737,7738
and|7739,7742
limits|7743,7749
evaluation|7750,7760
for|7761,7764
free|7765,7769
<EOL>|7770,7771
intraperitoneal|7771,7786
air|7787,7790
.|7790,7791
If|7793,7795
free|7796,7800
intraperitoneal|7801,7816
air|7817,7820
is|7821,7823
suspected|7824,7833
<EOL>|7834,7835
clinically|7835,7845
,|7845,7846
a|7847,7848
left|7849,7853
lateral|7854,7861
decubitus|7862,7871
view|7872,7876
of|7877,7879
the|7880,7883
abdomen|7884,7891
would|7892,7897
<EOL>|7898,7899
be|7899,7901
recommended|7902,7913
.|7913,7914
<EOL>|7914,7915
<EOL>|7916,7917
Ms.|7940,7943
_|7944,7945
_|7945,7946
_|7946,7947
is|7948,7950
a|7951,7952
_|7953,7954
_|7954,7955
_|7955,7956
with|7957,7961
metastatic|7962,7972
cancer|7973,7979
of|7980,7982
unknown|7983,7990
primary|7991,7998
,|7998,7999
<EOL>|8000,8001
including|8001,8010
lesions|8011,8018
in|8019,8021
the|8022,8025
liver|8026,8031
and|8032,8035
lungs|8036,8041
,|8041,8042
who|8043,8046
initially|8047,8056
<EOL>|8057,8058
presented|8058,8067
with|8068,8072
shortness|8073,8082
of|8083,8085
breath|8086,8092
,|8092,8093
likely|8094,8100
due|8101,8104
to|8105,8107
worsening|8108,8117
<EOL>|8118,8119
intrapulmonary|8119,8133
tumor|8134,8139
burden|8140,8146
,|8146,8147
and|8148,8151
later|8152,8157
underwent|8158,8167
percutaneous|8168,8180
<EOL>|8181,8182
liver|8182,8187
biopsy|8188,8194
with|8195,8199
pathology|8200,8209
consistent|8210,8220
with|8221,8225
metastatic|8226,8236
colon|8237,8242
<EOL>|8243,8244
cancer|8244,8250
,|8250,8251
prompting|8252,8261
transfer|8262,8270
to|8271,8273
the|8274,8277
oncology|8278,8286
service|8287,8294
and|8295,8298
<EOL>|8299,8300
eventually|8300,8310
discharged|8311,8321
home|8322,8326
with|8327,8331
hospice|8332,8339
.|8339,8340
<EOL>|8340,8341
<EOL>|8341,8342
Active|8342,8348
Issues|8349,8355
:|8355,8356
<EOL>|8356,8357
(|8357,8358
1|8358,8359
)|8359,8360
Metastatic|8361,8371
colon|8372,8377
adenocarcinoma|8378,8392
:|8392,8393
CTA|8394,8397
to|8398,8400
exclude|8401,8408
pulmonary|8409,8418
<EOL>|8419,8420
embolus|8420,8427
and|8428,8431
right|8432,8437
upper|8438,8443
quadrant|8444,8452
ultrasound|8453,8463
on|8464,8466
admission|8467,8476
<EOL>|8477,8478
demonstrated|8478,8490
progression|8491,8502
of|8503,8505
previously|8506,8516
recognized|8517,8527
metastatic|8528,8538
<EOL>|8539,8540
cancer|8540,8546
of|8547,8549
unknown|8550,8557
primary|8558,8565
involving|8566,8575
the|8576,8579
liver|8580,8585
and|8586,8589
lungs|8590,8595
,|8595,8596
which|8597,8602
<EOL>|8603,8604
had|8604,8607
evaded|8608,8614
diagnosis|8615,8624
in|8625,8627
the|8628,8631
outpatient|8632,8642
setting|8643,8650
due|8651,8654
to|8655,8657
patient|8658,8665
<EOL>|8666,8667
reluctance|8667,8677
to|8678,8680
engage|8681,8687
with|8688,8692
care|8693,8697
.|8697,8698
Percutaneous|8699,8711
liver|8712,8717
biopsy|8718,8724
<EOL>|8725,8726
ultimately|8726,8736
revealed|8737,8745
primary|8746,8753
colonic|8754,8761
adenocarcinoma|8762,8776
.|8776,8777
Following|8778,8787
<EOL>|8788,8789
discussion|8789,8799
with|8800,8804
her|8805,8808
outpatient|8809,8819
oncology|8820,8828
providers|8829,8838
,|8838,8839
she|8840,8843
was|8844,8847
<EOL>|8848,8849
transferred|8849,8860
to|8861,8863
the|8864,8867
inpatient|8868,8877
oncology|8878,8886
service|8887,8894
for|8895,8898
potential|8899,8908
<EOL>|8909,8910
trial|8910,8915
of|8916,8918
FLOX|8919,8923
.|8923,8924
However|8925,8932
,|8932,8933
given|8934,8939
the|8940,8943
patient|8944,8951
's|8951,8953
very|8954,8958
poor|8959,8963
functional|8964,8974
<EOL>|8975,8976
and|8976,8979
nutritional|8980,8991
status|8992,8998
a|8999,9000
goals|9001,9006
of|9007,9009
care|9010,9014
discussion|9015,9025
was|9026,9029
held|9030,9034
with|9035,9039
<EOL>|9040,9041
the|9041,9044
patient|9045,9052
's|9052,9054
HCP|9055,9058
,|9058,9059
_|9060,9061
_|9061,9062
_|9062,9063
and|9064,9067
it|9068,9070
was|9071,9074
decided|9075,9082
to|9083,9085
focus|9086,9091
<EOL>|9092,9093
goals|9093,9098
of|9099,9101
care|9102,9106
of|9107,9109
comfort|9110,9117
and|9118,9121
symptom|9122,9129
management|9130,9140
and|9141,9144
the|9145,9148
patient|9149,9156
<EOL>|9157,9158
was|9158,9161
discharged|9162,9172
home|9173,9177
with|9178,9182
home|9183,9187
hospice|9188,9195
.|9195,9196
<EOL>|9197,9198
<EOL>|9198,9199
(|9199,9200
2|9200,9201
)|9201,9202
Left|9203,9207
thigh|9208,9213
weakness|9214,9222
/|9222,9223
spinous|9223,9230
tenderness|9231,9241
:|9241,9242
She|9243,9246
was|9247,9250
found|9251,9256
to|9257,9259
<EOL>|9260,9261
have|9261,9265
focal|9266,9271
left|9272,9276
thigh|9277,9282
weakness|9283,9291
in|9292,9294
association|9295,9306
with|9307,9311
diffuse|9312,9319
<EOL>|9320,9321
spinous|9321,9328
tenderness|9329,9339
of|9340,9342
unclear|9343,9350
chronicity|9351,9361
in|9362,9364
the|9365,9368
setting|9369,9376
of|9377,9379
<EOL>|9380,9381
preserved|9381,9390
rectal|9391,9397
tone|9398,9402
without|9403,9410
saddle|9411,9417
anesthesia|9418,9428
.|9428,9429
She|9430,9433
was|9434,9437
noted|9438,9443
<EOL>|9444,9445
to|9445,9447
be|9448,9450
incontinent|9451,9462
of|9463,9465
urine|9466,9471
,|9471,9472
but|9473,9476
not|9477,9480
feces|9481,9486
.|9486,9487
Given|9488,9493
underlying|9494,9504
<EOL>|9505,9506
malignancy|9506,9516
,|9516,9517
there|9518,9523
was|9524,9527
concern|9528,9535
for|9536,9539
bony|9540,9544
metastases|9545,9555
or|9556,9558
cord|9559,9563
<EOL>|9564,9565
involvement|9565,9576
,|9576,9577
with|9578,9582
alternative|9583,9594
consideration|9595,9608
given|9609,9614
to|9615,9617
epidural|9618,9626
<EOL>|9627,9628
abscess|9628,9635
,|9635,9636
prompting|9637,9646
transient|9647,9656
initiation|9657,9667
of|9668,9670
empiric|9671,9678
antibiotic|9679,9689
<EOL>|9690,9691
coverage|9691,9699
with|9700,9704
vancomycin|9705,9715
/|9715,9716
cefepim|9716,9723
_|9724,9725
_|9725,9726
_|9726,9727
to|9728,9730
_|9731,9732
_|9732,9733
_|9733,9734
.|9734,9735
Despite|9736,9743
<EOL>|9744,9745
frequent|9745,9753
persuasive|9754,9764
efforts|9765,9772
,|9772,9773
she|9774,9777
declined|9778,9786
multiple|9787,9795
attempts|9796,9804
at|9805,9807
<EOL>|9808,9809
lumbosacral|9809,9820
MRI|9821,9824
,|9824,9825
including|9826,9835
with|9836,9840
lorazepam|9841,9850
premedication|9851,9864
,|9864,9865
citing|9866,9872
<EOL>|9873,9874
claustrophobia|9874,9888
.|9888,9889
Neuro|9890,9895
exam|9896,9900
was|9901,9904
monitored|9905,9914
and|9915,9918
remained|9919,9927
stable|9928,9934
.|9934,9935
<EOL>|9935,9936
<EOL>|9936,9937
(|9937,9938
3|9938,9939
)|9939,9940
Abdominal|9941,9950
pain|9951,9955
:|9955,9956
She|9957,9960
experienced|9961,9972
intermittent|9973,9985
abdominal|9986,9995
pain|9996,10000
<EOL>|10001,10002
and|10002,10005
tenderness|10006,10016
without|10017,10024
peritoneal|10025,10035
signs|10036,10041
,|10041,10042
concerning|10043,10053
for|10054,10057
<EOL>|10058,10059
obstruction|10059,10070
in|10071,10073
the|10074,10077
setting|10078,10085
of|10086,10088
intraabdominal|10089,10103
malignancy|10104,10114
,|10114,10115
<EOL>|10116,10117
particularly|10117,10129
given|10130,10135
episodes|10136,10144
of|10145,10147
emesis|10148,10154
/|10154,10155
hematemesis|10155,10166
as|10167,10169
below|10170,10175
.|10175,10176
<EOL>|10177,10178
While|10178,10183
multiple|10184,10192
KUBs|10193,10197
were|10198,10202
negative|10203,10211
for|10212,10215
obstruction|10216,10227
,|10227,10228
CT|10229,10231
abdomen|10232,10239
<EOL>|10240,10241
was|10241,10244
planned|10245,10252
to|10253,10255
evaluate|10256,10264
for|10265,10268
alternative|10269,10280
sources|10281,10288
of|10289,10291
<EOL>|10292,10293
intraabdominal|10293,10307
pathology|10308,10317
,|10317,10318
but|10319,10322
she|10323,10326
declined|10327,10335
on|10336,10338
multiple|10339,10347
<EOL>|10348,10349
occasions|10349,10358
.|10358,10359
Pain|10360,10364
was|10365,10368
controlled|10369,10379
with|10380,10384
acetaminophen|10385,10398
and|10399,10402
tramadol|10403,10411
<EOL>|10412,10413
as|10413,10415
needed|10416,10422
.|10422,10423
<EOL>|10423,10424
<EOL>|10424,10425
(|10425,10426
4|10426,10427
)|10427,10428
?|10429,10430
Hematemesis|10431,10442
:|10442,10443
She|10444,10447
experienced|10448,10459
a|10460,10461
single|10462,10468
episode|10469,10476
of|10477,10479
small|10480,10485
<EOL>|10486,10487
volume|10487,10493
emesis|10494,10500
,|10500,10501
reportedly|10502,10512
approximately|10513,10526
100cc|10527,10532
,|10532,10533
streaked|10534,10542
with|10543,10547
<EOL>|10548,10549
blood|10549,10554
and|10555,10558
found|10559,10564
to|10565,10567
be|10568,10570
guiac|10571,10576
positive|10577,10585
.|10585,10586
Vital|10587,10592
signs|10593,10598
and|10599,10602
hematocrit|10603,10613
<EOL>|10614,10615
remained|10615,10623
stable|10624,10630
.|10630,10631
IV|10632,10634
pantoprazole|10635,10647
was|10648,10651
initiated|10652,10661
for|10662,10665
<EOL>|10666,10667
gastrointestinal|10667,10683
prophylaxis|10684,10695
,|10695,10696
with|10697,10701
subsequent|10702,10712
discontinuation|10713,10728
of|10729,10731
<EOL>|10732,10733
PPI|10733,10736
given|10737,10742
no|10743,10745
recurrence|10746,10756
and|10757,10760
questionable|10761,10773
if|10774,10776
first|10777,10782
episode|10783,10790
was|10791,10794
<EOL>|10795,10796
true|10796,10800
blood|10801,10806
vs.|10807,10810
red|10811,10814
popsicle|10815,10823
was|10824,10827
eating|10828,10834
at|10835,10837
time|10838,10842
.|10842,10843
<EOL>|10844,10845
Esophagogastroduodenoscopy|10845,10871
was|10872,10875
deferred|10876,10884
in|10885,10887
the|10888,10891
absence|10892,10899
of|10900,10902
<EOL>|10903,10904
recurrent|10904,10913
hematemesis|10914,10925
;|10925,10926
no|10927,10929
prior|10930,10935
EGDs|10936,10940
were|10941,10945
available|10946,10955
in|10956,10958
OMR|10959,10962
.|10962,10963
<EOL>|10964,10965
<EOL>|10965,10966
(|10966,10967
5|10967,10968
)|10968,10969
Altered|10970,10977
mental|10978,10984
status|10985,10991
:|10991,10992
She|10993,10996
was|10997,11000
intermittently|11001,11015
altered|11016,11023
<EOL>|11024,11025
throughout|11025,11035
admission|11036,11045
,|11045,11046
never|11047,11052
oriented|11053,11061
to|11062,11064
more|11065,11069
than|11070,11074
person|11075,11081
and|11082,11085
<EOL>|11086,11087
place|11087,11092
,|11092,11093
with|11094,11098
occasional|11099,11109
difficulty|11110,11120
following|11121,11130
simple|11131,11137
commands|11138,11146
as|11147,11149
<EOL>|11150,11151
compared|11151,11159
to|11160,11162
an|11163,11165
uncertain|11166,11175
baseline|11176,11184
.|11184,11185
Infectious|11186,11196
work|11197,11201
up|11202,11204
,|11204,11205
including|11206,11215
<EOL>|11216,11217
blood|11217,11222
and|11223,11226
urine|11227,11232
cultures|11233,11241
and|11242,11245
CTA|11246,11249
on|11250,11252
admission|11253,11262
with|11263,11267
subsequent|11268,11278
<EOL>|11279,11280
CXRs|11280,11284
,|11284,11285
was|11286,11289
unrevealing|11290,11301
.|11301,11302
Noncontrast|11303,11314
head|11315,11319
CT|11320,11322
was|11323,11326
negative|11327,11335
for|11336,11339
<EOL>|11340,11341
acute|11341,11346
intracranial|11347,11359
process|11360,11367
.|11367,11368
Brain|11369,11374
MRI|11375,11378
for|11379,11382
definitive|11383,11393
exclusion|11394,11403
<EOL>|11404,11405
of|11405,11407
metastases|11408,11418
could|11419,11424
not|11425,11428
be|11429,11431
obtained|11432,11440
due|11441,11444
to|11445,11447
claustrophobia|11448,11462
/|11462,11463
MRI|11463,11466
<EOL>|11467,11468
aversion|11468,11476
as|11477,11479
above|11480,11485
.|11485,11486
ABG|11488,11491
on|11492,11494
_|11495,11496
_|11496,11497
_|11497,11498
without|11499,11506
signs|11507,11512
of|11513,11515
CO2|11516,11519
retention|11520,11529
.|11529,11530
<EOL>|11531,11532
History|11532,11539
of|11540,11542
opiates|11543,11550
making|11551,11557
patient|11558,11565
sleepy|11566,11572
per|11573,11576
HCP|11577,11580
as|11581,11583
possible|11584,11592
<EOL>|11593,11594
contributing|11594,11606
factor|11607,11613
and|11614,11617
therefore|11618,11627
these|11628,11633
were|11634,11638
discontinued|11639,11651
.|11651,11652
<EOL>|11653,11654
Hepatic|11654,11661
encephalopathy|11662,11676
also|11677,11681
on|11682,11684
differential|11685,11697
given|11698,11703
metastatic|11704,11714
<EOL>|11715,11716
lesions|11716,11723
to|11724,11726
liver|11727,11732
and|11733,11736
asterixis|11737,11746
on|11747,11749
exam|11750,11754
.|11754,11755
AMS|11757,11760
could|11761,11766
also|11767,11771
be|11772,11774
_|11775,11776
_|11776,11777
_|11777,11778
<EOL>|11779,11780
to|11780,11782
severe|11783,11789
depression|11790,11800
.|11800,11801
Mental|11802,11808
status|11809,11815
monitored|11816,11825
and|11826,11829
remained|11830,11838
<EOL>|11839,11840
stable|11840,11846
and|11847,11850
patient|11851,11858
at|11859,11861
baseline|11862,11870
per|11871,11874
HCP|11875,11878
on|11879,11881
discharge|11882,11891
.|11891,11892
<EOL>|11892,11893
<EOL>|11893,11894
(|11894,11895
6|11895,11896
)|11896,11897
Shortness|11898,11907
of|11908,11910
breath|11911,11917
:|11917,11918
She|11919,11922
presented|11923,11932
with|11933,11937
acute|11938,11943
onset|11944,11949
<EOL>|11950,11951
shortness|11951,11960
of|11961,11963
breath|11964,11970
without|11971,11978
frank|11979,11984
hypoxia|11985,11992
.|11992,11993
CTA|11994,11997
on|11998,12000
admission|12001,12010
was|12011,12014
<EOL>|12015,12016
negative|12016,12024
for|12025,12028
pulmonary|12029,12038
embolus|12039,12046
,|12046,12047
though|12048,12054
(|12055,12056
subsegmental|12056,12068
clot|12069,12073
could|12074,12079
<EOL>|12080,12081
not|12081,12084
be|12085,12087
excluded|12088,12096
definitively|12097,12109
)|12109,12110
,|12110,12111
pleural|12112,12119
effusion|12120,12128
,|12128,12129
or|12130,12132
focal|12133,12138
<EOL>|12139,12140
infiltrate|12140,12150
.|12150,12151
EKG|12152,12155
and|12156,12159
cardiac|12160,12167
enzymes|12168,12175
were|12176,12180
reassuring|12181,12191
against|12192,12199
<EOL>|12200,12201
acute|12201,12206
coronary|12207,12215
syndrome|12216,12224
.|12224,12225
Low|12227,12230
voltages|12231,12239
on|12240,12242
EKG|12243,12246
were|12247,12251
consistent|12252,12262
<EOL>|12263,12264
with|12264,12268
prior|12269,12274
,|12274,12275
hence|12276,12281
limited|12282,12289
suspicion|12290,12299
for|12300,12303
pericardial|12304,12315
effusion|12316,12324
.|12324,12325
<EOL>|12326,12327
Shortness|12327,12336
of|12337,12339
breath|12340,12346
resolved|12347,12355
over|12356,12360
the|12361,12364
course|12365,12371
of|12372,12374
admission|12375,12384
<EOL>|12385,12386
without|12386,12393
dedicated|12394,12403
treatment|12404,12413
,|12413,12414
with|12415,12419
the|12420,12423
exception|12424,12433
of|12434,12436
nebulizers|12437,12447
<EOL>|12448,12449
and|12449,12452
expectorants|12453,12465
as|12466,12468
needed|12469,12475
.|12475,12476
<EOL>|12476,12477
<EOL>|12477,12478
(|12478,12479
7|12479,12480
)|12480,12481
Leukocytosis|12482,12494
:|12494,12495
White|12496,12501
blood|12502,12507
cell|12508,12512
count|12513,12518
was|12519,12522
elevated|12523,12531
and|12532,12535
peaked|12536,12542
<EOL>|12543,12544
at|12544,12546
20.6|12547,12551
,|12551,12552
consistent|12553,12563
with|12564,12568
recent|12569,12575
baseline|12576,12584
,|12584,12585
likely|12586,12592
reflecting|12593,12603
<EOL>|12604,12605
underlying|12605,12615
malignancy|12616,12626
.|12626,12627
As|12628,12630
noted|12631,12636
above|12637,12642
,|12642,12643
infectious|12644,12654
work|12655,12659
up|12660,12662
<EOL>|12663,12664
including|12664,12673
CTA|12674,12677
,|12677,12678
urine|12679,12684
and|12685,12688
blood|12689,12694
cultures|12695,12703
,|12703,12704
and|12705,12708
CXRs|12709,12713
,|12713,12714
was|12715,12718
<EOL>|12719,12720
unrevealing|12720,12731
.|12731,12732
She|12733,12736
remained|12737,12745
afebrile|12746,12754
,|12754,12755
with|12756,12760
the|12761,12764
exception|12765,12774
of|12775,12777
<EOL>|12778,12779
isolated|12779,12787
transient|12788,12797
fever|12798,12803
to|12804,12806
100|12807,12810
,|12810,12811
with|12812,12816
stable|12817,12823
vital|12824,12829
signs|12830,12835
.|12835,12836
<EOL>|12837,12838
<EOL>|12838,12839
(|12839,12840
8|12840,12841
)|12842,12843
Liver|12843,12848
function|12849,12857
test|12858,12862
abnormalities|12863,12876
:|12876,12877
AST|12878,12881
remained|12882,12890
elevated|12891,12899
_|12900,12901
_|12901,12902
_|12902,12903
<EOL>|12904,12905
to|12905,12907
_|12908,12909
_|12909,12910
_|12910,12911
,|12911,12912
alkaline|12913,12921
phosphatase|12922,12933
260s|12934,12938
to|12939,12941
380s|12942,12946
,|12946,12947
and|12948,12951
total|12952,12957
bilirubin|12958,12967
<EOL>|12968,12969
2.1|12969,12972
to|12973,12975
2.6|12976,12979
,|12979,12980
likely|12981,12987
due|12988,12991
to|12992,12994
hepatic|12995,13002
infiltration|13003,13015
of|13016,13018
malignancy|13019,13029
.|13029,13030
<EOL>|13031,13032
Right|13032,13037
upper|13038,13043
quadrant|13044,13052
ultrasound|13053,13063
was|13064,13067
negative|13068,13076
for|13077,13080
cholecystitis|13081,13094
<EOL>|13095,13096
or|13096,13098
obstructive|13099,13110
process|13111,13118
.|13118,13119
The|13120,13123
possibility|13124,13135
of|13136,13138
superimposed|13139,13151
<EOL>|13152,13153
intraabdominal|13153,13167
process|13168,13175
,|13175,13176
such|13177,13181
as|13182,13184
infection|13185,13194
,|13194,13195
could|13196,13201
not|13202,13205
be|13206,13208
excluded|13209,13217
<EOL>|13218,13219
in|13219,13221
the|13222,13225
setting|13226,13233
of|13234,13236
abdominal|13237,13246
pain|13247,13251
with|13252,13256
emesis|13257,13263
as|13264,13266
above|13267,13272
,|13272,13273
but|13274,13277
she|13278,13281
<EOL>|13282,13283
declined|13283,13291
CT|13292,13294
for|13295,13298
further|13299,13306
evaluation|13307,13317
.|13317,13318
<EOL>|13318,13319
<EOL>|13319,13320
(|13320,13321
9|13321,13322
)|13322,13323
Elevated|13324,13332
lactate|13333,13340
:|13340,13341
Lactate|13342,13349
was|13350,13353
found|13354,13359
to|13360,13362
be|13363,13365
2.7|13366,13369
-|13369,13370
3.8|13370,13373
throughout|13374,13384
<EOL>|13385,13386
admission|13386,13395
despite|13396,13403
copious|13404,13411
IV|13412,13414
fluids|13415,13421
,|13421,13422
likely|13423,13429
reflecting|13430,13440
<EOL>|13441,13442
compromised|13442,13453
hepatic|13454,13461
clearance|13462,13471
in|13472,13474
the|13475,13478
setting|13479,13486
of|13487,13489
malignant|13490,13499
<EOL>|13500,13501
infiltration|13501,13513
.|13513,13514
<EOL>|13515,13516
<EOL>|13516,13517
(|13517,13518
10|13518,13520
)|13520,13521
Sinus|13522,13527
tachycardia|13528,13539
:|13539,13540
She|13541,13544
remained|13545,13553
persistently|13554,13566
tachycardic|13567,13578
<EOL>|13579,13580
100s|13580,13584
to|13585,13587
115s|13588,13592
throughout|13593,13603
admission|13604,13613
in|13614,13616
the|13617,13620
setting|13621,13628
of|13629,13631
poor|13632,13636
PO|13637,13639
<EOL>|13640,13641
intake|13641,13647
,|13647,13648
but|13649,13652
incompletely|13653,13665
responsive|13666,13676
to|13677,13679
copious|13680,13687
IV|13688,13690
fluids|13691,13697
.|13697,13698
<EOL>|13699,13700
Tachycardia|13700,13711
has|13712,13715
been|13716,13720
present|13721,13728
since|13729,13734
at|13735,13737
least|13738,13743
_|13744,13745
_|13745,13746
_|13746,13747
.|13747,13748
Despite|13749,13756
<EOL>|13757,13758
concurrent|13758,13768
leukocytosis|13769,13781
and|13782,13785
elevated|13786,13794
lactate|13795,13802
,|13802,13803
there|13804,13809
was|13810,13813
no|13814,13816
clear|13817,13822
<EOL>|13823,13824
infectious|13824,13834
source|13835,13841
,|13841,13842
hence|13843,13848
low|13849,13852
suspicion|13853,13862
for|13863,13866
sepsis|13867,13873
.|13873,13874
Subsegmental|13875,13887
<EOL>|13888,13889
pulmonary|13889,13898
embolus|13899,13906
could|13907,13912
not|13913,13916
be|13917,13919
excluded|13920,13928
on|13929,13931
the|13932,13935
basis|13936,13941
of|13942,13944
<EOL>|13945,13946
admission|13946,13955
CTA|13956,13959
,|13959,13960
but|13961,13964
shortness|13965,13974
of|13975,13977
breath|13978,13984
was|13985,13988
short|13989,13994
lived|13995,14000
,|14000,14001
and|14002,14005
she|14006,14009
<EOL>|14010,14011
was|14011,14014
never|14015,14020
hypoxic|14021,14028
.|14028,14029
Hematocrit|14030,14040
remained|14041,14049
stable|14050,14056
without|14057,14064
signs|14065,14070
of|14071,14073
<EOL>|14074,14075
active|14075,14081
bleeding|14082,14090
,|14090,14091
with|14092,14096
the|14097,14100
exception|14101,14110
of|14111,14113
transient|14114,14123
hematemesis|14124,14135
as|14136,14138
<EOL>|14139,14140
above|14140,14145
.|14145,14146
<EOL>|14146,14147
<EOL>|14147,14148
(|14148,14149
11|14149,14151
)|14151,14152
Depression|14153,14163
:|14163,14164
She|14165,14168
appeared|14169,14177
depressed|14178,14187
with|14188,14192
flat|14193,14197
affect|14198,14204
and|14205,14208
<EOL>|14209,14210
seeming|14210,14217
anhedonia|14218,14227
throughout|14228,14238
admission|14239,14248
,|14248,14249
with|14250,14254
underlying|14255,14265
<EOL>|14266,14267
depression|14267,14277
likely|14278,14284
affecting|14285,14294
motivation|14295,14305
to|14306,14308
seek|14309,14313
diagnosis|14314,14323
and|14324,14327
<EOL>|14328,14329
treatment|14329,14338
of|14339,14341
known|14342,14347
malignancy|14348,14358
.|14358,14359
She|14360,14363
denied|14364,14370
active|14371,14377
suicidal|14378,14386
<EOL>|14387,14388
ideation|14388,14396
and|14397,14400
frequently|14401,14411
declined|14412,14420
home|14421,14425
sertraline|14426,14436
,|14436,14437
particularly|14438,14450
<EOL>|14451,14452
prior|14452,14457
to|14458,14460
liver|14461,14466
biopsy|14467,14473
,|14473,14474
believing|14475,14484
that|14485,14489
it|14490,14492
was|14493,14496
supposed|14497,14505
to|14506,14508
be|14509,14511
held|14512,14516
<EOL>|14517,14518
preprocedurally|14518,14533
despite|14534,14541
explanation|14542,14553
to|14554,14556
the|14557,14560
contrary|14561,14569
.|14569,14570
She|14571,14574
was|14575,14578
<EOL>|14579,14580
seen|14580,14584
by|14585,14587
social|14588,14594
work|14595,14599
throughout|14600,14610
admission|14611,14620
.|14620,14621
<EOL>|14621,14622
<EOL>|14622,14623
(|14623,14624
12|14624,14626
)|14626,14627
Normocytic|14628,14638
anemia|14639,14645
:|14645,14646
Hematocrit|14647,14657
remained|14658,14666
stable|14667,14673
and|14674,14677
<EOL>|14678,14679
consistent|14679,14689
with|14690,14694
recent|14695,14701
baseline|14702,14710
at|14711,14713
27|14714,14716
to|14717,14719
33|14720,14722
throughout|14723,14733
<EOL>|14734,14735
admission|14735,14744
,|14744,14745
seemingly|14746,14755
due|14756,14759
to|14760,14762
anemia|14763,14769
of|14770,14772
chronic|14773,14780
disease|14781,14788
on|14789,14791
the|14792,14795
<EOL>|14796,14797
basis|14797,14802
of|14803,14805
preadmission|14806,14818
labs|14819,14823
.|14823,14824
Vital|14825,14830
signs|14831,14836
remained|14837,14845
stable|14846,14852
,|14852,14853
with|14854,14858
<EOL>|14859,14860
the|14860,14863
exception|14864,14873
of|14874,14876
persistent|14877,14887
tachycardia|14888,14899
,|14899,14900
without|14901,14908
signs|14909,14914
of|14915,14917
active|14918,14924
<EOL>|14925,14926
bleeding|14926,14934
apart|14935,14940
from|14941,14945
isolated|14946,14954
blood|14955,14960
streaked|14961,14969
emesis|14970,14976
as|14977,14979
above|14980,14985
.|14985,14986
<EOL>|14986,14987
<EOL>|14987,14988
(|14988,14989
13|14989,14991
)|14991,14992
Coagulopathy|14993,15005
:|15005,15006
INR|15007,15010
of|15011,15013
1.2|15014,15017
to|15018,15020
1.8|15021,15024
was|15025,15028
felt|15029,15033
to|15034,15036
reflect|15037,15044
<EOL>|15045,15046
synthetic|15046,15055
dysfunction|15056,15067
in|15068,15070
the|15071,15074
setting|15075,15082
of|15083,15085
hepatic|15086,15093
infiltration|15094,15106
of|15107,15109
<EOL>|15110,15111
malignancy|15111,15121
,|15121,15122
as|15123,15125
well|15126,15130
as|15131,15133
poor|15134,15138
oral|15139,15143
intake|15144,15150
.|15150,15151
There|15152,15157
were|15158,15162
no|15163,15165
signs|15166,15171
of|15172,15174
<EOL>|15175,15176
active|15176,15182
bleeding|15183,15191
,|15191,15192
with|15193,15197
the|15198,15201
exception|15202,15211
of|15212,15214
transient|15215,15224
hematemesis|15225,15236
as|15237,15239
<EOL>|15240,15241
above|15241,15246
.|15246,15247
<EOL>|15247,15248
<EOL>|15248,15249
Transitional|15249,15261
Issues|15262,15268
:|15268,15269
<EOL>|15269,15270
-|15270,15271
Patient|15271,15278
discharge|15279,15288
home|15289,15293
with|15294,15298
home|15299,15303
hospice|15304,15311
<EOL>|15311,15312
<EOL>|15313,15314
Medications|15314,15325
on|15326,15328
Admission|15329,15338
:|15338,15339
<EOL>|15339,15340
The|15340,15343
Preadmission|15344,15356
Medication|15357,15367
list|15368,15372
may|15373,15376
be|15377,15379
inaccurate|15380,15390
and|15391,15394
requires|15395,15403
<EOL>|15404,15405
futher|15405,15411
investigation|15412,15425
.|15425,15426
<EOL>|15426,15427
1.|15427,15429
Albuterol|15430,15439
Inhaler|15440,15447
_|15448,15449
_|15449,15450
_|15450,15451
PUFF|15452,15456
IH|15457,15459
Q6H|15460,15463
:|15463,15464
PRN|15464,15467
SOB|15468,15471
<EOL>|15472,15473
2.|15473,15475
BuPROPion|15476,15485
150|15486,15489
mg|15490,15492
PO|15493,15495
DAILY|15496,15501
<EOL>|15502,15503
3.|15503,15505
Gabapentin|15506,15516
300|15517,15520
mg|15521,15523
PO|15524,15526
HS|15527,15529
<EOL>|15530,15531
4.|15531,15533
Sertraline|15534,15544
200|15545,15548
mg|15549,15551
PO|15552,15554
DAILY|15555,15560
<EOL>|15561,15562
5.|15562,15564
traZODONE|15565,15574
100|15575,15578
mg|15579,15581
PO|15582,15584
HS|15585,15587
:|15587,15588
PRN|15588,15591
sleep|15592,15597
<EOL>|15598,15599
6.|15599,15601
Ondansetron|15602,15613
4|15614,15615
mg|15616,15618
PO|15619,15621
Q8H|15622,15625
:|15625,15626
PRN|15626,15629
nausea|15630,15636
<EOL>|15637,15638
7.|15638,15640
Bisacodyl|15641,15650
10|15651,15653
mg|15654,15656
PO|15657,15659
/|15659,15660
PR|15660,15662
DAILY|15663,15668
:|15668,15669
PRN|15669,15672
constipation|15673,15685
<EOL>|15686,15687
8.|15687,15689
OxycoDONE|15690,15699
(|15700,15701
Immediate|15701,15710
Release|15711,15718
)|15718,15719
5|15721,15722
mg|15723,15725
PO|15726,15728
Q6H|15729,15732
:|15732,15733
PRN|15733,15736
pain|15737,15741
<EOL>|15742,15743
please|15743,15749
hold|15750,15754
for|15755,15758
sedation|15759,15767
,|15767,15768
RR|15769,15771
<|15771,15772
10|15772,15774
<EOL>|15775,15776
9.|15776,15778
Enoxaparin|15779,15789
Sodium|15790,15796
40|15797,15799
mg|15800,15802
SC|15803,15805
DAILY|15806,15811
<EOL>|15812,15813
<EOL>|15813,15814
<EOL>|15815,15816
Discharge|15816,15825
Medications|15826,15837
:|15837,15838
<EOL>|15838,15839
1.|15839,15841
BuPROPion|15842,15851
150|15852,15855
mg|15856,15858
PO|15859,15861
DAILY|15862,15867
<EOL>|15868,15869
2.|15869,15871
Ondansetron|15872,15883
4|15884,15885
mg|15886,15888
PO|15889,15891
Q8H|15892,15895
:|15895,15896
PRN|15896,15899
nausea|15900,15906
<EOL>|15907,15908
3.|15908,15910
TraMADOL|15911,15919
(|15920,15921
Ultram|15921,15927
)|15927,15928
50|15929,15931
mg|15932,15934
PO|15935,15937
Q4H|15938,15941
:|15941,15942
PRN|15942,15945
pain|15946,15950
<EOL>|15951,15952
RX|15952,15954
*|15955,15956
tramadol|15956,15964
50|15965,15967
mg|15968,15970
1|15971,15972
tablet|15973,15979
(|15979,15980
s|15980,15981
)|15981,15982
by|15983,15985
mouth|15986,15991
every|15992,15997
four|15998,16002
(|16003,16004
4|16004,16005
)|16005,16006
hours|16007,16012
<EOL>|16013,16014
Disp|16014,16018
#|16019,16020
*|16020,16021
60|16021,16023
Tablet|16024,16030
Refills|16031,16038
:|16038,16039
*|16039,16040
0|16040,16041
<EOL>|16041,16042
4.|16042,16044
Senna|16045,16050
1|16051,16052
TAB|16053,16056
PO|16057,16059
BID|16060,16063
:|16063,16064
PRN|16064,16067
constipation|16068,16080
<EOL>|16081,16082
RX|16082,16084
*|16085,16086
sennosides|16086,16096
[|16097,16098
_|16098,16099
_|16099,16100
_|16100,16101
]|16101,16102
8.6|16103,16106
mg|16107,16109
1|16110,16111
tablet|16112,16118
by|16119,16121
mouth|16122,16127
twice|16128,16133
a|16134,16135
<EOL>|16136,16137
day|16137,16140
Disp|16141,16145
#|16146,16147
*|16147,16148
60|16148,16150
Tablet|16151,16157
Refills|16158,16165
:|16165,16166
*|16166,16167
0|16167,16168
<EOL>|16168,16169
5.|16169,16171
Omeprazole|16172,16182
20|16183,16185
mg|16186,16188
PO|16189,16191
DAILY|16192,16197
<EOL>|16198,16199
RX|16199,16201
*|16202,16203
omeprazole|16203,16213
20|16214,16216
mg|16217,16219
1|16220,16221
capsule|16222,16229
,|16229,16230
delayed|16230,16237
_|16238,16239
_|16239,16240
_|16240,16241
by|16242,16244
<EOL>|16245,16246
mouth|16246,16251
Daily|16252,16257
Disp|16258,16262
#|16263,16264
*|16264,16265
30|16265,16267
Capsule|16268,16275
Refills|16276,16283
:|16283,16284
*|16284,16285
0|16285,16286
<EOL>|16286,16287
6.|16287,16289
Hospital|16290,16298
Bed|16299,16302
<EOL>|16302,16303
Bariatric|16303,16312
Hospital|16313,16321
Bed|16322,16325
and|16326,16329
<EOL>|16329,16330
Therapeutic|16330,16341
Mattress|16342,16350
:|16350,16351
BariMaxxII|16352,16362
<EOL>|16362,16363
<EOL>|16363,16364
7.|16364,16366
Hospice|16367,16374
Order|16375,16380
<EOL>|16380,16381
Please|16381,16387
Screen|16388,16394
and|16395,16398
Admit|16399,16404
to|16405,16407
Hospice|16408,16415
.|16415,16416
<EOL>|16416,16417
8.|16417,16419
Bisacodyl|16420,16429
10|16430,16432
mg|16433,16435
PO|16436,16438
/|16438,16439
PR|16439,16441
DAILY|16442,16447
:|16447,16448
PRN|16448,16451
constipation|16452,16464
<EOL>|16465,16466
9.|16466,16468
Docusate|16469,16477
Sodium|16478,16484
100|16485,16488
mg|16489,16491
PO|16492,16494
BID|16495,16498
<EOL>|16499,16500
10.|16500,16503
Sertraline|16504,16514
200|16515,16518
mg|16519,16521
PO|16522,16524
DAILY|16525,16530
<EOL>|16531,16532
11.|16532,16535
traZODONE|16536,16545
100|16546,16549
mg|16550,16552
PO|16553,16555
HS|16556,16558
:|16558,16559
PRN|16559,16562
sleep|16563,16568
<EOL>|16569,16570
12.|16570,16573
Polyethylene|16574,16586
Glycol|16587,16593
17|16594,16596
g|16597,16598
PO|16599,16601
DAILY|16602,16607
:|16607,16608
PRN|16608,16611
constipation|16612,16624
<EOL>|16625,16626
<EOL>|16626,16627
<EOL>|16628,16629
Discharge|16629,16638
Disposition|16639,16650
:|16650,16651
<EOL>|16651,16652
Home|16652,16656
With|16657,16661
Service|16662,16669
<EOL>|16669,16670
<EOL>|16671,16672
Facility|16672,16680
:|16680,16681
<EOL>|16681,16682
_|16682,16683
_|16683,16684
_|16684,16685
<EOL>|16685,16686
<EOL>|16687,16688
Discharge|16688,16697
Diagnosis|16698,16707
:|16707,16708
<EOL>|16708,16709
Primary|16709,16716
:|16716,16717
<EOL>|16717,16718
Metastatic|16718,16728
colon|16729,16734
adenocarcinoma|16735,16749
<EOL>|16749,16750
<EOL>|16750,16751
<EOL>|16752,16753
Mental|16774,16780
Status|16781,16787
:|16787,16788
Confused|16789,16797
-|16798,16799
sometimes|16800,16809
.|16809,16810
<EOL>|16810,16811
Level|16811,16816
of|16817,16819
Consciousness|16820,16833
:|16833,16834
Alert|16835,16840
and|16841,16844
interactive|16845,16856
.|16856,16857
<EOL>|16857,16858
Activity|16858,16866
Status|16867,16873
:|16873,16874
Bedbound|16875,16883
.|16883,16884
<EOL>|16884,16885
<EOL>|16885,16886
<EOL>|16887,16888
Dear|16912,16916
Ms.|16917,16920
_|16921,16922
_|16922,16923
_|16923,16924
,|16924,16925
<EOL>|16925,16926
It|16926,16928
was|16929,16932
a|16933,16934
pleasure|16935,16943
taking|16944,16950
part|16951,16955
in|16956,16958
your|16959,16963
care|16964,16968
during|16969,16975
your|16976,16980
admission|16981,16990
<EOL>|16991,16992
to|16992,16994
_|16995,16996
_|16996,16997
_|16997,16998
.|16998,16999
As|17000,17002
you|17003,17006
know|17007,17011
,|17011,17012
you|17013,17016
were|17017,17021
<EOL>|17022,17023
admitted|17023,17031
for|17032,17035
shortness|17036,17045
of|17046,17048
breath|17049,17055
,|17055,17056
likely|17057,17063
due|17064,17067
to|17068,17070
your|17071,17075
underlying|17076,17086
<EOL>|17087,17088
cancer|17088,17094
,|17094,17095
and|17096,17099
there|17100,17105
was|17106,17109
no|17110,17112
evidence|17113,17121
of|17122,17124
pneumonia|17125,17134
or|17135,17137
blood|17138,17143
clot|17144,17148
in|17149,17151
<EOL>|17152,17153
the|17153,17156
blood|17157,17162
vessels|17163,17170
of|17171,17173
your|17174,17178
lungs|17179,17184
.|17184,17185
Your|17186,17190
shortness|17191,17200
of|17201,17203
breath|17204,17210
<EOL>|17211,17212
resolved|17212,17220
,|17220,17221
but|17222,17225
you|17226,17229
were|17230,17234
found|17235,17240
to|17241,17243
have|17244,17248
weakness|17249,17257
in|17258,17260
your|17261,17265
left|17266,17270
thigh|17271,17276
<EOL>|17277,17278
and|17278,17281
abdominal|17282,17291
pain|17292,17296
.|17296,17297
You|17298,17301
declined|17302,17310
imaging|17311,17318
studies|17319,17326
for|17327,17330
further|17331,17338
<EOL>|17339,17340
investigation|17340,17353
of|17354,17356
these|17357,17362
findings|17363,17371
.|17371,17372
You|17373,17376
underwent|17377,17386
biopsy|17387,17393
of|17394,17396
your|17397,17401
<EOL>|17402,17403
liver|17403,17408
that|17409,17413
revealed|17414,17422
that|17423,17427
the|17428,17431
cancer|17432,17438
known|17439,17444
to|17445,17447
affect|17448,17454
your|17455,17459
liver|17460,17465
<EOL>|17466,17467
and|17467,17470
lungs|17471,17476
originated|17477,17487
in|17488,17490
your|17491,17495
colon|17496,17501
(|17502,17503
large|17503,17508
bowel|17509,17514
)|17514,17515
.|17515,17516
You|17517,17520
were|17521,17525
<EOL>|17526,17527
transferred|17527,17538
to|17539,17541
the|17542,17545
oncology|17546,17554
service|17555,17562
,|17562,17563
but|17564,17567
unfortunately|17568,17581
<EOL>|17582,17583
chemotherapy|17583,17595
would|17596,17601
do|17602,17604
more|17605,17609
harm|17610,17614
for|17615,17618
you|17619,17622
than|17623,17627
good|17628,17632
.|17632,17633
After|17635,17640
a|17641,17642
long|17643,17647
<EOL>|17648,17649
discussion|17649,17659
with|17660,17664
you|17665,17668
and|17669,17672
your|17673,17677
health|17678,17684
care|17685,17689
proxy|17690,17695
,|17695,17696
it|17697,17699
was|17700,17703
decided|17704,17711
<EOL>|17712,17713
that|17713,17717
you|17718,17721
will|17722,17726
go|17727,17729
home|17730,17734
to|17735,17737
be|17738,17740
with|17741,17745
your|17746,17750
family|17751,17757
and|17758,17761
loved|17762,17767
ones|17768,17772
.|17772,17773
We|17775,17777
<EOL>|17778,17779
will|17779,17783
also|17784,17788
set|17789,17792
up|17793,17795
hospice|17796,17803
services|17804,17812
for|17813,17816
you|17817,17820
so|17821,17823
that|17824,17828
they|17829,17833
can|17834,17837
help|17838,17842
<EOL>|17843,17844
with|17844,17848
any|17849,17852
issues|17853,17859
that|17860,17864
arise|17865,17870
while|17871,17876
you|17877,17880
are|17881,17884
at|17885,17887
home|17888,17892
.|17892,17893
<EOL>|17895,17896
<EOL>|17897,17898
Followup|17898,17906
Instructions|17907,17919
:|17919,17920
<EOL>|17920,17921
_|17921,17922
_|17922,17923
_|17923,17924
<EOL>|17924,17925

