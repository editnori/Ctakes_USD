CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|false|false||Drugsnull|Drugs - dental services|Procedure|false|false||Drugsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Abdomen distended|Finding|false|false||Abdominal distentionnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Distention|Finding|false|false||distention
null|Pathological Dilatation|Finding|false|false||distentionnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Paracentesis|Procedure|false|false||Paracentesisnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Very|Modifier|false|false||verynull|Nitroglycerin/Sodium Citrate/Ethanol Solution|Drug|false|false||nice
null|Nitroglycerin/Sodium Citrate/Ethanol Solution|Drug|false|false||nicenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Alcohol abuse|Disorder|false|false||ETOH abusenull|ethanol|Drug|false|false||ETOH
null|ethanol|Drug|false|false||ETOHnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Constipation|Finding|false|false||constipationnull|Abdomen distended|Finding|false|false||abdominal distentionnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Distention|Finding|false|false||distention
null|Pathological Dilatation|Finding|false|false||distentionnull|10 days|Time|false|false||10 daysnull|day|Time|false|false||daysnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Eyeglasses|Device|false|false||glassesnull|Wine|Drug|false|false||winenull|Night time|Time|false|false||nightnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Binge Drinking|Finding|false|false||binge drinkingnull|Binge eating behavior|Finding|false|false||bingenull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|1 Month|Time|false|false||1 monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Abdomen distended|Finding|false|false||abdominal distensionnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Progressive|Finding|false|false||progressivenull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Solid Dose Form|Drug|false|false||solid
null|solid substance|Drug|false|false||solidnull|Solid|Modifier|false|false||solidnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|Dyspnea|Finding|false|false||SOBnull|Dyspnea on exertion|Finding|false|false||DOEnull|Department of Energy|Subject|false|false||DOEnull|Adult female goat|Entity|false|false||DOEnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Physiologic tolerance|Finding|false|false||tolerance
null|Mental tolerance|Finding|false|false||tolerance
null|Immune Tolerance|Finding|false|false||tolerance
null|Drug Tolerance|Finding|false|false||tolerancenull|Tolerance|Modifier|false|false||tolerancenull|Recent|Time|false|false||recentnull|travel|Finding|false|false||travelnull|travel charge|Procedure|false|false||travelnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|true|false||NSAIDs
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|true|false||NSAIDsnull|Tylenol|Drug|true|false||Tylenol
null|Tylenol|Drug|true|false||Tylenolnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|null|Drug|true|false||medications othernull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Infrequent|Time|false|false||occasionalnull|Menstruation|Finding|false|false||periodsnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Fatty Liver|Disorder|false|false||fatty liver
null|Steatohepatitis|Disorder|false|false||fatty livernull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Hepatic|Anatomy|false|false||portalnull|Flow|Phenomenon|false|false||flownull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Valium|Drug|false|false||valium
null|Valium|Drug|false|false||valiumnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false||IVFnull|SCN5A wt Allele|Finding|false|false||IVF
null|SCN5A gene|Finding|false|false||IVFnull|Assisted Reproductive Technologies|Procedure|false|false||IVF
null|Fertilization in Vitro|Procedure|false|false||IVFnull|Structure of interventricular foramen|Anatomy|false|false||IVFnull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Alcohol abuse|Disorder|false|false||Alcohol abusenull|Alcohols|Drug|false|false||Alcohol
null|Alcohols|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||Alcoholnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Chronic back pain|Finding|false|false||Chronic back painnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Malignant neoplasm of breast|Disorder|false|true||Breast Canull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||Breastnull|Breast problem|Finding|false|false||Breastnull|Procedures on breast|Procedure|false|false||Breastnull|Breast|Anatomy|false|false||Breastnull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|ibudilast|Drug|true|false||IBD
null|ibudilast|Drug|true|false||IBDnull|Inflammatory Bowel Diseases|Disorder|true|false||IBD
null|Irritable Bowel Syndrome|Disorder|true|false||IBDnull|ACAD8 wt Allele|Finding|true|false||IBDnull|Liver Failure|Disorder|true|false||liver failurenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Failure (biologic function)|Finding|true|false||failure
null|Failure|Finding|true|false||failure
null|Personal failure|Finding|true|false||failurenull|Numerous|LabModifier|false|false||Multiplenull|Relative (related person)|Subject|false|false||relativesnull|Alcoholic Intoxication, Chronic|Disorder|false|false||alcoholismnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|Pleasant|Finding|false|false||pleasantnull|Appropriate|Modifier|false|false||appropriatenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|HEENT|Anatomy|false|false||HEENTnull|Facial wasting|Disorder|true|false||temporal wastingnull|Temporal wasting|Finding|true|false||temporal wastingnull|Temporal - Temporal Qualifier|Time|false|false||temporalnull|Temporal Anatomic Qualifier|Modifier|false|false||temporalnull|Wasting|Disorder|true|false||wastingnull|Cachexia|Finding|true|false||wastingnull|Jugular venous engorgement|Finding|true|false||JVDnull|Neck>Neck veins|Anatomy|false|false||neck veins
null|Structure of vein of neck|Anatomy|false|false||neck veinsnull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Fill|Event|false|false||fillnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|MAS1L gene|Finding|true|false||MRGnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|cetrimonium bromide|Drug|false|false||CTABnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Dilated|Finding|false|false||Distendednull|Distended|Modifier|false|false||Distendednull|Tights|Device|false|false||tightnull|Tightness sensation quality|Modifier|false|false||tightnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Flatulence|Finding|false|false||flatulencenull|Limb structure|Anatomy|false|false||LIMBSnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Lewis Blood-Group System|Finding|false|false||LEsnull|Inferior esophageal sphincter structure|Anatomy|false|false||LEsnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Asterixis|Finding|true|false||asterixisnull|Very mild|Finding|true|false||very mildnull|Very|Modifier|false|false||verynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||generalnull|General medical service|Procedure|false|false||generalnull|Generalized|Modifier|false|false||generalnull|Tremor|Finding|false|false||tremornull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Gamma-glutamyl transferase|Drug|false|false||GGT
null|Gamma-glutamyl transferase|Drug|false|false||GGTnull|GGT2P gene|Finding|false|false||GGT
null|GGT1 gene|Finding|false|false||GGTnull|Gamma glutamyl transferase measurement|Procedure|false|false||GGTnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Greater|LabModifier|false|false||GREATERnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|T4 free measurement|Procedure|false|false||Free T4null|Free of (attribute)|Finding|false|false||Freenull|Empty (qualifier)|Modifier|false|false||Freenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Hepatitis B Surface Antigens|Drug|false|false||HBsAg
null|Hepatitis B Surface Antigens|Drug|false|false||HBsAg
null|Hepatitis B Surface Antigens|Drug|false|false||HBsAg
null|Hepatitis B Antigen Vaccine|Drug|false|false||HBsAg
null|Hepatitis B Antigen Vaccine|Drug|false|false||HBsAg
null|Hepatitis B Antigen Vaccine|Drug|false|false||HBsAgnull|Hepatitis B surface antigen measurement|Procedure|false|false||HBsAgnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Hepatitis B Virus Surface Antibody|Drug|false|false||HBsAb
null|Hepatitis B Virus Surface Antibody|Drug|false|false||HBsAbnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Antibody to hepatitis B core antigen|Drug|false|false||HBcAb
null|Antibody to hepatitis B core antigen|Drug|false|false||HBcAb
null|Antibody to hepatitis B core antigen|Drug|false|false||HBcAbnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Hepatitis A|Disorder|false|false||HAVnull|AB(S) hearing assessment list|Device|false|false||Abnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Immunoglobulin M|Drug|false|false||IgM
null|Immunoglobulin M|Drug|false|false||IgMnull|CD40LG wt Allele|Finding|false|false||IgMnull|Immunoglobulin M measurement|Procedure|false|false||IgMnull|Hepatitis A|Disorder|false|false||HAVnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Recombinant Human Chorionic Gonadotropin|Drug|false|false||HCG
null|human chorionic gonadotropin|Drug|false|false||HCG
null|human chorionic gonadotropin|Drug|false|false||HCG
null|human chorionic gonadotropin|Drug|false|false||HCG
null|Recombinant Human Chorionic Gonadotropin|Drug|false|false||HCG
null|Recombinant Human Chorionic Gonadotropin|Drug|false|false||HCGnull|HYPERTRICHOSIS, CONGENITAL GENERALIZED, 2|Disorder|false|false||HCGnull|CGA wt Allele|Finding|false|false||HCG
null|HTC2 gene|Finding|false|false||HCG
null|CGA gene|Finding|false|false||HCG
null|CGB5 gene|Finding|false|false||HCGnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Against Medical Advice|Finding|false|false||AMAnull|cytarabine/melphalan|Procedure|false|false||AMAnull|American Medical Association|Entity|false|false||AMAnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Smooth|Modifier|false|false||Smoothnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|AB(S) hearing assessment list|Device|true|false||Abnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Hold - dosing instruction fragment|Finding|false|false||HOLD
null|hold - Data Operation|Finding|false|false||HOLDnull|Hold (action)|Event|false|false||HOLDnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Hold - dosing instruction fragment|Finding|false|false||HOLD
null|hold - Data Operation|Finding|false|false||HOLDnull|Hold (action)|Event|false|false||HOLDnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|AB(S) hearing assessment list|Device|false|false||Abnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Ceruloplasmin|Drug|false|false||CERULOPLASMIN
null|Ceruloplasmin|Drug|false|false||CERULOPLASMIN
null|CP protein, human|Drug|false|false||CERULOPLASMIN
null|CP protein, human|Drug|false|false||CERULOPLASMINnull|ferroxidase activity|Finding|false|false||CERULOPLASMIN
null|CP gene|Finding|false|false||CERULOPLASMINnull|Ceruloplasmin measurement|Procedure|false|false||CERULOPLASMINnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|alpha 1-antitrypsin|Drug|false|false||ALPHA-1-ANTITRYPSIN
null|SERPINA1 protein, human|Drug|false|false||ALPHA-1-ANTITRYPSIN
null|SERPINA1 protein, human|Drug|false|false||ALPHA-1-ANTITRYPSIN
null|alpha 1-antitrypsin|Drug|false|false||ALPHA-1-ANTITRYPSIN
null|alpha 1-antitrypsin|Drug|false|false||ALPHA-1-ANTITRYPSINnull|SERPINA1 gene|Finding|false|false||ALPHA-1-ANTITRYPSINnull|Alpha-1-antitrypsin measurement|Procedure|false|false||ALPHA-1-ANTITRYPSINnull|Alpha-1|Drug|false|false||ALPHA-1null|ALPHA (substance)|Drug|false|false||ALPHA
null|ALPHA (substance)|Drug|false|false||ALPHAnull|Greek letter alpha (qualifier value)|Finding|false|false||ALPHAnull|Alpha Value|Modifier|false|false||ALPHAnull|SERPINA5 protein, human|Drug|false|false||ANTITRYPSIN
null|SERPINA5 protein, human|Drug|false|false||ANTITRYPSINnull|SERPINA1 gene|Finding|false|false||ANTITRYPSINnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|null|Attribute|false|false||US abdnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Echogenic|Finding|false|false||echogenicnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Fatty infiltration|Finding|false|false||fatty infiltrationnull|Infiltration Route of Administration|Finding|false|false||infiltration
null|Infiltration|Finding|false|false||infiltration
null|Spread by direct extension|Finding|false|false||infiltrationnull|Infiltration (procedure)|Procedure|false|false||infiltrationnull|Manufactured form|Device|false|false||formsnull|Qualitative form|Modifier|false|false||formsnull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|More|LabModifier|false|false||morenull|Advanced phase|Modifier|false|false||advancednull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Fibrosis|Finding|false|false||fibrosisnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|anatomical layer|Anatomy|false|false||Layeringnull|Physiological sludge|Finding|false|false||sludgenull|Environmental sludge|Phenomenon|false|false||sludgenull|examination of gallbladder|Procedure|false|false||gallbladdernull|Gallbladder (MMHCC)|Anatomy|false|false||gallbladder
null|Gallbladder|Anatomy|false|false||gallbladder
null|Abdomen>Gallbladder|Anatomy|false|false||gallbladdernull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|examination of gallbladder|Procedure|false|false||gallbladdernull|Gallbladder (MMHCC)|Anatomy|false|false||gallbladder
null|Gallbladder|Anatomy|false|false||gallbladder
null|Abdomen>Gallbladder|Anatomy|false|false||gallbladdernull|Walls of a building|Device|false|false||wallnull|Thickened|Finding|false|false||thickeningnull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Legal patent|Finding|false|false||Patentnull|Open|Modifier|false|false||Patentnull|Portal Venous System|Anatomy|false|false||portal venous systemnull|Hepatic|Anatomy|false|false||portalnull|Venous system|Anatomy|false|false||venous systemnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|System (basic dose form)|Drug|false|false||systemnull|System, LOINC Axis 4|Finding|false|false||system
null|System|Finding|false|false||systemnull|Device system|Device|false|false||system
null|System - kit|Device|false|false||systemnull|System (unit of presentation)|LabModifier|false|false||systemnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Encounter Special Courtesy - staff|Finding|false|false||staffnull|Staff|Subject|false|false||staffnull|On Staff|Modifier|false|false||staffnull|Procedure Practitioner Identifier Code Type - Radiologist|Finding|false|false||radiologistnull|radiologist|Subject|false|false||radiologistnull|null|Attribute|false|false||CT abdnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|LARGE1 wt Allele|Finding|false|false||Large
null|LARGE1 gene|Finding|false|false||Largenull|Large|LabModifier|false|false||Largenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Enlargement procedure|Procedure|false|false||enlargednull|Enlarged|Modifier|false|false||enlargednull|Edema|Finding|false|false||edematousnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Acute hepatitis|Disorder|false|false||acute hepatitisnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Small|LabModifier|false|false||Smallnull|Bilateral|Modifier|false|false||bilateralnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Left atrial structure|Anatomy|false|false||left atriumnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false||atriumnull|Right atrial structure|Anatomy|false|false||right atriumnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Heart Atrium|Anatomy|false|false||atriumnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|cardiac evaluation of ventricular wall thickness|Finding|false|false||ventricular wall thicknessnull|Wall of ventricle|Anatomy|false|false||ventricular wallnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Thick|Modifier|false|false||thicknessnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Tissue Specimen Code|Finding|false|false||tissuenull|Body tissue|Anatomy|false|false||tissuenull|Doppler studies|Procedure|false|false||Dopplernull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Diastole|Attribute|false|false||diastolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pulmonary Wedge Pressure|Attribute|false|false||PCWPnull|Ventricular Septal Defects|Disorder|false|false||ventricular septal defectnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Congenital septal defect of heart|Disorder|false|false||septal defect
null|Heart Septal Defects|Disorder|false|false||septal defectnull|Septal|Modifier|false|false||septalnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Diameter (qualifier value)|LabModifier|false|false||diametersnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Sequencing - Ascending|Finding|false|false||ascending
null|Ascend (action)|Finding|false|false||ascendingnull|Ascending|Modifier|false|false||ascendingnull|Age-Related Clonal Hematopoiesis|Finding|false|false||arch
null|ZBTB8OS gene|Finding|false|false||archnull|Arch of foot|Anatomy|false|false||arch
null|Structure of nucleus infundibularis hypothalami|Anatomy|false|false||arch
null|ARCH|Anatomy|false|false||archnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Leaflet|Finding|false|false||leafletnull|Leaflet Device|Device|false|false||leafletnull|Aortic Valve Insufficiency|Disorder|true|false||aortic regurgitationnull|Aorta|Anatomy|false|false||aorticnull|Regurgitation|Finding|true|false||regurgitation
null|Regurgitates after swallowing|Finding|true|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|true|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mitral Valve Prolapse Syndrome|Disorder|true|false||mitral valve prolapsenull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Ptosis|Disorder|true|false||prolapsenull|Pericardial effusion|Disorder|true|false||pericardial effusionnull|Pericardial effusion body substance|Finding|true|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|true|false||effusion
null|null|Finding|true|false||effusion
null|effusion|Finding|true|false||effusionnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|biventricular|Modifier|false|false||biventricularnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Diastolic dysfunction|Finding|true|false||diastolic dysfunctionnull|Diastole|Attribute|false|false||diastolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|true|false||dysfunctionnull|Dysfunction|Finding|true|false||dysfunction
null|physiopathological|Finding|true|false||dysfunction
null|Functional disorder|Finding|true|false||dysfunctionnull|Pulmonary Hypertension|Finding|true|false||pulmonary hypertensionnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Hypertensive disease|Disorder|true|false||hypertensionnull|Pathologic|Finding|false|false||pathologicnull|Valvular disease|Disorder|false|false||valvular diseasenull|Disease|Disorder|false|false||diseasenull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|ethanol|Drug|false|false||EtOH
null|ethanol|Drug|false|false||EtOHnull|year|Time|false|false||yearsnull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|new onset|Finding|false|false||new onsetnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Liver Failure|Disorder|false|false||liver failurenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Ascites|Disorder|false|false||ASCITESnull|Peritoneal Effusion|Finding|false|false||ASCITESnull|new onset|Finding|false|false||New onsetnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Serum-Ascites Albumin Gradient|Lab|false|false||SAAGnull|Supportive assistance|Finding|false|false||supportivenull|Portal Hypertension|Disorder|false|false||portal hypertensionnull|Hepatic|Anatomy|false|false||portalnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|alcoholic hepatitis with ascites|Disorder|false|false||alcoholic hepatitis with ascitesnull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Steroids|Drug|false|false||Steroids
null|Steroids|Drug|false|false||Steroidsnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Discriminate|Modifier|false|false||discriminatenull|Mathematical Factor|Finding|false|false||factor
null|Factor|Finding|false|false||factor
null|Feelings about Genomic Testing Results|Finding|false|false||factornull|Etiology aspects|Finding|false|false||etiologiesnull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Iron panel|Procedure|false|false||iron panelnull|null|Attribute|false|false||iron panelnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Groups|Finding|false|false||panelnull|Panel Device|Device|false|false||panelnull|Consistent with|Finding|true|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|true|false||consistentnull|HEMOCHROMATOSIS, TYPE 1|Disorder|false|false||hemochromatosis
null|Hemochromatosis|Disorder|false|false||hemochromatosisnull|HFE gene|Finding|false|false||hemochromatosisnull|Against Medical Advice|Finding|false|false||AMAnull|cytarabine/melphalan|Procedure|false|false||AMAnull|American Medical Association|Entity|false|false||AMAnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Autoimmune reaction|Finding|false|false||autoimmune
null|Autoimmune|Finding|false|false||autoimmunenull|Etiology aspects|Finding|false|false||causes
null|Etiology|Finding|false|false||causesnull|alpha 1-antitrypsin|Drug|false|false||Alpha 1 antitrypsin
null|alpha 1-proteinase inhibitor, human|Drug|false|false||Alpha 1 antitrypsin
null|alpha 1-proteinase inhibitor, human|Drug|false|false||Alpha 1 antitrypsin
null|alpha 1-proteinase inhibitor, human|Drug|false|false||Alpha 1 antitrypsin
null|alpha 1-antitrypsin|Drug|false|false||Alpha 1 antitrypsin
null|alpha 1-antitrypsin|Drug|false|false||Alpha 1 antitrypsinnull|ALPHA (substance)|Drug|false|false||Alpha
null|ALPHA (substance)|Drug|false|false||Alphanull|Greek letter alpha (qualifier value)|Finding|false|false||Alphanull|Alpha Value|Modifier|false|false||Alphanull|SERPINA5 protein, human|Drug|false|false||antitrypsin
null|SERPINA5 protein, human|Drug|false|false||antitrypsinnull|SERPINA1 gene|Finding|false|false||antitrypsinnull|Ceruloplasmin|Drug|false|false||ceruloplasmin
null|Ceruloplasmin|Drug|false|false||ceruloplasmin
null|CP protein, human|Drug|false|false||ceruloplasmin
null|CP protein, human|Drug|false|false||ceruloplasminnull|ferroxidase activity|Finding|false|false||ceruloplasmin
null|CP gene|Finding|false|false||ceruloplasminnull|Ceruloplasmin measurement|Procedure|false|false||ceruloplasminnull|Viral studies (procedure)|Procedure|false|false||Viral studiesnull|null|Attribute|false|false||Viral studiesnull|Viral|Finding|false|false||Viralnull|Scientific Study|Procedure|false|false||studiesnull|Immune response|Finding|false|false||immunity
null|Immune status|Finding|false|false||immunitynull|EPHB6 protein, human|Drug|false|false||Hep
null|EPHB6 protein, human|Drug|false|false||Hepnull|Hepatoerythropoietic Porphyria|Disorder|false|false||Hepnull|EPHB6 wt Allele, Human|Finding|false|false||Hep
null|EPHB6 gene|Finding|false|false||Hep
null|EPHB6 protein, human|Finding|false|false||Hep
null|HPSE wt Allele|Finding|false|false||Hep
null|DNLZ gene|Finding|false|false||Hepnull|HEP (body structure)|Anatomy|false|false||Hepnull|Histamine Equivalent Prick Unit|LabModifier|false|false||Hepnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|null|Attribute|false|false||CT abdnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Obstructed|Finding|false|false||obstructivenull|Lesion|Finding|false|false||lesionsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Paracentesis|Procedure|false|false||paracentesisnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Low-Dose Treatment|Procedure|false|false||Low-dosenull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Alcoholic Intoxication, Chronic|Disorder|false|false||ALCOHOLISMnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Ethanol measurement|Procedure|false|false||alcohol levelnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|clinical institute withdrawal assessment (CIWA) for alcohol|Finding|false|false||CIWAnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|MVI Regimen|Procedure|false|false||MVInull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|folate|Drug|false|false||folate
null|folate|Drug|false|false||folate
null|folate|Drug|false|false||folatenull|Folic acid measurement|Procedure|false|false||folatenull|Social Work (discipline)|Subject|false|false||social worknull|Social|Finding|false|false||socialnull|Work|Event|false|false||worknull|Contact Information|Finding|false|false||contact informationnull|Contact - HL7 Attribution|Finding|false|false||contact
null|Contact with|Finding|false|false||contact
null|Communication Contact|Finding|false|false||contactnull|contact person|Subject|false|false||contactnull|Physical contact|Phenomenon|false|false||contactnull|Personal Contact|Event|false|false||contactnull|Acknowledgement Detail Type - Information|Finding|false|false||information
null|Error severity - Information|Finding|false|false||information
null|Information|Finding|false|false||information
null|control act - information|Finding|false|false||informationnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Health Services, Outpatient|Procedure|false|false||outpatient treatment
null|Ambulatory Care|Procedure|false|false||outpatient treatmentnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Addictive Behavior|Disorder|false|false||addictionnull|Numerous|LabModifier|false|false||multiplenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Back Pain|Finding|false|false||BACK PAINnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Lidocaine Patch|Drug|false|false||lidocaine patchnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Breakthrough Pain|Finding|false|false||breakthrough painnull|Breakthrough|Modifier|false|false||breakthroughnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Leukocytosis|Disorder|false|false||LEUKOCYTOSISnull|Blood leukocyte number above reference range|Finding|false|false||LEUKOCYTOSISnull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|ciprofloxacin|Drug|false|false||ciprofloxacin
null|ciprofloxacin|Drug|false|false||ciprofloxacinnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Patient Discharge|Procedure|false|false||discharge, patientnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Polyarteritis Nodosa|Disorder|false|false||pannull|ADA2 wt Allele|Finding|false|false||pannull|proteasome-activating nucleotidase complex|Anatomy|false|false||pannull|Pansexuality|Subject|false|false||pannull|Pan <Homininae>|Entity|false|false||pan
null|Public Affairs Network of Cancer Centers|Entity|false|false||pan
null|Punjabi language|Entity|false|false||pannull|Plain chest X-ray|Procedure|false|false||CXRnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Cipro|Drug|false|false||Cipro
null|Cipro|Drug|false|false||Cipronull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Anemia, Macrocytic|Disorder|false|false||MACROCYTIC ANEMIAnull|TCN2 gene|Finding|false|false||MACROCYTIC ANEMIAnull|Mean corpuscular volume above reference range|Finding|false|false||MACROCYTICnull|Anemia|Disorder|false|false||ANEMIAnull|Anemia <Anemiaceae>|Entity|false|false||ANEMIAnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|folate|Drug|false|false||folate
null|folate|Drug|false|false||folate
null|folate|Drug|false|false||folatenull|Folic acid measurement|Procedure|false|false||folatenull|null|Attribute|false|false||nutritionalnull|Nutritional|Modifier|false|false||nutritionalnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Alcoholic Intoxication, Chronic|Disorder|false|false||alcoholismnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|Folate supplementation|Procedure|false|false||folate supplementationnull|folate|Drug|false|false||folate
null|folate|Drug|false|false||folate
null|folate|Drug|false|false||folatenull|Folic acid measurement|Procedure|false|false||folatenull|Dietary Supplementation|Procedure|false|false||supplementationnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Anxiety Disorders|Disorder|false|false||ANXIETY
null|Anxiety|Disorder|false|false||ANXIETYnull|Anxiety symptoms|Finding|false|false||ANXIETYnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Marked|Modifier|false|false||marked
null|Massive|Modifier|false|false||markednull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Benefit|LabModifier|false|false||benefitnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Selective Serotonin Reuptake Inhibitors|Drug|false|false||SSRI
null|Serotonin Reuptake Inhibitor [EPC]|Drug|false|false||SSRInull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Sinus Tachycardia|Disorder|false|false||SINUS TACHYCARDIAnull|continuous electrocardiogram sinus tachycardia|Finding|false|false||SINUS TACHYCARDIA
null|Sinus Tachycardia by ECG Finding|Finding|false|false||SINUS TACHYCARDIAnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||SINUS
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||SINUSnull|pathologic fistula|Disorder|false|false||SINUSnull|Sinus - general anatomical term|Anatomy|false|false||SINUS
null|Nasal sinus|Anatomy|false|false||SINUSnull|Tachycardia by ECG Finding|Finding|false|false||TACHYCARDIA
null|Tachycardia|Finding|false|false||TACHYCARDIAnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Application Context|Finding|false|false||context
null|Context|Finding|false|false||context
null|contextual factors|Finding|false|false||contextnull|Decompensated|Modifier|false|false||decompensatednull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Telemetry|Procedure|false|false||telemetrynull|Hospitalization|Procedure|false|false||hospitalizationnull|Constipation|Finding|false|false||CONSTIPATIONnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|sennosides, USP|Drug|false|false||senna
null|sennosides, USP|Drug|false|false||sennanull|Senna alexandrina|Entity|false|false||senna
null|Senna Plant|Entity|false|false||sennanull|Colace|Drug|false|false||colace
null|Colace|Drug|false|false||colacenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Multivitamin tablet|Drug|false|false||Multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acidnull|Folic acid measurement|Procedure|false|false||Folic Acidnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HClnull|Thiamine Drug Class|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|Thiamine Drug Class|Drug|false|false||Thiaminenull|Thiamine measurement|Procedure|false|false||Thiaminenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|ADHESIVE PATCH, MEDICATED|Device|false|false||Adhesive Patch, Medicatednull|Adhesives|Device|false|false||Adhesivenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Medicated|Drug|false|false||Medicatednull|Medicated (finding)|Finding|false|false||Medicatednull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|ADHESIVE PATCH, MEDICATED|Device|false|false||Adhesive Patch, Medicatednull|Adhesives|Device|false|false||Adhesivenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Medicated|Drug|false|false||Medicatednull|Medicated (finding)|Finding|false|false||Medicatednull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Apply (administration method)|Finding|false|false||Apply
null|Apply (instruction)|Finding|false|false||Apply
null|null|Finding|false|false||Apply
null|Apply|Finding|false|false||Applynull|Affected Area|Finding|false|false||affected areanull|Affected area of body|Anatomy|false|false||affected areanull|Involvement with|Finding|false|false||affected
null|Affecting|Finding|false|false||affectednull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|ADHESIVE PATCH, MEDICATED|Device|false|false||Adhesive Patch, Medicatednull|Adhesives|Device|false|false||Adhesivenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Medicated|Drug|false|false||Medicatednull|Medicated (finding)|Finding|false|false||Medicatednull|refill|Finding|false|false||Refillsnull|nicotine|Drug|true|false||Nicotine
null|nicotine|Drug|true|false||Nicotinenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Transdermal Route of Administration|Finding|false|false||Transdermal
null|transdermal|Finding|false|false||Transdermal
null|Transdermal (intended site)|Finding|false|false||Transdermalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|refill|Finding|false|false||Refillsnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|levofloxacin|Drug|false|false||Levofloxacin
null|levofloxacin|Drug|false|false||Levofloxacinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|Blood specimen|Finding|false|false||blood samplesnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|complete blood count with differential|Procedure|false|false||CBC with differentialnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Amount type - Differential|Finding|false|false||differentialnull|Differential (qualifier value)|Modifier|false|false||differential
null|Different|Modifier|false|false||differential
null|Differential - view|Modifier|false|false||differentialnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|Bilirubin|Drug|false|false||total bilirubin
null|Bilirubin|Drug|false|false||total bilirubinnull|Total bilirubin metabolic function|Finding|false|false||total bilirubinnull|Bilirubin, total measurement|Procedure|false|false||total bilirubinnull|Total bilirubin level|Lab|false|false||total bilirubinnull|Total|Modifier|false|false||totalnull|bilirubin preparation|Drug|false|false||bilirubin
null|bilirubin preparation|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubinnull|Bilirubin, total measurement|Procedure|false|false||bilirubin
null|blood bilirubin level test|Procedure|false|false||bilirubinnull|Alkaline Phosphatase|Drug|false|false||alkaline phosphatase
null|Alkaline Phosphatase|Drug|false|false||alkaline phosphatasenull|Alkaline phosphatase metabolic function|Finding|false|false||alkaline phosphatasenull|Alkaline phosphatase measurement|Procedure|false|false||alkaline phosphatasenull|Phosphoric Monoester Hydrolases|Drug|false|false||phosphatase
null|Phosphoric Monoester Hydrolases|Drug|false|false||phosphatasenull|phosphoric monoester hydrolase activity|Finding|false|false||phosphatasenull|Phosphatase (disposition)|Modifier|false|false||phosphatasenull|Albumin|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumin|Drug|false|false||albuminnull|Albumin metabolic function|Finding|false|false||albumin
null|ALB gene|Finding|false|false||albuminnull|Albumin measurement|Procedure|false|false||albuminnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|MT-CO3 gene|Finding|false|false||CO3null|Renal function|Finding|false|false||renal functionnull|Kidney Function Tests|Procedure|false|false||renal functionnull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucosenull|Glucose measurement|Procedure|false|false||glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||glucosenull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis|Procedure|false|false||Diagnosesnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Inflammation|Finding|false|false||inflammationnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|alcohol consumption (history)|Finding|false|false||alcohol consumption
null|Alcohol consumption|Finding|false|false||alcohol consumptionnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Consumption-archaic term for TB|Disorder|false|false||consumptionnull|biologic consumption|Finding|false|false||consumptionnull|Consumption of goods|Event|false|false||consumptionnull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Alcohol withdrawal syndrome|Disorder|false|false||alcohol withdrawalnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Withdrawal (dysfunction)|Disorder|false|false||withdrawalnull|Withdrawal - birth control|Procedure|false|false||withdrawalnull|Withdraw (activity)|Event|false|false||withdrawalnull|Liver function|Finding|false|false||liver functionnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Daily|Time|false|false||dailynull|Hematologic Tests|Procedure|false|false||blood testsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Tests (qualifier value)|Finding|false|false||testsnull|Laboratory Procedures|Procedure|false|false||testsnull|Liver function|Finding|false|false||liver functionnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Urinary tract infection|Disorder|false|false||urinary tract infectionnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Pneumonia|Disorder|false|false||pneumonianull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|More|LabModifier|false|false||morenull|day|Time|false|false||daysnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Infection of musculoskeletal system|Disorder|false|false||infectionsnull|Infection|Finding|false|false||infectionsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Abdomen|Anatomy|false|false||abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Leg|Anatomy|false|false||legsnull|null|Attribute|false|false||legsnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Work|Event|false|false||worknull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Heart Atrium|Anatomy|false|false||Atriumnull|Suite|Device|false|false||Suitenull|First floor|Modifier|false|false||first floornull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Sixth floor|Modifier|false|false||sixth floornull|Sixth|LabModifier|false|false||sixthnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Maxillary right canine mesial prosthesis|Device|false|false||6pmnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|folate|Drug|false|false||folate
null|folate|Drug|false|false||folate
null|folate|Drug|false|false||folatenull|Folic acid measurement|Procedure|false|false||folatenull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||generalnull|General medical service|Procedure|false|false||generalnull|Generalized|Modifier|false|false||generalnull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Lidocaine Patch|Drug|false|false||lidocaine patchnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Nicotine Transdermal Patch|Drug|false|false||nicotine patchnull|nicotine|Drug|false|false||nicotine
null|nicotine|Drug|false|false||nicotinenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Antibiotics|Drug|false|false||antibioticnull|Pneumonia|Disorder|false|false||pneumonianull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Accumulation|Finding|false|false||accumulationnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Appointments|Event|false|false||appointmentsnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions