 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Event|Event|Allergies|189,198|false|false|false|||Attending
Finding|Functional Concept|Allergies|189,198|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|224,229|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Chief Complaint|224,229|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Chief Complaint|224,238|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|Chief Complaint|230,238|false|false|false|||pressure
Finding|Finding|Chief Complaint|230,238|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Chief Complaint|230,238|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Chief Complaint|230,238|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Chief Complaint|230,238|false|false|false|C0033095||pressure
Finding|Classification|Chief Complaint|241,246|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|247,255|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|247,255|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|259,277|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|268,277|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|268,277|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|268,277|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|268,277|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|268,277|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|279,286|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Chief Complaint|279,286|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|History of Present Illness|365,385|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|past medical history
Finding|Functional Concept|History of Present Illness|370,377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|370,377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|370,377|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|370,377|false|false|false|C0199168|Medical service|medical
Finding|Finding|History of Present Illness|370,385|false|false|false|C0262926|Medical History|medical history
Finding|Finding|History of Present Illness|370,388|false|false|false|C0262926|Medical History|medical history of
Event|Event|History of Present Illness|378,385|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|378,385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|378,385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|378,385|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|378,388|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|390,393|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|390,393|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|390,393|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|390,393|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|390,393|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|390,393|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|390,393|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|390,393|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Location or Region|History of Present Illness|403,409|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|403,409|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|History of Present Illness|410,414|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|410,414|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|423,426|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|423,426|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|History of Present Illness|423,426|false|false|false|||LAD
Finding|Gene or Genome|History of Present Illness|423,426|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|History of Present Illness|439,447|false|false|false|||presents
Anatomy|Body Location or Region|History of Present Illness|454,459|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|454,459|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|454,468|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|History of Present Illness|460,468|false|false|false|||pressure
Finding|Finding|History of Present Illness|460,468|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|460,468|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|460,468|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|460,468|false|false|false|C0033095||pressure
Event|Event|History of Present Illness|475,479|false|false|false|||woke
Anatomy|Body Location or Region|History of Present Illness|507,512|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|507,512|false|false|false|C0741025|Chest problem|chest
Event|Event|History of Present Illness|514,522|false|false|false|||pressure
Finding|Finding|History of Present Illness|514,522|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|514,522|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|514,522|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|514,522|false|false|false|C0033095||pressure
Event|Event|History of Present Illness|532,538|false|false|false|||severe
Finding|Finding|History of Present Illness|532,538|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|532,538|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|History of Present Illness|563,566|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|History of Present Illness|563,566|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Drug|Organic Chemical|History of Present Illness|576,582|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|576,582|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|History of Present Illness|576,582|false|false|false|||relief
Finding|Finding|History of Present Illness|576,582|false|false|false|C0564405|Feeling relief|relief
Finding|Finding|History of Present Illness|595,607|false|false|false|C0425946|Short menstrual periods|short period
Event|Event|History of Present Illness|601,607|false|false|false|||period
Finding|Organism Function|History of Present Illness|601,607|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|History of Present Illness|601,607|false|false|false|C2347804|Clinical Trial Period|period
Finding|Finding|History of Present Illness|611,615|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|611,615|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|611,615|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|625,633|false|false|false|||radiated
Finding|Functional Concept|History of Present Illness|625,633|false|false|false|C0332301|Radiating to|radiated
Finding|Functional Concept|History of Present Illness|642,647|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|673,682|false|false|false|C0230348|Both upper arms|both arms
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|678,682|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|History of Present Illness|678,682|false|false|false|C5782111||arms
Disorder|Neoplastic Process|History of Present Illness|678,682|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|History of Present Illness|678,682|false|false|false|||arms
Finding|Gene or Genome|History of Present Illness|678,682|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|History of Present Illness|678,682|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|History of Present Illness|689,696|false|false|false|||reports
Event|Event|History of Present Illness|698,709|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|698,709|false|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|History of Present Illness|715,721|false|false|false|||denied
Attribute|Clinical Attribute|History of Present Illness|733,739|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|733,739|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|733,739|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|741,749|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|741,749|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|752,767|true|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|752,767|true|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|771,780|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|771,780|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|787,794|false|false|false|||reports
Event|Event|History of Present Illness|808,812|false|false|false|||felt
Event|Event|History of Present Illness|821,824|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|821,824|false|false|false|C0013404|Dyspnea|SOB
Disorder|Disease or Syndrome|History of Present Illness|842,851|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|History of Present Illness|842,851|false|false|false|||pneumonia
Finding|Gene or Genome|History of Present Illness|886,889|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|897,903|false|false|false|||denied
Event|Event|History of Present Illness|904,913|true|false|false|||worsening
Event|Event|History of Present Illness|914,921|true|false|false|||dyspnea
Finding|Finding|History of Present Illness|914,921|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|914,921|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|History of Present Illness|928,933|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|928,933|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|928,933|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|928,933|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|939,947|false|false|false|||improved
Event|Event|History of Present Illness|974,981|false|false|false|||minimal
Finding|Finding|History of Present Illness|990,994|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|990,994|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|990,994|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1002,1006|false|false|false|||went
Disorder|Disease or Syndrome|History of Present Illness|1014,1017|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1014,1017|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1014,1017|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1014,1017|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1014,1017|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1014,1017|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1014,1017|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1014,1017|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1014,1017|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1014,1017|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1014,1017|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|1020,1026|false|false|false|||office
Finding|Idea or Concept|History of Present Illness|1020,1026|false|false|false|C1549636|Address type - Office|office
Event|Event|History of Present Illness|1035,1040|false|false|false|||found
Finding|Finding|History of Present Illness|1051,1054|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1051,1054|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|History of Present Illness|1051,1059|false|false|false|C3844356|New LBBB|new LBBB
Disorder|Disease or Syndrome|History of Present Illness|1055,1059|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|History of Present Illness|1055,1059|false|false|false|||LBBB
Lab|Laboratory or Test Result|History of Present Illness|1055,1059|false|false|false|C0344420||LBBB
Disorder|Disease or Syndrome|History of Present Illness|1065,1073|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|History of Present Illness|1065,1073|false|false|false|||anterior
Event|Event|History of Present Illness|1077,1087|false|false|false|||elevations
Event|Event|History of Present Illness|1098,1109|false|false|false|||transferred
Drug|Organic Chemical|History of Present Illness|1135,1141|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|History of Present Illness|1135,1141|false|false|false|C0633084|Plavix|Plavix
Drug|Organic Chemical|History of Present Illness|1149,1156|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|History of Present Illness|1149,1156|false|false|false|C0004057|aspirin|Aspirin
Event|Event|History of Present Illness|1158,1165|false|false|false|||boluses
Drug|Biologically Active Substance|History of Present Illness|1169,1176|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|History of Present Illness|1169,1176|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|History of Present Illness|1169,1176|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|History of Present Illness|1169,1176|false|false|false|||heparin
Event|Event|History of Present Illness|1182,1193|false|false|false|||integrillin
Disorder|Disease or Syndrome|History of Present Illness|1200,1205|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|History of Present Illness|1200,1205|false|false|false|||STEMI
Finding|Finding|History of Present Illness|1200,1205|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Event|Event|History of Present Illness|1210,1216|false|false|false|||called
Event|Event|History of Present Illness|1221,1225|false|false|false|||went
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1233,1237|false|false|false|C0007430|Catheterization|cath
Event|Event|History of Present Illness|1238,1241|false|false|false|||lab
Finding|Gene or Genome|History of Present Illness|1238,1241|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|History of Present Illness|1238,1241|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|History of Present Illness|1245,1249|false|false|false|||Cath
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1245,1249|false|false|false|C0007430|Catheterization|Cath
Event|Event|History of Present Illness|1250,1256|false|false|false|||showed
Finding|Finding|History of Present Illness|1257,1265|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|History of Present Illness|1257,1265|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Event|Event|History of Present Illness|1266,1269|false|false|false|||SVG
Finding|Functional Concept|History of Present Illness|1271,1277|false|false|false|C0302891|Native (qualifier value)|Native
Finding|Finding|History of Present Illness|1283,1291|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|History of Present Illness|1283,1291|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Attribute|Clinical Attribute|History of Present Illness|1292,1300|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1301,1304|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|1301,1304|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|History of Present Illness|1301,1304|false|false|false|||LAD
Finding|Gene or Genome|History of Present Illness|1301,1304|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1318,1321|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|1318,1321|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|History of Present Illness|1318,1321|false|false|false|||LAD
Finding|Gene or Genome|History of Present Illness|1318,1321|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|History of Present Illness|1326,1335|false|false|false|||difficult
Finding|Finding|History of Present Illness|1326,1335|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|History of Present Illness|1350,1357|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1350,1357|false|false|false|C2699424|Concern|concern
Finding|Finding|History of Present Illness|1367,1375|false|false|false|C0332149|Possible|possible
Event|Event|History of Present Illness|1376,1386|false|false|false|||dissection
Finding|Pathologic Function|History of Present Illness|1376,1386|false|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1376,1386|false|false|false|C0012737|Tissue Dissection|dissection
Disorder|Disease or Syndrome|History of Present Illness|1392,1395|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|History of Present Illness|1392,1395|false|false|false|||BMS
Event|Event|History of Present Illness|1400,1406|false|false|false|||placed
Attribute|Clinical Attribute|History of Present Illness|1414,1422|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1423,1426|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|1423,1426|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|History of Present Illness|1423,1426|false|false|false|||LAD
Finding|Gene or Genome|History of Present Illness|1423,1426|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|History of Present Illness|1429,1435|false|false|false|C4522154|Distal Resection Margin|Distal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1436,1439|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|1436,1439|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|History of Present Illness|1436,1439|false|false|false|||LAD
Finding|Gene or Genome|History of Present Illness|1436,1439|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|History of Present Illness|1443,1453|false|false|false|C3842384|Diminutive|diminutive
Finding|Functional Concept|History of Present Illness|1474,1478|false|false|false|C1704338|diagnosis aspects|diag
Procedure|Diagnostic Procedure|History of Present Illness|1474,1478|false|false|false|C0011900|Diagnosis|diag
Event|Event|History of Present Illness|1479,1487|false|false|false|||branches
Finding|Finding|History of Present Illness|1505,1527|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|History of Present Illness|1521,1527|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1521,1527|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|History of Present Illness|1547,1550|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1547,1550|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|1547,1550|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|History of Present Illness|1547,1550|false|false|false|||SBP
Finding|Gene or Genome|History of Present Illness|1547,1550|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|1547,1550|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Anatomy|Anatomical Structure|History of Present Illness|1570,1575|false|false|false|C3714591|Floor (anatomic)|floor
Anatomy|Body Location or Region|History of Present Illness|1594,1599|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1594,1599|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1594,1604|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1594,1604|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1600,1604|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1600,1604|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1600,1604|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1600,1604|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|1600,1609|false|false|false|C0908489|Pain-Free|pain free
Event|Event|History of Present Illness|1605,1609|false|false|false|||free
Finding|Functional Concept|History of Present Illness|1605,1609|false|false|false|C0332296|Free of (attribute)|free
Event|Event|History of Present Illness|1615,1620|false|false|false|||feels
Event|Event|History of Present Illness|1621,1625|false|false|false|||well
Finding|Finding|History of Present Illness|1621,1625|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|1639,1645|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|1639,1645|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|1639,1645|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|1639,1648|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|1639,1656|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|1639,1656|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|History of Present Illness|1649,1656|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|1649,1656|false|false|false|C0449913|System|systems
Event|Event|History of Present Illness|1662,1668|true|false|false|||denies
Event|Event|History of Present Illness|1679,1686|true|false|false|||history
Finding|Conceptual Entity|History of Present Illness|1679,1686|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|1679,1686|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|1679,1686|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|1679,1689|true|false|false|C0262926|Medical History|history of
Attribute|Clinical Attribute|History of Present Illness|1690,1694|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1696,1702|true|false|false|C0042449|Veins|venous
Finding|Finding|History of Present Illness|1696,1713|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|History of Present Illness|1696,1713|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|History of Present Illness|1703,1713|true|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|1703,1713|true|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1715,1724|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|1715,1724|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|1715,1724|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|1715,1733|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|History of Present Illness|1725,1733|false|false|false|||embolism
Finding|Finding|History of Present Illness|1725,1733|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|History of Present Illness|1725,1733|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|History of Present Illness|1735,1743|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|1735,1743|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|History of Present Illness|1751,1755|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1751,1755|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1751,1755|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1760,1767|false|false|false|||surgery
Finding|Finding|History of Present Illness|1760,1767|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|1760,1767|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|1760,1767|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1760,1767|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|1769,1777|false|false|false|||myalgias
Finding|Sign or Symptom|History of Present Illness|1769,1777|false|false|false|C0231528|Myalgia|myalgias
Anatomy|Body Space or Junction|History of Present Illness|1779,1784|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|History of Present Illness|1779,1784|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|History of Present Illness|1779,1784|false|false|false|C0575044|Joint problem|joint
Finding|Sign or Symptom|History of Present Illness|1779,1790|false|false|false|C0003862|Arthralgia|joint pains
Event|Event|History of Present Illness|1785,1790|false|false|false|||pains
Finding|Sign or Symptom|History of Present Illness|1785,1790|false|false|false|C0030193|Pain|pains
Drug|Organic Chemical|History of Present Illness|1792,1797|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1792,1797|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1792,1797|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1792,1797|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1799,1809|false|false|false|||hemoptysis
Finding|Sign or Symptom|History of Present Illness|1799,1809|false|false|false|C0019079|Hemoptysis|hemoptysis
Finding|Pathologic Function|History of Present Illness|1811,1823|false|false|false|C0025222;C0474585|Melena|black stools
Finding|Sign or Symptom|History of Present Illness|1811,1823|false|false|false|C0025222;C0474585|Melena|black stools
Attribute|Clinical Attribute|History of Present Illness|1817,1823|false|false|false|C0489144||stools
Event|Event|History of Present Illness|1817,1823|false|false|false|||stools
Finding|Body Substance|History of Present Illness|1817,1823|false|false|false|C0015733|Feces|stools
Finding|Finding|History of Present Illness|1828,1831|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|History of Present Illness|1828,1831|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Sign or Symptom|History of Present Illness|1828,1838|false|false|false|C0278012|Red stools|red stools
Attribute|Clinical Attribute|History of Present Illness|1832,1838|false|false|false|C0489144||stools
Event|Event|History of Present Illness|1832,1838|false|false|false|||stools
Finding|Body Substance|History of Present Illness|1832,1838|false|false|false|C0015733|Feces|stools
Event|Event|History of Present Illness|1844,1850|false|false|false|||denies
Event|Event|History of Present Illness|1858,1864|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1858,1864|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1866,1872|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1866,1872|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|1876,1882|true|false|false|||rigors
Finding|Sign or Symptom|History of Present Illness|1876,1882|true|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Event|Event|History of Present Illness|1902,1908|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|1902,1908|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|1902,1908|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|1902,1911|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|1902,1919|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|1902,1919|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|History of Present Illness|1912,1919|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|1912,1919|false|false|false|C0449913|System|systems
Event|Event|History of Present Illness|1925,1933|false|false|false|||negative
Finding|Classification|History of Present Illness|1925,1933|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1925,1933|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1925,1933|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1941,1948|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|History of Present Illness|1941,1948|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|History of Present Illness|1949,1955|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|1949,1955|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|1949,1955|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|1949,1958|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|1949,1966|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|1949,1966|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|History of Present Illness|1959,1966|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|1959,1966|false|false|false|C0449913|System|systems
Event|Event|History of Present Illness|1970,1977|false|false|false|||notable
Disorder|Anatomical Abnormality|History of Present Illness|1982,1989|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|History of Present Illness|1982,1989|false|false|false|||absence
Finding|Functional Concept|History of Present Illness|1982,1989|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|History of Present Illness|1982,1992|false|false|false|C0332197|Absent|absence of
Anatomy|Body Location or Region|History of Present Illness|1993,1998|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1993,1998|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1993,2003|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1993,2003|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1999,2003|false|true|false|C2598155||pain
Event|Event|History of Present Illness|1999,2003|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1999,2003|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1999,2003|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2006,2013|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|2006,2013|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|2006,2013|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|2006,2025|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|History of Present Illness|2017,2025|false|false|false|C0015264|Exertion|exertion
Disorder|Disease or Syndrome|History of Present Illness|2027,2055|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|paroxysmal nocturnal dyspnea
Event|Event|History of Present Illness|2048,2055|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|2048,2055|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|2048,2055|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|2057,2066|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|2057,2066|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|2057,2066|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Anatomy|Body Location or Region|History of Present Illness|2069,2074|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|History of Present Illness|2069,2074|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Finding|Pathologic Function|History of Present Illness|2069,2080|false|false|false|C0235439|Ankle edema (finding)|ankle edema
Attribute|Clinical Attribute|History of Present Illness|2075,2080|false|false|false|C1717255||edema
Event|Event|History of Present Illness|2075,2080|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2075,2080|false|false|false|C0013604|Edema|edema
Event|Event|History of Present Illness|2082,2094|false|false|false|||palpitations
Finding|Finding|History of Present Illness|2082,2094|false|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|2096,2103|false|false|false|||syncope
Finding|Sign or Symptom|History of Present Illness|2096,2103|false|false|false|C0039070|Syncope|syncope
Finding|Finding|History of Present Illness|2096,2117|false|false|false|C3807340|Presyncope or syncope|syncope or presyncope
Event|Event|History of Present Illness|2107,2117|false|false|false|||presyncope
Finding|Sign or Symptom|History of Present Illness|2107,2117|false|false|false|C0700200|Presyncope|presyncope
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2149,2156|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Past Medical History|2149,2156|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|Past Medical History|2149,2161|false|false|false|C3176821|CARD.RISK|CARDIAC RISK
Finding|Finding|Past Medical History|2149,2169|false|false|false|C2024776|cardiac risk factors|CARDIAC RISK FACTORS
Event|Event|Past Medical History|2157,2161|false|false|false|||RISK
Finding|Idea or Concept|Past Medical History|2157,2161|false|false|false|C0035647|Risk|RISK
Attribute|Clinical Attribute|Past Medical History|2157,2169|false|false|false|C1830376||RISK FACTORS
Finding|Finding|Past Medical History|2157,2169|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Finding|Intellectual Product|Past Medical History|2157,2169|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Event|Event|Past Medical History|2162,2169|false|false|false|||FACTORS
Disorder|Disease or Syndrome|Past Medical History|2173,2181|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Past Medical History|2173,2181|false|false|false|||Diabetes
Disorder|Disease or Syndrome|Past Medical History|2185,2197|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Past Medical History|2185,2197|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|2202,2214|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|2202,2214|false|false|false|||Hypertension
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2220,2227|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Past Medical History|2220,2227|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|Patient History|2240,2244|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Patient History|2240,2244|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Location or Region|Patient History|2281,2287|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Patient History|2281,2287|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|Patient History|2288,2292|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Patient History|2288,2292|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Patient History|2299,2302|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|2299,2302|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Patient History|2299,2302|false|false|false|||LAD
Finding|Gene or Genome|Patient History|2299,2302|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Functional Concept|Patient History|2304,2316|false|false|false|C1522243|Percutaneous Route of Drug Administration|PERCUTANEOUS
Procedure|Therapeutic or Preventive Procedure|Patient History|2304,2339|false|false|false|C1532338|Percutaneous Coronary Intervention|PERCUTANEOUS CORONARY INTERVENTIONS
Anatomy|Body Part, Organ, or Organ Component|Patient History|2317,2325|false|false|false|C0018787|Heart|CORONARY
Attribute|Clinical Attribute|Patient History|2326,2339|false|false|false|C2979881||INTERVENTIONS
Event|Event|Patient History|2326,2339|false|false|false|||INTERVENTIONS
Procedure|Health Care Activity|Patient History|2326,2339|false|false|false|C0886296;C1273869|Intervention regimes;Nursing interventions|INTERVENTIONS
Finding|Individual Behavior|Patient History|2348,2354|true|false|false|C0562458|Pacing up and down|PACING
Disorder|Disease or Syndrome|Patient History|2355,2358|true|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|Patient History|2355,2358|true|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Event|Event|Patient History|2355,2358|true|false|false|||ICD
Finding|Gene or Genome|Patient History|2355,2358|true|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|Patient History|2355,2358|true|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|Patient History|2355,2358|true|false|false|C5575277|Icd Regimen|ICD
Event|Event|Patient History|2380,2387|true|false|false|||MEDICAL
Finding|Functional Concept|Patient History|2380,2387|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Idea or Concept|Patient History|2380,2387|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Intellectual Product|Patient History|2380,2387|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Procedure|Health Care Activity|Patient History|2380,2387|true|false|false|C0199168|Medical service|MEDICAL
Disorder|Disease or Syndrome|Patient History|2401,2404|true|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Patient History|2401,2404|true|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Patient History|2401,2404|true|false|false|||CVA
Finding|Functional Concept|Patient History|2413,2417|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|Patient History|2418,2427|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|Patient History|2436,2443|false|false|false|||infarct
Finding|Pathologic Function|Patient History|2436,2443|false|false|false|C0021308|Infarction|infarct
Drug|Biomedical or Dental Material|Patient History|2476,2479|false|false|false|C0039225|Tablet Dosage Form|tab
Event|Event|Patient History|2476,2479|false|false|false|||tab
Drug|Organic Chemical|Patient History|2483,2489|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Patient History|2483,2489|false|false|false|C0633084|Plavix|plavix
Event|Event|Patient History|2483,2489|false|false|false|||plavix
Disorder|Disease or Syndrome|Patient History|2498,2518|false|false|false|C0020443|Hypercholesterolemia|hypercholesterolemia
Event|Event|Patient History|2498,2518|false|false|false|||hypercholesterolemia
Finding|Finding|Patient History|2498,2518|false|false|false|C1522133|Hypercholesterolemia result|hypercholesterolemia
Event|Event|Patient History|2530,2533|false|false|false|||PFO
Event|Event|Patient History|2545,2557|false|false|false|||Degereration
Finding|Conceptual Entity|Family Medical History|2600,2606|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|2600,2606|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|Family Medical History|2607,2611|false|false|false|||died
Disorder|Disease or Syndrome|Family Medical History|2619,2622|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2619,2622|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|2619,2622|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|2619,2622|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|2619,2622|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|2619,2622|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|2619,2622|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2619,2622|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|Family Medical History|2626,2629|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|2626,2629|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|2626,2629|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|2626,2629|false|false|false|||age
Finding|Idea or Concept|Family Medical History|2640,2646|false|false|false|C1546508|Relationship - Mother|mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2651,2658|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|2651,2658|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|2651,2658|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Family Medical History|2651,2658|false|false|false|||stomach
Finding|Finding|Family Medical History|2651,2658|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2651,2658|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|2651,2665|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|Family Medical History|2659,2665|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|2659,2665|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2670,2674|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|Family Medical History|2670,2674|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|Family Medical History|2670,2674|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Neoplastic Process|Family Medical History|2670,2681|false|false|false|C0279530;C0585442|Malignant Bone Neoplasm;Osteosarcoma of bone|bone cancer
Disorder|Neoplastic Process|Family Medical History|2675,2681|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|2675,2681|false|false|false|||cancer
Event|Event|General Exam|2700,2707|false|false|false|||GENERAL
Finding|Classification|General Exam|2700,2707|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2700,2707|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|2709,2713|false|false|false|||WDWN
Disorder|Disease or Syndrome|General Exam|2717,2720|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2717,2720|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2717,2720|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2717,2720|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2717,2720|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2717,2720|false|false|false|||NAD
Finding|Finding|General Exam|2717,2720|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|General Exam|2722,2730|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|General Exam|2735,2739|false|false|false|C2713234||Mood
Event|Event|General Exam|2735,2739|false|false|false|||Mood
Finding|Conceptual Entity|General Exam|2735,2739|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|2735,2739|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|2735,2739|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|General Exam|2741,2747|false|false|false|||affect
Event|Event|General Exam|2748,2759|false|false|false|||appropriate
Anatomy|Body Location or Region|General Exam|2763,2768|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|2770,2774|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|General Exam|2776,2782|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|2776,2782|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|2776,2782|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|2776,2782|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|2783,2792|false|false|false|||anicteric
Finding|Finding|General Exam|2783,2792|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|2794,2799|false|false|false|||PERRL
Finding|Finding|General Exam|2794,2799|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|2801,2805|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|2807,2818|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|2807,2818|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|2807,2818|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|General Exam|2807,2818|true|false|false|||Conjunctiva
Finding|Body Substance|General Exam|2807,2818|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|2807,2818|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|2807,2818|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|General Exam|2834,2840|true|false|false|||pallor
Finding|Finding|General Exam|2834,2840|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|General Exam|2844,2852|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|2844,2852|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|2860,2864|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|2860,2864|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|2860,2864|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|2860,2864|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|2860,2871|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|2865,2871|true|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|2865,2871|true|false|false|C1561514||mucosa
Event|Event|General Exam|2876,2887|true|false|false|||xanthalesma
Anatomy|Body Location or Region|General Exam|2892,2896|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2892,2896|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2892,2896|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|2898,2904|false|false|false|||Supple
Finding|Functional Concept|General Exam|2898,2904|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|2910,2913|false|false|false|||JVP
Finding|Finding|General Exam|2910,2913|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|2925,2932|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|2925,2932|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|2934,2937|false|false|false|||PMI
Finding|Finding|General Exam|2934,2937|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|General Exam|2934,2937|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|General Exam|2953,2970|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|General Exam|2965,2970|false|false|false|C0282173|Space (Astronomy)|space
Event|Event|General Exam|2972,2985|false|false|false|||midclavicular
Drug|Biologically Active Substance|General Exam|2987,2991|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2987,2991|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|General Exam|2987,2991|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|General Exam|2987,2991|false|false|false|||line
Finding|Intellectual Product|General Exam|2987,2991|false|false|false|C1546701|line source specimen code|line
Event|Event|General Exam|3019,3020|true|false|false|||g
Event|Event|General Exam|3025,3032|true|false|false|||thrills
Finding|Finding|General Exam|3025,3032|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|General Exam|3034,3039|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|General Exam|3057,3062|false|false|false|C0024109|Lung|LUNGS
Anatomy|Body Location or Region|General Exam|3067,3072|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|3067,3072|true|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|General Exam|3067,3077|true|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|3067,3077|true|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Disorder|Anatomical Abnormality|General Exam|3067,3089|true|false|false|C3164427|Deformity of chest wall|chest wall deformities
Disorder|Congenital Abnormality|General Exam|3078,3089|true|false|false|C0000768|Congenital Abnormality|deformities
Event|Event|General Exam|3078,3089|true|false|false|||deformities
Disorder|Acquired Abnormality|General Exam|3091,3100|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Congenital Abnormality|General Exam|3091,3100|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Disease or Syndrome|General Exam|3091,3100|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Event|Event|General Exam|3091,3100|true|false|false|||scoliosis
Disorder|Acquired Abnormality|General Exam|3104,3112|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Anatomical Abnormality|General Exam|3104,3112|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Congenital Abnormality|General Exam|3104,3112|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Event|Event|General Exam|3104,3112|true|false|false|||kyphosis
Finding|Finding|General Exam|3104,3112|true|false|false|C2115817|kyphosis|kyphosis
Attribute|Clinical Attribute|General Exam|3114,3118|true|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|3114,3118|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|General Exam|3114,3118|true|false|false|||Resp
Event|Event|General Exam|3125,3134|true|false|false|||unlabored
Finding|Functional Concept|General Exam|3125,3134|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|General Exam|3139,3155|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|3139,3159|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|3149,3155|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|3149,3155|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|3156,3159|true|false|false|||use
Finding|Functional Concept|General Exam|3156,3159|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|3156,3159|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Amino Acid, Peptide, or Protein|General Exam|3161,3164|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|3161,3164|true|false|false|||CTA
Finding|Gene or Genome|General Exam|3161,3164|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|3161,3164|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|General Exam|3181,3189|true|false|false|||crackles
Finding|Finding|General Exam|3181,3189|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|General Exam|3191,3198|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3191,3198|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3202,3209|true|false|false|||rhonchi
Finding|Finding|General Exam|3202,3209|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|3213,3220|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3213,3220|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3213,3220|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3213,3220|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3222,3226|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|3222,3226|false|false|false|||Soft
Event|Event|General Exam|3228,3232|false|false|false|||NTND
Event|Event|General Exam|3237,3240|true|false|false|||HSM
Finding|Gene or Genome|General Exam|3237,3240|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|General Exam|3244,3254|true|false|false|||tenderness
Finding|Mental Process|General Exam|3244,3254|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3244,3254|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|General Exam|3256,3259|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|3256,3259|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|General Exam|3260,3265|true|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|3260,3265|true|false|false|C0869784|Procedure on aorta|aorta
Event|Event|General Exam|3271,3279|true|false|false|||enlarged
Event|Event|General Exam|3283,3292|true|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|3283,3292|true|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|3308,3314|true|false|false|||bruits
Finding|Finding|General Exam|3308,3314|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|General Exam|3318,3329|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|General Exam|3341,3348|false|false|false|C0015811|Femur|Femoral
Anatomy|Body Part, Organ, or Organ Component|General Exam|3349,3355|false|false|false|C0227952|Foreskin of penis|sheath
Event|Activity|General Exam|3359,3364|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|3359,3364|false|false|false|||place
Finding|Functional Concept|General Exam|3359,3364|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3359,3364|false|false|false|C1533810||place
Finding|Functional Concept|General Exam|3368,3373|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|3374,3379|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|groin
Anatomy|Body System|General Exam|3383,3387|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3383,3387|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3383,3387|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|3383,3387|false|false|false|||SKIN
Finding|Body Substance|General Exam|3383,3387|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3383,3387|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|General Exam|3392,3398|true|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|3392,3409|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|3399,3409|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|General Exam|3399,3409|true|false|false|||dermatitis
Event|Event|General Exam|3411,3417|true|false|false|||ulcers
Finding|Pathologic Function|General Exam|3411,3417|true|false|false|C0041582|Ulcer|ulcers
Event|Event|General Exam|3419,3424|true|false|false|||scars
Finding|Finding|General Exam|3419,3424|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|General Exam|3419,3424|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|General Exam|3429,3438|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|General Exam|3429,3438|false|false|false|||xanthomas
Drug|Food|General Exam|3442,3448|false|false|false|C5890763||PULSES
Event|Event|General Exam|3442,3448|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|3442,3448|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3442,3448|false|false|false|C0034107|Pulse taking|PULSES
Finding|Functional Concept|General Exam|3452,3457|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|3459,3466|false|false|false|C0007272|Carotid Arteries|Carotid
Finding|Functional Concept|General Exam|3485,3489|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3491,3498|false|false|false|C0007272|Carotid Arteries|Carotid
Event|Event|General Exam|3538,3541|false|false|false|||EKG
Finding|Intellectual Product|General Exam|3538,3541|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|3538,3541|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|General Exam|3544,3547|false|false|false|||new
Finding|Finding|General Exam|3544,3547|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|3544,3547|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|General Exam|3544,3552|false|false|false|C3844356|New LBBB|new LBBB
Disorder|Disease or Syndrome|General Exam|3548,3552|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Event|Event|General Exam|3548,3552|false|false|false|||LBBB
Lab|Laboratory or Test Result|General Exam|3548,3552|false|false|false|C0344420||LBBB
Event|Event|General Exam|3558,3561|false|false|false|||STE
Finding|Gene or Genome|General Exam|3558,3561|false|false|false|C1420459;C3811127|SULT1E1 gene;SULT1E1 wt Allele|STE
Procedure|Diagnostic Procedure|General Exam|3608,3617|false|false|false|C0039451|Telemetry|TELEMETRY
Finding|Molecular Function|General Exam|3619,3622|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|General Exam|3619,3622|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Procedure|Diagnostic Procedure|General Exam|3644,3658|false|false|false|C0013516|Echocardiography|ECHOCARDIOGRAM
Event|Event|General Exam|3661,3668|false|false|false|||pending
Finding|Idea or Concept|General Exam|3661,3668|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Disorder|Neoplastic Process|General Exam|3669,3672|false|false|false|C1266159|Trophoblastic tumor, epithelioid|ETT
Event|Event|General Exam|3669,3672|false|false|false|||ETT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3683,3690|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3683,3690|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Diagnostic Procedure|General Exam|3683,3695|false|false|false|C0018795|Cardiac Catheterization Procedures|CARDIAC CATH
Event|Event|General Exam|3691,3695|false|false|false|||CATH
Procedure|Therapeutic or Preventive Procedure|General Exam|3691,3695|false|false|false|C0007430|Catheterization|CATH
Drug|Organic Chemical|General Exam|3699,3703|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Pharmacologic Substance|General Exam|3699,3703|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Vitamin|General Exam|3699,3703|false|false|false|C2828271|levomefolate calcium|LMCA
Event|Event|General Exam|3699,3703|false|false|false|||LMCA
Attribute|Clinical Attribute|General Exam|3709,3715|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3716,3719|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3716,3719|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3716,3719|false|false|false|||LAD
Finding|Gene or Genome|General Exam|3716,3719|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|General Exam|3721,3729|false|false|false|C0028778;C1947917|Obstruction;Occluded|Occluded
Finding|Functional Concept|General Exam|3721,3729|false|false|false|C0028778;C1947917|Obstruction;Occluded|Occluded
Event|Event|General Exam|3730,3739|false|false|false|||difficult
Finding|Finding|General Exam|3730,3739|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|General Exam|3754,3761|false|false|false|||crossed
Attribute|Clinical Attribute|General Exam|3778,3786|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3787,3790|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3787,3790|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3787,3790|false|false|false|||LAD
Finding|Gene or Genome|General Exam|3787,3790|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|General Exam|3793,3799|false|false|false|C4522154|Distal Resection Margin|Distal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3800,3803|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3800,3803|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3800,3803|false|false|false|||LAD
Finding|Gene or Genome|General Exam|3800,3803|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|3812,3820|false|false|false|||diseased
Drug|Amino Acid, Peptide, or Protein|General Exam|3824,3827|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Drug|Enzyme|General Exam|3824,3827|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Event|Event|General Exam|3824,3827|false|false|false|||LCX
Finding|Gene or Genome|General Exam|3824,3827|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCX
Finding|Finding|General Exam|3829,3837|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|General Exam|3829,3837|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Drug|Amino Acid, Peptide, or Protein|General Exam|3847,3850|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Drug|Enzyme|General Exam|3847,3850|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Event|Event|General Exam|3847,3850|false|false|false|||LCX
Finding|Gene or Genome|General Exam|3847,3850|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCX
Event|Event|General Exam|3851,3854|false|false|false|||RCA
Finding|Finding|General Exam|3856,3864|false|false|false|C0028778;C1947917|Obstruction;Occluded|Occluded
Finding|Functional Concept|General Exam|3856,3864|false|false|false|C0028778;C1947917|Obstruction;Occluded|Occluded
Event|Event|Hospital Course|3920,3927|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|3920,3927|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3920,3927|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|3920,3927|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3920,3930|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|3931,3934|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3931,3934|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3931,3934|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3931,3934|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3931,3934|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3931,3934|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3931,3934|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3931,3934|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|3940,3949|false|false|false|||presented
Disorder|Disease or Syndrome|Hospital Course|3958,3963|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|Hospital Course|3958,3963|false|false|false|||STEMI
Finding|Finding|Hospital Course|3958,3963|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Event|Event|Hospital Course|3968,3983|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3968,3983|false|false|false|C0007430|Catheterization|catheterization
Event|Event|Hospital Course|4006,4011|false|false|false|||found
Finding|Finding|Hospital Course|4020,4046|false|false|false|C0748164|Multiple Pulmonary Nodules|multiple pulmonary nodules
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4029,4038|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|4029,4038|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|4029,4038|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|Hospital Course|4029,4046|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|Hospital Course|4039,4046|false|false|false|||nodules
Event|Event|Hospital Course|4047,4057|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|4047,4057|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|4047,4062|false|false|false|C0332290|Consistent with|consistent with
Disorder|Neoplastic Process|Hospital Course|4064,4078|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|4064,4078|false|false|false|||adenocarcinoma
Disorder|Disease or Syndrome|Hospital Course|4086,4091|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|Hospital Course|4086,4091|false|false|false|||STEMI
Finding|Finding|Hospital Course|4086,4091|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Event|Event|Hospital Course|4096,4105|false|false|false|||presented
Disorder|Disease or Syndrome|Hospital Course|4114,4122|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Disorder|Disease or Syndrome|Hospital Course|4123,4128|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|Hospital Course|4123,4128|false|false|false|||STEMI
Finding|Finding|Hospital Course|4123,4128|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Event|Event|Hospital Course|4140,4144|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|4140,4144|false|false|false|C0035647|Risk|risk
Event|Event|Hospital Course|4146,4151|false|false|false|||score
Finding|Finding|Hospital Course|4146,4151|false|false|false|C0449820|Score|score
Event|Event|Hospital Course|4158,4168|false|false|false|||indicating
Event|Event|Hospital Course|4175,4179|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|4175,4179|false|false|false|C0035647|Risk|risk
Event|Event|Hospital Course|4194,4203|false|false|false|||mortality
Event|Event|Hospital Course|4205,4208|false|false|false|||new
Finding|Finding|Hospital Course|4205,4208|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|4205,4208|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Hospital Course|4213,4222|false|false|false|||recurrent
Finding|Finding|Hospital Course|4230,4236|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|4230,4236|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Hospital Course|4247,4255|false|false|false|||ischemia
Finding|Pathologic Function|Hospital Course|4247,4255|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4247,4255|false|false|false|C4321499|Ischemia Procedure|ischemia
Event|Event|Hospital Course|4266,4272|false|false|false|||urgent
Finding|Intellectual Product|Hospital Course|4266,4272|false|false|false|C1546403;C1546845;C1547230;C1561556|Admission Type - Urgent;Certification patient type - Urgent;Triage Code - Urgent;Visit Priority Code - Urgent|urgent
Event|Event|Hospital Course|4274,4291|false|false|false|||revascularization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4274,4291|false|false|false|C0581603||revascularization
Event|Event|Hospital Course|4298,4301|false|false|false|||SVG
Event|Event|Hospital Course|4302,4307|false|false|false|||found
Finding|Intellectual Product|Hospital Course|4314,4324|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|Hospital Course|4325,4333|false|false|false|||occluded
Finding|Finding|Hospital Course|4325,4333|false|true|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|Hospital Course|4325,4333|false|true|false|C0028778;C1947917|Obstruction;Occluded|occluded
Disorder|Disease or Syndrome|Hospital Course|4341,4344|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Hospital Course|4341,4344|false|false|false|||BMS
Event|Event|Hospital Course|4349,4355|false|false|false|||placed
Attribute|Clinical Attribute|Hospital Course|4363,4371|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4372,4375|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|4372,4375|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Hospital Course|4372,4375|false|false|false|||LAD
Finding|Gene or Genome|Hospital Course|4372,4375|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|Hospital Course|4389,4395|false|false|false|||timing
Finding|Intellectual Product|Hospital Course|4389,4395|false|false|false|C1704250|Timing, LOINC Axis 3|timing
Event|Event|Hospital Course|4408,4417|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|4408,4417|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4408,4417|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Gene or Genome|Hospital Course|4433,4436|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|4445,4452|false|false|false|||thought
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4462,4465|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|4462,4465|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|4462,4465|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|Hospital Course|4471,4478|false|false|false|||managed
Finding|Idea or Concept|Hospital Course|4482,4486|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|Hospital Course|4482,4486|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Event|Event|Hospital Course|4487,4500|false|false|false|||revascularize
Event|Event|Hospital Course|4519,4527|false|false|false|||supplied
Event|Event|Hospital Course|4536,4539|false|false|false|||RCA
Event|Event|Hospital Course|4550,4557|false|false|false|||started
Event|Event|Hospital Course|4561,4568|false|false|false|||routine
Finding|Idea or Concept|Hospital Course|4561,4568|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|Hospital Course|4561,4568|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|Hospital Course|4561,4568|false|false|false|C1979801|Routine coag|routine
Anatomy|Body Space or Junction|Hospital Course|4569,4572|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|Hospital Course|4569,4572|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4569,4572|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|Hospital Course|4569,4572|false|false|false|C4042561|ACSS2 protein, human|ACS
Finding|Gene or Genome|Hospital Course|4569,4572|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|Hospital Course|4569,4572|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|Hospital Course|4569,4572|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Attribute|Clinical Attribute|Hospital Course|4573,4584|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4573,4584|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|4573,4584|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|4573,4584|false|false|false|C4284232|Medications|medications
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4586,4598|false|false|false|C0253563|eptifibatide|eptifibatide
Drug|Pharmacologic Substance|Hospital Course|4586,4598|false|false|false|C0253563|eptifibatide|eptifibatide
Event|Event|Hospital Course|4586,4598|false|false|false|||eptifibatide
Disorder|Disease or Syndrome|Hospital Course|4607,4610|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4607,4610|false|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|Hospital Course|4607,4610|false|false|false|C1568891|HGS protein, human|hrs
Event|Event|Hospital Course|4607,4610|false|false|false|||hrs
Finding|Gene or Genome|Hospital Course|4607,4610|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Drug|Organic Chemical|Hospital Course|4612,4618|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|4612,4618|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|4612,4618|false|false|false|||plavix
Drug|Organic Chemical|Hospital Course|4626,4633|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|4626,4633|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|4634,4639|false|false|false|||325mg
Drug|Organic Chemical|Hospital Course|4641,4651|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|4641,4651|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|4641,4651|false|false|false|||metoprolol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4653,4662|false|false|false|C0006938|captopril|captopril
Drug|Pharmacologic Substance|Hospital Course|4653,4662|false|false|false|C0006938|captopril|captopril
Event|Event|Hospital Course|4653,4662|false|false|false|||captopril
Drug|Organic Chemical|Hospital Course|4669,4681|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|4669,4681|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|4669,4681|false|false|false|||atorvastatin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4684,4691|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|4684,4691|false|false|false|C1314974|Cardiac attachment|Cardiac
Attribute|Clinical Attribute|Hospital Course|4684,4699|false|false|false|C2926589||Cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4684,4699|false|false|false|C0443763|Cardiac enzymes|Cardiac enzymes
Drug|Enzyme|Hospital Course|4684,4699|false|false|false|C0443763|Cardiac enzymes|Cardiac enzymes
Procedure|Laboratory Procedure|Hospital Course|4684,4699|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|Cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4692,4699|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|Hospital Course|4692,4699|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|Hospital Course|4692,4699|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Event|Event|Hospital Course|4692,4699|false|false|false|||enzymes
Finding|Functional Concept|Hospital Course|4692,4699|false|false|false|C0014445|enzymology|enzymes
Event|Event|Hospital Course|4700,4707|false|false|false|||trended
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4745,4749|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CKMB
Drug|Enzyme|Hospital Course|4745,4749|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CKMB
Event|Event|Hospital Course|4745,4749|false|false|false|||CKMB
Event|Event|Hospital Course|4778,4785|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|4778,4785|false|false|false|C2699424|Concern|concern
Finding|Intellectual Product|Hospital Course|4791,4796|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|4791,4810|false|false|false|C0264714|Acute heart failure|acute heart failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4797,4802|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|4797,4802|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|4797,4802|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Hospital Course|4797,4810|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Hospital Course|4803,4810|false|false|false|||failure
Finding|Functional Concept|Hospital Course|4803,4810|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|4803,4810|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|4803,4810|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Functional Concept|Hospital Course|4816,4824|false|false|false|C0475224|Ischemic|ischemic
Drug|Biologically Active Substance|Hospital Course|4832,4838|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|4832,4838|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|4832,4838|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4832,4838|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|4839,4850|false|false|false|||requirement
Finding|Functional Concept|Hospital Course|4839,4850|false|false|false|C1514873|Requirement|requirement
Event|Event|Hospital Course|4871,4876|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4892,4895|true|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|Hospital Course|4892,4895|true|false|false|C5703311|Radiolucent Lines|RLL
Disorder|Disease or Syndrome|Hospital Course|4896,4905|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|4896,4905|true|false|false|||pneumonia
Finding|Idea or Concept|Hospital Course|4914,4925|true|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4926,4935|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|4926,4935|true|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|4926,4935|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|4926,4941|true|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|4936,4941|true|false|false|C1717255||edema
Event|Event|Hospital Course|4936,4941|true|false|false|||edema
Finding|Pathologic Function|Hospital Course|4936,4941|true|false|false|C0013604|Edema|edema
Event|Event|Hospital Course|4943,4946|true|false|false|||see
Event|Event|Hospital Course|4956,4960|false|false|false|||ECHO
Procedure|Health Care Activity|Hospital Course|4956,4960|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4956,4960|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|Hospital Course|4961,4967|false|false|false|||showed
Event|Event|Hospital Course|4968,4976|false|false|false|||moderate
Finding|Finding|Hospital Course|4968,4976|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|4968,4976|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|Hospital Course|4981,4987|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|4981,4987|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|Hospital Course|4997,5001|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|Hospital Course|4997,5034|false|false|false|C1277187|Left ventricular systolic dysfunction|left ventricular systolic dysfunction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5002,5013|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|Hospital Course|5014,5022|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|Hospital Course|5014,5034|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|Hospital Course|5023,5034|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|5023,5034|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|5023,5034|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|5023,5034|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|5023,5034|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Disorder|Disease or Syndrome|Hospital Course|5041,5049|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Hospital Course|5041,5049|false|false|false|||anterior
Event|Event|Hospital Course|5067,5075|false|false|false|||akinesis
Event|Event|Hospital Course|5080,5088|false|false|false|||inferior
Finding|Social Behavior|Hospital Course|5080,5088|false|false|false|C0678975|inferiority|inferior
Event|Event|Hospital Course|5104,5115|false|false|false|||hypokinesis
Finding|Finding|Hospital Course|5104,5115|false|false|false|C0086439|Hypokinesia|hypokinesis
Finding|Body Substance|Hospital Course|5129,5136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5129,5136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5129,5136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5142,5149|false|false|false|||started
Drug|Organic Chemical|Hospital Course|5153,5161|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|5153,5161|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Hospital Course|5153,5161|false|false|false|||coumadin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5167,5178|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|Hospital Course|5167,5187|false|false|false|C0876993|Cardiac ventricular thrombosis|ventricular thrombus
Event|Event|Hospital Course|5179,5187|false|false|false|||thrombus
Finding|Pathologic Function|Hospital Course|5179,5187|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|Hospital Course|5188,5199|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5188,5199|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|5228,5240|false|false|false|||discontinued
Event|Event|Hospital Course|5244,5248|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|5244,5248|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|Hospital Course|5244,5251|false|false|false|C0035647|Risk|risk of
Finding|Finding|Hospital Course|5244,5260|false|false|false|C3251812|Bleeding risk|risk of bleeding
Event|Event|Hospital Course|5252,5260|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|5252,5260|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|5272,5279|false|false|false|||benefit
Finding|Finding|Hospital Course|5285,5292|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|Hospital Course|5285,5292|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Event|Event|Hospital Course|5300,5315|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|5300,5315|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Body Substance|Hospital Course|5317,5324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5317,5324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5317,5324|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5329,5338|false|false|false|||maintaing
Event|Event|Hospital Course|5340,5351|false|false|false|||saturations
Phenomenon|Natural Phenomenon or Process|Hospital Course|5340,5351|false|false|false|C0522534|Saturated|saturations
Finding|Finding|Hospital Course|5355,5358|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|5355,5358|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Biomedical or Dental Material|Hospital Course|5374,5382|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|5374,5382|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|5374,5382|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|5395,5398|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|5395,5398|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|5400,5406|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5407,5410|false|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|Hospital Course|5407,5410|false|false|false|C5703311|Radiolucent Lines|RLL
Disorder|Disease or Syndrome|Hospital Course|5411,5420|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|5411,5420|false|false|false|||pneumonia
Event|Event|Hospital Course|5426,5433|false|false|false|||patient
Finding|Body Substance|Hospital Course|5426,5433|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5426,5433|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5426,5433|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5451,5458|false|false|false|||started
Drug|Antibiotic|Hospital Course|5463,5474|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|5463,5474|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|5463,5474|false|false|false|||ceftriaxone
Drug|Antibiotic|Hospital Course|5476,5488|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|5476,5488|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|5476,5488|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|5476,5488|false|false|false|||azithromycin
Drug|Organic Chemical|Hospital Course|5490,5503|false|false|false|C0025872|metronidazole|metronidazole
Drug|Pharmacologic Substance|Hospital Course|5490,5503|false|false|false|C0025872|metronidazole|metronidazole
Event|Event|Hospital Course|5490,5503|false|false|false|||metronidazole
Finding|Body Substance|Hospital Course|5513,5520|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5513,5520|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5513,5520|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5526,5533|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5526,5533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5526,5533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5526,5533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5544,5547|false|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|Hospital Course|5544,5547|false|false|false|C5703311|Radiolucent Lines|RLL
Disorder|Disease or Syndrome|Hospital Course|5548,5557|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|5548,5557|false|false|false|||pneumonia
Procedure|Diagnostic Procedure|Hospital Course|5561,5568|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|5564,5568|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|5564,5568|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|5589,5595|false|false|false|||showed
Finding|Finding|Hospital Course|5596,5602|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|5596,5602|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|Hospital Course|5603,5608|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5603,5619|false|false|false|C1261075|Structure of right lower lobe of lung|right lower lobe
Anatomy|Body Location or Region|Hospital Course|5609,5614|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|5609,5614|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5609,5619|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5615,5619|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|5615,5619|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|Hospital Course|5620,5633|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Hospital Course|5620,5633|false|false|false|||consolidation
Finding|Finding|Hospital Course|5649,5652|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|5649,5652|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|Hospital Course|5662,5666|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5662,5666|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|5662,5666|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|5662,5666|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Hospital Course|5662,5674|false|false|false|C0034079||lung nodules
Event|Event|Hospital Course|5667,5674|false|false|false|||nodules
Finding|Body Substance|Hospital Course|5681,5687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|5681,5687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Finding|Hospital Course|5681,5696|false|false|false|C0551076|Sputum cytology (finding)|sputum cytology
Procedure|Laboratory Procedure|Hospital Course|5681,5696|false|false|false|C1521752|Sputum Cytology Screening|sputum cytology
Lab|Laboratory or Test Result|Hospital Course|5681,5705|false|false|false|C0580411|Abnormality detected in sputum by cytology|sputum cytology positive
Event|Event|Hospital Course|5688,5696|false|false|false|||cytology
Procedure|Laboratory Procedure|Hospital Course|5688,5696|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|cytology
Disorder|Cell or Molecular Dysfunction|Hospital Course|5697,5705|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|5697,5705|false|false|false|||positive
Finding|Classification|Hospital Course|5697,5705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|5697,5705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|5697,5709|false|false|false|C1446409|Positive|positive for
Disorder|Neoplastic Process|Hospital Course|5711,5725|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|5711,5725|false|false|false|||adenocarcinoma
Event|Event|Hospital Course|5728,5735|false|false|false|||Hypoxia
Finding|Finding|Hospital Course|5728,5735|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|Hospital Course|5728,5735|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Event|Event|Hospital Course|5750,5754|false|false|false|||felt
Event|Event|Hospital Course|5763,5774|false|false|false|||combination
Finding|Finding|Hospital Course|5763,5774|false|false|false|C3811910|combination - answer to question|combination
Disorder|Disease or Syndrome|Hospital Course|5779,5804|false|false|false|C0747690|Postobstructive pneumonia|postobstructive pneumonia
Disorder|Disease or Syndrome|Hospital Course|5795,5804|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|5795,5804|false|false|false|||pneumonia
Disorder|Neoplastic Process|Hospital Course|5809,5814|false|false|false|C0027651|Neoplasms|tumor
Event|Event|Hospital Course|5809,5814|false|false|false|||tumor
Finding|Finding|Hospital Course|5809,5814|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|Hospital Course|5809,5814|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Procedure|Diagnostic Procedure|Hospital Course|5809,5821|false|false|false|C1449699|Tumor Burden|tumor burden
Event|Event|Hospital Course|5815,5821|false|false|false|||burden
Finding|Idea or Concept|Hospital Course|5815,5821|false|false|false|C2828008|Burden|burden
Disorder|Neoplastic Process|Hospital Course|5828,5842|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|5828,5842|false|false|false|||adenocarcinoma
Drug|Antibiotic|Hospital Course|5845,5856|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|Hospital Course|5845,5856|false|false|false|||Antibiotics
Event|Event|Hospital Course|5862,5869|false|false|false|||changed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5873,5883|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|5873,5883|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|Hospital Course|5873,5883|false|false|false|||vancomycin
Procedure|Laboratory Procedure|Hospital Course|5873,5883|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|Hospital Course|5886,5898|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|5886,5898|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|5886,5898|false|false|false|||levofloxacin
Drug|Organic Chemical|Hospital Course|5903,5909|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|Hospital Course|5903,5909|false|false|false|C0699678|Flagyl|flagyl
Event|Event|Hospital Course|5903,5909|false|false|false|||flagyl
Event|Event|Hospital Course|5923,5932|false|false|false|||completed
Finding|Idea or Concept|Hospital Course|5938,5941|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5938,5941|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5942,5948|false|false|false|||course
Procedure|Diagnostic Procedure|Hospital Course|5959,5966|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|5962,5966|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|5962,5966|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|5967,5973|false|false|false|||showed
Disorder|Disease or Syndrome|Hospital Course|5974,5980|false|false|false|C0023882|Little's Disease|little
Finding|Finding|Hospital Course|5974,5980|false|false|false|C3889124|Only a Little|little
Finding|Intellectual Product|Hospital Course|5981,5989|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|Hospital Course|5990,6001|false|false|false|||improvement
Finding|Conceptual Entity|Hospital Course|5990,6001|false|false|false|C2986411|Improvement|improvement
Finding|Functional Concept|Hospital Course|6005,6010|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|6011,6016|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|6011,6016|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6018,6022|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|6018,6022|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Hospital Course|6023,6033|false|false|false|||infiltrate
Finding|Functional Concept|Hospital Course|6023,6033|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Hospital Course|6023,6033|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Hospital Course|6023,6033|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Attribute|Clinical Attribute|Hospital Course|6036,6047|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|Hospital Course|6036,6047|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|Hospital Course|6036,6047|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|Hospital Course|6036,6047|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Attribute|Clinical Attribute|Hospital Course|6036,6054|false|false|false|C2598168||Respiratory status
Finding|Finding|Hospital Course|6036,6054|false|false|false|C1998827|Respiratory Status|Respiratory status
Attribute|Clinical Attribute|Hospital Course|6048,6054|false|false|false|C5889824||status
Event|Event|Hospital Course|6048,6054|false|false|false|||status
Finding|Idea or Concept|Hospital Course|6048,6054|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|6064,6071|false|false|false|||tenuous
Finding|Body Substance|Hospital Course|6073,6080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6073,6080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6073,6080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6082,6091|false|false|false|||requiring
Finding|Finding|Hospital Course|6092,6096|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|6092,6096|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|6092,6096|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Phenomenon|Natural Phenomenon or Process|Hospital Course|6097,6101|false|false|false|C0806140|Flow|flow
Event|Event|Hospital Course|6120,6133|false|false|false|||desaturations
Finding|Finding|Hospital Course|6137,6141|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|6137,6141|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|6137,6141|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Activity|Hospital Course|6152,6160|false|false|false|C0441655|Activities|activity
Event|Event|Hospital Course|6152,6160|false|false|false|||activity
Finding|Daily or Recreational Activity|Hospital Course|6152,6160|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Hospital Course|6152,6160|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Hospital Course|6172,6181|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6172,6181|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6172,6181|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6172,6181|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6172,6181|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6185,6196|false|false|false|||requirement
Finding|Functional Concept|Hospital Course|6185,6196|false|false|false|C1514873|Requirement|requirement
Event|Event|Hospital Course|6201,6203|false|false|false|||5L
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6208,6213|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|6208,6213|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|6208,6213|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|6208,6213|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|6208,6213|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|6208,6213|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6214,6221|false|false|false|C1550232|Body Parts - Cannula|cannula
Event|Event|Hospital Course|6214,6221|false|false|false|||cannula
Finding|Body Substance|Hospital Course|6214,6221|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Hospital Course|6214,6221|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Event|Event|Hospital Course|6232,6241|false|false|false|||breathing
Drug|Biologically Active Substance|Hospital Course|6259,6265|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|6259,6265|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|6259,6265|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|6259,6265|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6259,6265|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|6267,6277|false|false|false|||saturation
Phenomenon|Natural Phenomenon or Process|Hospital Course|6267,6277|false|false|false|C0522534|Saturated|saturation
Finding|Finding|Hospital Course|6285,6288|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6285,6288|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Hospital Course|6312,6320|false|false|false|||continue
Event|Event|Hospital Course|6328,6337|false|false|false|||necessary
Finding|Finding|Hospital Course|6347,6351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|6347,6351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|6347,6351|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|6363,6367|false|false|false|||mask
Finding|Gene or Genome|Hospital Course|6363,6367|false|false|false|C1538279;C1555580;C1845191|ANKHD1 gene;STK26 gene;masked - No information|mask
Finding|Idea or Concept|Hospital Course|6363,6367|false|false|false|C1538279;C1555580;C1845191|ANKHD1 gene;STK26 gene;masked - No information|mask
Event|Event|Hospital Course|6375,6379|false|false|false|||used
Event|Event|Hospital Course|6383,6389|false|false|false|||assist
Finding|Social Behavior|Hospital Course|6383,6389|false|false|false|C0018896|Helping Behavior|assist
Procedure|Health Care Activity|Hospital Course|6383,6389|false|false|false|C0557034|Assisting (procedure)|assist
Event|Event|Hospital Course|6396,6407|false|false|false|||oxygenation
Finding|Cell Function|Hospital Course|6396,6407|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Organ or Tissue Function|Hospital Course|6396,6407|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Event|Event|Hospital Course|6411,6417|false|false|false|||needed
Anatomy|Body Location or Region|Hospital Course|6427,6431|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6427,6431|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|Hospital Course|6427,6431|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|Hospital Course|6427,6431|false|false|false|C0740941|Lung Problem|Lung
Finding|Finding|Hospital Course|6427,6439|false|false|false|C0034079||Lung nodules
Event|Event|Hospital Course|6432,6439|false|false|false|||nodules
Disorder|Neoplastic Process|Hospital Course|6458,6467|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|6458,6467|false|false|false|||carcinoma
Procedure|Diagnostic Procedure|Hospital Course|6469,6476|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|6472,6476|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|6472,6476|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6491,6500|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6491,6500|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6491,6500|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|Hospital Course|6491,6508|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|Hospital Course|6501,6508|false|false|false|||nodules
Finding|Body Substance|Hospital Course|6513,6519|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|6513,6519|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Finding|Hospital Course|6513,6528|false|false|false|C0551076|Sputum cytology (finding)|sputum cytology
Procedure|Laboratory Procedure|Hospital Course|6513,6528|false|false|false|C1521752|Sputum Cytology Screening|sputum cytology
Lab|Laboratory or Test Result|Hospital Course|6513,6537|false|false|false|C0580411|Abnormality detected in sputum by cytology|sputum cytology positive
Event|Event|Hospital Course|6520,6528|false|false|false|||cytology
Procedure|Laboratory Procedure|Hospital Course|6520,6528|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|cytology
Disorder|Cell or Molecular Dysfunction|Hospital Course|6529,6537|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|6529,6537|false|false|false|||positive
Finding|Classification|Hospital Course|6529,6537|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6529,6537|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6529,6541|false|false|false|C1446409|Positive|positive for
Disorder|Neoplastic Process|Hospital Course|6543,6557|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|6543,6557|false|false|false|||adenocarcinoma
Event|Event|Hospital Course|6560,6568|false|false|false|||Etiology
Finding|Conceptual Entity|Hospital Course|6560,6568|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|Hospital Course|6560,6568|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Event|Event|Hospital Course|6573,6577|false|false|false|||felt
Event|Event|Hospital Course|6593,6609|false|false|false|||bronchioalveolar
Finding|Functional Concept|Hospital Course|6613,6623|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6624,6631|false|false|false|C0040132|Thyroid Gland|thyroid
Disorder|Disease or Syndrome|Hospital Course|6624,6631|false|false|false|C0040128|Thyroid Diseases|thyroid
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6624,6631|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Hormone|Hospital Course|6624,6631|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6624,6631|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Organic Chemical|Hospital Course|6624,6631|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Pharmacologic Substance|Hospital Course|6624,6631|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Event|Event|Hospital Course|6624,6631|false|false|false|||thyroid
Procedure|Health Care Activity|Hospital Course|6624,6631|false|false|false|C2228489|examination of thyroid|thyroid
Finding|Finding|Hospital Course|6648,6656|false|false|false|C0332149|Possible|possible
Disorder|Neoplastic Process|Hospital Course|6674,6683|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|6674,6683|false|false|false|||carcinoma
Finding|Idea or Concept|Hospital Course|6694,6701|true|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|Hospital Course|6694,6701|true|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|Hospital Course|6694,6701|true|false|false|C1979801|Routine coag|routine
Disorder|Neoplastic Process|Hospital Course|6702,6708|true|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Diagnostic Procedure|Hospital Course|6702,6718|true|false|false|C0199230|Screening for cancer|cancer screening
Event|Event|Hospital Course|6709,6718|true|false|false|||screening
Finding|Finding|Hospital Course|6709,6718|true|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|Hospital Course|6709,6718|true|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|Hospital Course|6709,6718|true|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|Hospital Course|6709,6718|true|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|Hospital Course|6709,6718|true|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Anatomy|Tissue|Hospital Course|6743,6749|true|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Hospital Course|6743,6749|true|false|false|C1547928|Tissue Specimen Code|tissue
Finding|Finding|Hospital Course|6743,6759|true|false|false|C1546905|Tissue diagnosis|tissue diagnosis
Attribute|Clinical Attribute|Hospital Course|6750,6759|true|false|false|C0945731||diagnosis
Event|Event|Hospital Course|6750,6759|true|false|false|||diagnosis
Finding|Classification|Hospital Course|6750,6759|true|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|6750,6759|true|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6750,6759|true|false|false|C0011900|Diagnosis|diagnosis
Finding|Body Substance|Hospital Course|6788,6795|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6788,6795|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6788,6795|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|6798,6802|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|6798,6802|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|6798,6802|true|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Biologically Active Substance|Hospital Course|6803,6809|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|6803,6809|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|6803,6809|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6803,6809|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|6810,6821|false|false|false|||requirement
Finding|Functional Concept|Hospital Course|6810,6821|false|false|false|C1514873|Requirement|requirement
Event|Event|Hospital Course|6826,6841|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|6826,6841|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|6826,6841|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6826,6841|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Drug|Organic Chemical|Hospital Course|6848,6854|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|6848,6854|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|6848,6854|false|false|false|||plavix
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6855,6858|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Enzyme|Hospital Course|6855,6858|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Organic Chemical|Hospital Course|6855,6858|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Pharmacologic Substance|Hospital Course|6855,6858|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Event|Event|Hospital Course|6855,6858|false|false|false|||asa
Finding|Gene or Genome|Hospital Course|6855,6858|false|false|false|C1412553|ARSA gene|asa
Finding|Mental Process|Hospital Course|6866,6873|false|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|6888,6897|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|6888,6897|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6888,6897|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Body Substance|Hospital Course|6910,6917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6910,6917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6910,6917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6931,6938|true|false|false|||imaging
Finding|Finding|Hospital Course|6931,6938|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|6931,6938|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Anatomy|Body Location or Region|Hospital Course|6946,6950|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6946,6950|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|6946,6950|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6946,6950|true|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|6952,6959|true|false|false|||staging
Finding|Functional Concept|Hospital Course|6952,6959|true|false|false|C0332305|With staging|staging
Event|Event|Hospital Course|6969,6971|false|false|false|||CT
Disorder|Virus|Hospital Course|6983,6987|false|false|false|C4697913|Venezuelan equine encephalitis virus subtype IIIA|IIIa
Event|Event|Hospital Course|6983,6987|false|false|false|||IIIa
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6993,7002|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6993,7002|true|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6993,7002|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|Hospital Course|6993,7010|true|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|Hospital Course|7003,7010|true|false|false|||nodules
Anatomy|Body Location or Region|Hospital Course|7019,7023|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7019,7023|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|7019,7023|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|7019,7023|true|false|false|C0740941|Lung Problem|lung
Attribute|Clinical Attribute|Hospital Course|7048,7054|true|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7055,7058|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|7055,7058|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Hospital Course|7055,7058|true|false|false|||LAD
Finding|Gene or Genome|Hospital Course|7055,7058|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Neoplastic Process|Hospital Course|7062,7072|true|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastasis
Event|Event|Hospital Course|7062,7072|true|false|false|||metastasis
Finding|Finding|Hospital Course|7062,7072|true|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Finding|Pathologic Function|Hospital Course|7062,7072|true|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Event|Event|Hospital Course|7083,7090|false|false|false|||therapy
Finding|Finding|Hospital Course|7083,7090|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|7083,7090|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7083,7090|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Hospital Course|7097,7103|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Drug|Chemical Viewed Functionally|Hospital Course|7104,7109|false|false|false|C0450442;C1254351|Agent;Pharmacologic Substance|agent
Drug|Pharmacologic Substance|Hospital Course|7104,7109|false|false|false|C0450442;C1254351|Agent;Pharmacologic Substance|agent
Finding|Functional Concept|Hospital Course|7104,7109|false|false|false|C1521826;C1551364;C4763809|GDC Therapeutic Agent Terminology;Protocol Agent;agent - RoleClass|agent
Finding|Intellectual Product|Hospital Course|7104,7109|false|false|false|C1521826;C1551364;C4763809|GDC Therapeutic Agent Terminology;Protocol Agent;agent - RoleClass|agent
Event|Event|Hospital Course|7110,7122|false|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|7110,7122|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7110,7122|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Hospital Course|7127,7136|false|false|false|||initiated
Drug|Organic Chemical|Hospital Course|7150,7160|false|false|false|C0210657|pemetrexed|Pemetrexed
Drug|Pharmacologic Substance|Hospital Course|7150,7160|false|false|false|C0210657|pemetrexed|Pemetrexed
Event|Event|Hospital Course|7150,7160|false|false|false|||Pemetrexed
Event|Event|Hospital Course|7167,7176|false|false|false|||tolerated
Finding|Finding|Hospital Course|7182,7186|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|7193,7201|false|false|false|||received
Drug|Organic Chemical|Hospital Course|7203,7216|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|Hospital Course|7203,7216|false|false|false|C0011777|dexamethasone|dexamethasone
Event|Event|Hospital Course|7203,7216|false|false|false|||dexamethasone
Disorder|Disease or Syndrome|Hospital Course|7235,7239|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|Hospital Course|7235,7239|false|false|false|||rash
Finding|Pathologic Function|Hospital Course|7235,7239|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|Hospital Course|7235,7239|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Intellectual Product|Hospital Course|7247,7254|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|7247,7254|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|7247,7274|false|false|false|C0403447|Chronic Kidney Insufficiency|Chronic renal insufficiency
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7255,7260|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|7255,7260|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|7255,7274|false|false|false|C0035078;C1565489|Kidney Failure;Renal Insufficiency|renal insufficiency
Event|Event|Hospital Course|7261,7274|false|false|false|||insufficiency
Finding|Functional Concept|Hospital Course|7261,7274|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Body Substance|Hospital Course|7277,7284|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7277,7284|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7277,7284|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7290,7293|false|false|false|||GFR
Finding|Gene or Genome|Hospital Course|7290,7293|false|false|false|C1424601|RAPGEF5 gene|GFR
Attribute|Clinical Attribute|Hospital Course|7300,7311|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7300,7311|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7300,7311|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7300,7311|false|false|false|C4284232|Medications|Medications
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7335,7340|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|7335,7340|false|false|false|C0042075|Urologic Diseases|renal
Finding|Organ or Tissue Function|Hospital Course|7335,7349|false|false|false|C0232804|Renal function|renal function
Procedure|Laboratory Procedure|Hospital Course|7335,7349|false|false|false|C0022662|Kidney Function Tests|renal function
Event|Event|Hospital Course|7341,7349|false|false|false|||function
Finding|Finding|Hospital Course|7341,7349|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|7341,7349|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|7341,7349|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|7341,7349|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Hospital Course|7365,7373|false|false|false|||followed
Event|Event|Hospital Course|7384,7391|false|false|false|||treated
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7414,7422|false|false|false|C0699252|Mucomyst|mucomyst
Drug|Pharmacologic Substance|Hospital Course|7414,7422|false|false|false|C0699252|Mucomyst|mucomyst
Event|Event|Hospital Course|7414,7422|false|false|false|||mucomyst
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|7442,7453|false|false|false|C4072741|IV contrast|IV contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|7445,7453|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Hospital Course|7445,7453|false|false|false|||contrast
Event|Event|Hospital Course|7454,7458|false|false|false|||dose
Drug|Biologically Active Substance|Hospital Course|7461,7471|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|7461,7471|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|7461,7471|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|7461,7471|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|7461,7471|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|7472,7480|false|false|false|||remained
Event|Event|Hospital Course|7481,7487|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|7481,7487|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|7502,7514|false|false|false|||Hyperkalemia
Finding|Finding|Hospital Course|7502,7514|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Finding|Body Substance|Hospital Course|7521,7528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7521,7528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7521,7528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7540,7552|false|false|false|||hyperkalemic
Finding|Idea or Concept|Hospital Course|7557,7560|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7557,7560|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|7571,7580|true|false|false|||discharge
Finding|Body Substance|Hospital Course|7571,7580|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7571,7580|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7571,7580|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7571,7580|true|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|7596,7599|true|false|false|||EKG
Finding|Intellectual Product|Hospital Course|7596,7599|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|7596,7599|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|7600,7607|true|false|false|||changes
Finding|Functional Concept|Hospital Course|7600,7607|true|false|false|C0392747|Changing|changes
Drug|Organic Chemical|Hospital Course|7639,7649|false|false|false|C0124498|Kayexalate|kayexalate
Drug|Pharmacologic Substance|Hospital Course|7639,7649|false|false|false|C0124498|Kayexalate|kayexalate
Event|Event|Hospital Course|7639,7649|false|false|false|||kayexalate
Drug|Inorganic Chemical|Hospital Course|7652,7664|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Drug|Pharmacologic Substance|Hospital Course|7652,7664|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Event|Event|Hospital Course|7652,7664|false|false|false|||Electrolytes
Event|Event|Hospital Course|7675,7682|false|false|false|||checked
Event|Event|Hospital Course|7696,7702|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|7696,7702|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|7718,7722|false|false|false|||ACEI
Event|Event|Hospital Course|7732,7739|false|false|false|||stopped
Disorder|Disease or Syndrome|Hospital Course|7744,7747|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|7744,7747|false|false|false|||HTN
Event|Event|Hospital Course|7758,7770|false|false|false|||normotensive
Event|Event|Hospital Course|7774,7778|false|false|false|||ACEI
Event|Event|Hospital Course|7785,7792|false|false|false|||blocker
Attribute|Clinical Attribute|Hospital Course|7799,7810|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7799,7810|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7799,7810|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7799,7810|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|7799,7823|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|7814,7823|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|7814,7823|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|7827,7838|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|7827,7838|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|7840,7846|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|7840,7846|false|false|false|C0633084|Plavix|Plavix
Drug|Biomedical or Dental Material|Hospital Course|7854,7860|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|7872,7881|false|false|false|C1142985|ezetimibe|Ezetimibe
Drug|Pharmacologic Substance|Hospital Course|7872,7881|false|false|false|C1142985|ezetimibe|Ezetimibe
Drug|Pharmacologic Substance|Hospital Course|7872,7893|false|false|false|C1532737|ezetimibe / simvastatin|Ezetimibe-Simvastatin
Drug|Organic Chemical|Hospital Course|7882,7893|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|7882,7893|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|Hospital Course|7895,7902|false|false|false|C1527845|Vytorin|Vytorin
Drug|Pharmacologic Substance|Hospital Course|7895,7902|false|false|false|C1527845|Vytorin|Vytorin
Drug|Organic Chemical|Hospital Course|7937,7947|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|Hospital Course|7937,7947|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Organic Chemical|Hospital Course|7967,7980|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|7967,7980|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Biomedical or Dental Material|Hospital Course|7993,7998|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|7993,7998|false|false|false|||Patch
Finding|Finding|Hospital Course|7993,7998|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Biomedical or Dental Material|Hospital Course|8007,8012|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|Hospital Course|8007,8012|false|false|false|||patch
Finding|Finding|Hospital Course|8007,8012|false|false|false|C0332461|Plaque (lesion)|patch
Finding|Intellectual Product|Hospital Course|8013,8017|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|8013,8023|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|8020,8023|false|false|false|||day
Finding|Idea or Concept|Hospital Course|8020,8023|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8020,8023|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|8042,8052|true|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|sublingual
Finding|Functional Concept|Hospital Course|8042,8052|true|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|sublingual
Finding|Gene or Genome|Hospital Course|8058,8061|true|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8072,8076|true|false|false|||used
Event|Event|Hospital Course|8086,8091|true|false|false|||prior
Drug|Organic Chemical|Hospital Course|8104,8115|false|false|false|C0033497|propranolol|Propranolol
Drug|Pharmacologic Substance|Hospital Course|8104,8115|false|false|false|C0033497|propranolol|Propranolol
Drug|Biomedical or Dental Material|Hospital Course|8122,8128|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|8132,8136|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|8132,8142|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|8139,8142|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8139,8142|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|8155,8167|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|8155,8167|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|8155,8167|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Event|Event|Hospital Course|8170,8179|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8170,8179|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8170,8179|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8170,8179|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8170,8179|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8170,8191|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8170,8191|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8180,8191|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8180,8191|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8180,8191|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|8193,8201|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8193,8201|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|8193,8206|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|8202,8206|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|8202,8206|false|false|false|||Care
Finding|Finding|Hospital Course|8202,8206|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|8202,8206|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|8209,8217|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|8209,8217|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|8225,8234|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8225,8234|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8225,8234|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8225,8234|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8225,8234|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8225,8244|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|8235,8244|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|8235,8244|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|8235,8244|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8235,8244|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8235,8244|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Hospital Course|8255,8267|false|false|false|C0520886|ST segment elevation (finding)|ST elevation
Disorder|Disease or Syndrome|Hospital Course|8255,8289|false|false|false|C1536220|ST segment elevation myocardial infarction|ST elevation myocardial infarction
Event|Event|Hospital Course|8258,8267|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8258,8267|false|false|false|C0439775|Elevation procedure|elevation
Anatomy|Tissue|Hospital Course|8268,8278|false|false|false|C0027061|Myocardium|myocardial
Attribute|Clinical Attribute|Hospital Course|8268,8289|false|false|false|C2926063||myocardial infarction
Disorder|Disease or Syndrome|Hospital Course|8268,8289|false|false|false|C0027051|Myocardial Infarction|myocardial infarction
Event|Event|Hospital Course|8279,8289|false|false|false|||infarction
Finding|Pathologic Function|Hospital Course|8279,8289|false|false|false|C0021308|Infarction|infarction
Event|Event|Hospital Course|8290,8298|false|false|false|||Presumed
Disorder|Neoplastic Process|Hospital Course|8316,8325|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|8316,8325|false|false|false|||carcinoma
Event|Event|Discharge Condition|8350,8356|false|false|false|||stable
Finding|Intellectual Product|Discharge Condition|8350,8356|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Biologically Active Substance|Discharge Condition|8366,8372|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Condition|8366,8372|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Condition|8366,8372|false|false|false|C0030054|oxygen|oxygen
Event|Event|Discharge Condition|8366,8372|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|8366,8372|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Condition|8373,8384|false|false|false|||requirement
Finding|Functional Concept|Discharge Condition|8373,8384|false|false|false|C1514873|Requirement|requirement
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|8392,8395|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|Discharge Condition|8392,8395|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|Discharge Condition|8392,8395|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|Discharge Condition|8392,8395|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Finding|Discharge Condition|8403,8406|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Condition|8403,8406|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Discharge Instructions|8447,8455|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|8463,8471|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|8476,8481|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|8476,8481|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Discharge Instructions|8476,8490|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|Discharge Instructions|8482,8490|false|false|false|||pressure
Finding|Finding|Discharge Instructions|8482,8490|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|8482,8490|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|8482,8490|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|8482,8490|false|false|false|C0033095||pressure
Event|Event|Discharge Instructions|8495,8500|false|false|false|||found
Finding|Finding|Discharge Instructions|8495,8500|false|false|false|C0150312|Present|found
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8512,8517|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8512,8517|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8512,8517|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|8512,8524|false|false|false|C0027051|Myocardial Infarction|heart attack
Event|Event|Discharge Instructions|8518,8524|false|false|false|||attack
Finding|Finding|Discharge Instructions|8518,8524|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Discharge Instructions|8518,8524|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8537,8544|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Discharge Instructions|8537,8544|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|Discharge Instructions|8537,8560|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|Discharge Instructions|8537,8560|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|Discharge Instructions|8537,8560|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|Discharge Instructions|8537,8560|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|Discharge Instructions|8545,8560|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8545,8560|false|false|false|C0007430|Catheterization|catheterization
Drug|Inorganic Chemical|Discharge Instructions|8577,8582|false|false|false|C0025552|Metals|metal
Event|Event|Discharge Instructions|8583,8588|false|false|false|||stent
Event|Event|Discharge Instructions|8589,8595|false|false|false|||placed
Event|Event|Discharge Instructions|8623,8630|false|false|false|||trouble
Attribute|Clinical Attribute|Discharge Instructions|8632,8641|false|false|false|C5885990||breathing
Event|Event|Discharge Instructions|8632,8641|false|false|false|||breathing
Finding|Finding|Discharge Instructions|8632,8641|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|8632,8641|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|8632,8641|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|8632,8641|false|false|false|C1160636|respiratory system process|breathing
Event|Event|Discharge Instructions|8652,8656|false|false|false|||scan
Procedure|Diagnostic Procedure|Discharge Instructions|8652,8656|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Discharge Instructions|8662,8668|false|false|false|||showed
Event|Event|Discharge Instructions|8674,8681|false|false|false|||nodules
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8690,8695|false|false|false|C0024109|Lung|lungs
Finding|Body Substance|Discharge Instructions|8701,8707|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Discharge Instructions|8701,8707|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Body Substance|Discharge Instructions|8701,8714|false|false|false|C0444159|Sputum specimen|sputum sample
Drug|Substance|Discharge Instructions|8708,8714|false|false|false|C0370003|Specimen|sample
Event|Event|Discharge Instructions|8708,8714|false|false|false|||sample
Finding|Body Substance|Discharge Instructions|8708,8714|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Finding|Intellectual Product|Discharge Instructions|8708,8714|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Event|Event|Discharge Instructions|8719,8723|false|false|false|||sent
Anatomy|Cell|Discharge Instructions|8728,8743|false|false|false|C0334227|Tumor cells, malignant|malignant cells
Anatomy|Cell|Discharge Instructions|8738,8743|false|false|false|C0007634|Cells|cells
Event|Event|Discharge Instructions|8749,8753|false|false|false|||seen
Event|Event|Discharge Instructions|8765,8772|false|false|false|||thought
Anatomy|Body Location or Region|Discharge Instructions|8796,8800|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8796,8800|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|8796,8800|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|8796,8800|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Discharge Instructions|8796,8807|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Discharge Instructions|8801,8807|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Discharge Instructions|8801,8807|false|false|false|||cancer
Event|Event|Discharge Instructions|8823,8830|false|false|false|||treated
Event|Event|Discharge Instructions|8840,8844|false|false|false|||dose
Event|Event|Discharge Instructions|8848,8860|false|false|false|||chemotherapy
Finding|Functional Concept|Discharge Instructions|8848,8860|false|false|true|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8848,8860|false|false|true|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Discharge Instructions|8880,8886|false|false|false|||follow
Event|Event|Discharge Instructions|8906,8915|false|false|false|||determine
Event|Event|Discharge Instructions|8928,8937|false|false|false|||treatment
Finding|Conceptual Entity|Discharge Instructions|8928,8937|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Discharge Instructions|8928,8937|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Discharge Instructions|8928,8937|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8928,8937|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Discharge Instructions|8946,8952|false|false|false|||needed
Event|Event|Discharge Instructions|8985,8989|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|8996,9002|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|8996,9002|false|false|false|||weight
Finding|Finding|Discharge Instructions|8996,9002|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|8996,9002|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|8996,9002|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|9003,9007|false|false|false|||goes
Procedure|Laboratory Procedure|Discharge Instructions|9024,9027|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|9044,9051|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|9044,9051|false|false|false|C0392747|Changing|changes
Event|Event|Discharge Instructions|9057,9061|false|false|false|||made
Attribute|Clinical Attribute|Discharge Instructions|9070,9081|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9070,9081|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9070,9081|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9070,9081|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9095,9102|false|false|false|||started
Drug|Organic Chemical|Discharge Instructions|9106,9112|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Discharge Instructions|9106,9112|false|false|false|C0633084|Plavix|plavix
Event|Event|Discharge Instructions|9106,9112|false|false|false|||plavix
Drug|Pharmacologic Substance|Discharge Instructions|9116,9126|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|9116,9126|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|9116,9126|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|9130,9134|false|false|false|||thin
Disorder|Disease or Syndrome|Discharge Instructions|9140,9145|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|9140,9145|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|9140,9145|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|9157,9161|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|9167,9177|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|9167,9177|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|9167,9177|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|9184,9189|false|false|false|||month
Finding|Idea or Concept|Discharge Instructions|9184,9189|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Discharge Instructions|9184,9189|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Drug|Food|Discharge Instructions|9193,9199|true|false|false|C0218063|Ensure (product)|ensure
Event|Event|Discharge Instructions|9193,9199|true|false|false|||ensure
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9211,9216|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|9211,9216|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|9211,9216|true|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Discharge Instructions|9217,9222|true|false|false|||stent
Event|Event|Discharge Instructions|9232,9238|true|false|false|||become
Event|Event|Discharge Instructions|9239,9246|true|false|false|||blocked
Finding|Finding|Discharge Instructions|9239,9246|true|true|false|C0028778;C0332206|Blocking;Obstruction|blocked
Finding|Functional Concept|Discharge Instructions|9239,9246|true|true|false|C0028778;C0332206|Blocking;Obstruction|blocked
Procedure|Health Care Activity|Discharge Instructions|9251,9259|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9260,9272|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9260,9272|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9260,9272|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

