 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
MEDICINE|155,163
<EOL>|163,164
<EOL>|165,166
Allergies|166,175
:|175,176
<EOL>|177,178
Codeine|178,185
/|186,187
Augmentin|188,197
/|198,199
Topamax|200,207
<EOL>|207,208
<EOL>|209,210
Attending|210,219
:|219,220
_|221,222
_|222,223
_|223,224
.|224,225
<EOL>|225,226
<EOL>|227,228
Chief|228,233
Complaint|234,243
:|243,244
<EOL>|244,245
RLE|245,248
pain|249,253
and|254,257
swelling|258,266
<EOL>|266,267
<EOL>|268,269
Major|269,274
Surgical|275,283
or|284,286
Invasive|287,295
Procedure|296,305
:|305,306
<EOL>|306,307
Ultrasound|307,317
guided|318,324
steroid|325,332
injection|333,342
of|343,345
the|346,349
right|350,355
trochanteric|356,368
<EOL>|369,370
bursa|370,375
(|376,377
right|377,382
hip|383,386
)|386,387
<EOL>|387,388
<EOL>|388,389
<EOL>|390,391
History|391,398
of|399,401
Present|402,409
Illness|410,417
:|417,418
<EOL>|418,419
This|419,423
is|424,426
a|427,428
_|429,430
_|430,431
_|431,432
woman|433,438
with|439,443
a|444,445
history|446,453
of|454,456
breast|457,463
cancer|464,470
with|471,475
<EOL>|475,476
BRCA1|476,481
gene|482,486
mutation|487,495
,|495,496
COPD|497,501
,|501,502
cerebral|503,511
aneurysm|512,520
,|520,521
sleep|522,527
apnea|528,533
,|533,534
<EOL>|534,535
depression|535,545
,|545,546
hyperlipidemia|547,561
,|561,562
antiphospholipid|563,579
syndrome|580,588
with|589,593
hx|594,596
<EOL>|596,597
DVT|597,600
/|600,601
PE|601,603
_|604,605
_|605,606
_|606,607
ago|608,611
on|612,614
warfarin|615,623
who|624,627
presents|628,636
for|637,640
evaluation|641,651
of|652,654
severe|655,661
<EOL>|661,662
right|662,667
lower|668,673
extremity|674,683
pain|684,688
.|688,689
<EOL>|689,690
<EOL>|690,691
She|691,694
was|695,698
just|699,703
admitted|704,712
to|713,715
the|716,719
hospital|720,728
for|729,732
lumpectomy|733,743
<EOL>|743,744
(|744,745
infiltrating|745,757
ductal|758,764
carcinoma|765,774
of|775,777
left|778,782
breast|783,789
)|789,790
and|791,794
sentinel|795,803
<EOL>|804,805
lymph|805,810
<EOL>|810,811
node|811,815
biopsy|816,822
on|823,825
_|826,827
_|827,828
_|828,829
,|829,830
complicated|831,842
by|843,845
hematoma|846,854
status|855,861
post|862,866
<EOL>|866,867
evacuation|867,877
on|878,880
_|881,882
_|882,883
_|883,884
.|884,885
Prior|886,891
to|892,894
these|895,900
procedures|901,911
,|911,912
she|913,916
had|917,920
<EOL>|921,922
severe|922,928
<EOL>|928,929
right|929,934
lower|935,940
extremity|941,950
pain|951,955
similar|956,963
to|964,966
today|967,972
and|973,976
underwent|977,986
a|987,988
DVT|989,992
<EOL>|992,993
ultrasound|993,1003
on|1004,1006
_|1007,1008
_|1008,1009
_|1009,1010
which|1011,1016
was|1017,1020
negative|1021,1029
.|1029,1030
Her|1031,1034
anticoagulation|1035,1050
was|1051,1054
<EOL>|1054,1055
held|1055,1059
in|1060,1062
the|1063,1066
hospital|1067,1075
due|1076,1079
to|1080,1082
the|1083,1086
hematoma|1087,1095
,|1095,1096
and|1097,1100
she|1101,1104
had|1105,1108
DVT|1109,1112
<EOL>|1112,1113
prophylaxis|1113,1124
with|1125,1129
pneumoboots|1130,1141
.|1141,1142
<EOL>|1142,1143
<EOL>|1143,1144
During|1144,1150
her|1151,1154
postoperative|1155,1168
hematoma|1169,1177
her|1178,1181
anticoagulation|1182,1197
was|1198,1201
held|1202,1206
.|1206,1207
<EOL>|1207,1208
She|1208,1211
did|1212,1215
not|1216,1219
have|1220,1224
extremity|1225,1234
pain|1235,1239
during|1240,1246
her|1247,1250
time|1251,1255
in|1256,1258
the|1259,1262
hospital|1263,1271
.|1271,1272
<EOL>|1272,1273
However|1273,1280
,|1280,1281
upon|1282,1286
returning|1287,1296
home|1297,1301
,|1301,1302
she|1303,1306
developed|1307,1316
severe|1317,1323
pain|1324,1328
which|1329,1334
<EOL>|1335,1336
she|1336,1339
<EOL>|1339,1340
describes|1340,1349
as|1350,1352
cramps|1353,1359
in|1360,1362
her|1363,1366
mid|1367,1370
calf|1371,1375
on|1376,1378
the|1379,1382
right|1383,1388
.|1388,1389
She|1390,1393
also|1394,1398
has|1399,1402
<EOL>|1402,1403
pain|1403,1407
that|1408,1412
intermittently|1413,1427
occurs|1428,1434
in|1435,1437
the|1438,1441
right|1442,1447
thigh|1448,1453
which|1454,1459
she|1460,1463
<EOL>|1463,1464
describes|1464,1473
as|1474,1476
spasms|1477,1483
.|1483,1484
She|1485,1488
has|1489,1492
not|1493,1496
had|1497,1500
numbness|1501,1509
,|1509,1510
tingling|1511,1519
,|1519,1520
or|1521,1523
<EOL>|1523,1524
weakness|1524,1532
on|1533,1535
that|1536,1540
side|1541,1545
.|1545,1546
She|1547,1550
was|1551,1554
seen|1555,1559
in|1560,1562
breast|1563,1569
clinic|1570,1576
today|1577,1582
where|1583,1588
<EOL>|1588,1589
she|1589,1592
complained|1593,1603
of|1604,1606
this|1607,1611
pain|1612,1616
,|1616,1617
and|1618,1621
was|1622,1625
referred|1626,1634
to|1635,1637
the|1638,1641
ED|1642,1644
for|1645,1648
<EOL>|1648,1649
further|1649,1656
evaluation|1657,1667
.|1667,1668
She|1669,1672
initially|1673,1682
triggered|1683,1692
as|1693,1695
a|1696,1697
pulseless|1698,1707
<EOL>|1707,1708
extremity|1708,1717
because|1718,1725
of|1726,1728
nonpalpable|1729,1740
pulses|1741,1747
in|1748,1750
the|1751,1754
right|1755,1760
foot|1761,1765
.|1765,1766
She|1767,1770
<EOL>|1770,1771
has|1771,1774
been|1775,1779
taking|1780,1786
Tylenol|1787,1794
as|1795,1797
well|1798,1802
as|1803,1805
tramadol|1806,1814
with|1815,1819
minimal|1820,1827
pain|1828,1832
<EOL>|1832,1833
relief|1833,1839
.|1839,1840
<EOL>|1841,1842
<EOL>|1842,1843
Of|1843,1845
note|1846,1850
,|1850,1851
she|1852,1855
resumed|1856,1863
her|1864,1867
warfarin|1868,1876
without|1877,1884
any|1885,1888
enoxaparin|1889,1899
bridge|1900,1906
<EOL>|1906,1907
this|1907,1911
past|1912,1916
_|1917,1918
_|1918,1919
_|1919,1920
.|1920,1921
She|1922,1925
has|1926,1929
been|1930,1934
wearing|1935,1942
compression|1943,1954
stockings|1955,1964
and|1965,1968
<EOL>|1968,1969
elevating|1969,1978
her|1979,1982
leg|1983,1986
in|1987,1989
an|1990,1992
attempt|1993,2000
to|2001,2003
relieve|2004,2011
the|2012,2015
pain|2016,2020
.|2020,2021
<EOL>|2022,2023
<EOL>|2023,2024
In|2024,2026
the|2027,2030
ED|2031,2033
,|2033,2034
initial|2035,2042
vitals|2043,2049
:|2049,2050
<EOL>|2053,2054
T|2054,2055
98.7|2056,2060
HR|2062,2064
85|2065,2067
BP|2069,2071
175|2072,2075
/|2075,2076
77|2076,2078
RR|2080,2082
20|2083,2085
O2|2087,2089
Sat|2090,2093
98|2094,2096
%|2096,2097
RA|2098,2100
<EOL>|2101,2102
<EOL>|2102,2103
-|2103,2104
Exam|2105,2109
notable|2110,2117
for|2118,2121
:|2121,2122
<EOL>|2124,2125
Right|2125,2130
lower|2131,2136
extremity|2137,2146
with|2147,2151
dopplerable|2152,2163
pulses|2164,2170
,|2170,2171
palpable|2172,2180
pulses|2181,2187
<EOL>|2188,2189
in|2189,2191
<EOL>|2191,2192
the|2192,2195
left|2196,2200
lower|2201,2206
extremity|2207,2216
.|2216,2217
The|2218,2221
right|2222,2227
lower|2228,2233
extremity|2234,2243
is|2244,2246
warm|2247,2251
.|2251,2252
<EOL>|2252,2253
There|2253,2258
is|2259,2261
tenderness|2262,2272
to|2273,2275
palpation|2276,2285
of|2286,2288
the|2289,2292
right|2293,2298
calf|2299,2303
.|2303,2304
Tenderness|2305,2315
<EOL>|2316,2317
to|2317,2319
<EOL>|2319,2320
palpation|2320,2329
of|2330,2332
the|2333,2336
right|2337,2342
thigh|2343,2348
.|2348,2349
<EOL>|2349,2350
<EOL>|2350,2351
-|2351,2352
Labs|2353,2357
notable|2358,2365
for|2366,2369
:|2369,2370
<EOL>|2372,2373
Chem|2373,2377
panel|2378,2383
:|2383,2384
Unremarkable|2385,2397
with|2398,2402
Cr|2403,2405
0.8|2406,2409
<EOL>|2409,2410
CK|2410,2412
67|2413,2415
<EOL>|2415,2416
CBC|2416,2419
:|2419,2420
WBC|2421,2424
5.6|2425,2428
,|2428,2429
Hgb|2430,2433
10.8|2434,2438
with|2439,2443
MCV|2444,2447
93|2448,2450
,|2450,2451
Plt|2452,2455
264|2456,2459
<EOL>|2459,2460
Coags|2460,2465
:|2465,2466
_|2467,2468
_|2468,2469
_|2469,2470
14.8|2471,2475
,|2475,2476
PTT|2477,2480
28.2|2481,2485
,|2485,2486
INR|2487,2490
1.4|2491,2494
<EOL>|2494,2495
Lactate|2495,2502
1.1|2503,2506
<EOL>|2506,2507
UA|2507,2509
:|2509,2510
Mod|2511,2514
Leuk|2515,2519
,|2519,2520
few|2521,2524
bacteria|2525,2533
<EOL>|2533,2534
<EOL>|2534,2535
-|2535,2536
Imaging|2537,2544
notable|2545,2552
for|2553,2556
:|2556,2557
<EOL>|2559,2560
<EOL>|2560,2561
RLE|2561,2564
Ultrasound|2565,2575
_|2576,2577
_|2577,2578
_|2578,2579
<EOL>|2579,2580
Right|2580,2585
calf|2586,2590
veins|2591,2596
not|2597,2600
visualized|2601,2611
.|2611,2612
Otherwise|2613,2622
,|2622,2623
no|2624,2626
evidence|2627,2635
of|2636,2638
deep|2639,2643
<EOL>|2643,2644
venous|2644,2650
<EOL>|2650,2651
thrombosis|2651,2661
in|2662,2664
the|2665,2668
right|2669,2674
lower|2675,2680
extremity|2681,2690
veins|2691,2696
.|2696,2697
<EOL>|2697,2698
<EOL>|2698,2699
CT|2699,2701
Lower|2702,2707
Extremity|2708,2717
Right|2718,2723
_|2724,2725
_|2725,2726
_|2726,2727
<EOL>|2727,2728
Unremarkable|2728,2740
contrast|2741,2749
enhanced|2750,2758
CT|2759,2761
of|2762,2764
the|2765,2768
right|2769,2774
calf|2775,2779
with|2780,2784
a|2785,2786
two|2787,2790
<EOL>|2790,2791
vessel|2791,2797
runoff|2798,2804
to|2805,2807
the|2808,2811
foot|2812,2816
.|2816,2817
<EOL>|2817,2818
The|2818,2821
veins|2822,2827
of|2828,2830
the|2831,2834
lower|2835,2840
extremity|2841,2850
are|2851,2854
not|2855,2858
opacified|2859,2868
therefore|2869,2878
<EOL>|2878,2879
can|2879,2882
not|2882,2885
be|2886,2888
<EOL>|2888,2889
assessed|2889,2897
for|2898,2901
patency|2902,2909
.|2909,2910
Consider|2911,2919
repeat|2920,2926
ultrasound|2927,2937
to|2938,2940
more|2941,2945
fully|2946,2951
<EOL>|2951,2952
evaluate|2952,2960
.|2960,2961
<EOL>|2961,2962
No|2962,2964
focal|2965,2970
collection|2971,2981
or|2982,2984
obvious|2985,2992
muscular|2993,3001
abnormality|3002,3013
identified|3014,3024
<EOL>|3025,3026
by|3026,3028
<EOL>|3028,3029
CT|3029,3031
.|3031,3032
<EOL>|3032,3033
<EOL>|3033,3034
-|3034,3035
Pt|3036,3038
given|3039,3044
:|3044,3045
<EOL>|3047,3048
IV|3048,3050
Morphine|3051,3059
4mg|3060,3063
<EOL>|3063,3064
IV|3064,3066
APAP|3067,3071
1g|3072,3074
<EOL>|3074,3075
IV|3075,3077
NS|3078,3080
<EOL>|3080,3081
IV|3081,3083
Dilaudid|3084,3092
5|3093,3094
mg|3095,3097
total|3098,3103
(|3104,3105
1mg|3105,3108
x|3109,3110
5|3111,3112
)|3112,3113
<EOL>|3113,3114
Warfarin|3114,3122
7.5|3123,3126
mg|3126,3128
<EOL>|3128,3129
Atorvastatin|3129,3141
40mg|3142,3146
<EOL>|3146,3147
Omeprazole|3147,3157
20mg|3158,3162
<EOL>|3162,3163
<EOL>|3163,3164
Surgery|3164,3171
was|3172,3175
consulted|3176,3185
:|3185,3186
Recommend|3187,3196
vascular|3197,3205
surgery|3206,3213
consult|3214,3221
for|3222,3225
<EOL>|3225,3226
possible|3226,3234
dvt|3235,3238
with|3239,3243
history|3244,3251
of|3252,3254
multiple|3255,3263
vein|3264,3268
stripping|3269,3278
procedures|3279,3289
<EOL>|3289,3290
and|3290,3293
DVTs|3294,3298
.|3298,3299
Also|3300,3304
recommend|3305,3314
admission|3315,3324
to|3325,3327
medicine|3328,3336
for|3337,3340
pain|3341,3345
control|3346,3353
.|3353,3354
<EOL>|3355,3356
<EOL>|3356,3357
<EOL>|3357,3358
Vascular|3358,3366
surgery|3367,3374
was|3375,3378
consulted|3379,3388
:|3388,3389
There|3390,3395
is|3396,3398
no|3399,3401
clear|3402,3407
vascular|3408,3416
<EOL>|3416,3417
etiology|3417,3425
for|3426,3429
her|3430,3433
pain|3434,3438
.|3438,3439
<EOL>|3439,3440
<EOL>|3440,3441
-|3441,3442
Vitals|3443,3449
prior|3450,3455
to|3456,3458
transfer|3459,3467
:|3467,3468
<EOL>|3471,3472
T|3472,3473
98.3|3474,3478
HR|3480,3482
83|3483,3485
BP|3487,3489
140|3490,3493
/|3493,3494
55|3494,3496
RR|3498,3500
20|3501,3503
O2|3505,3507
Sat|3508,3511
100|3512,3515
%|3515,3516
RA|3517,3519
<EOL>|3520,3521
<EOL>|3521,3522
Upon|3522,3526
arrival|3527,3534
to|3535,3537
the|3538,3541
floor|3542,3547
,|3547,3548
the|3549,3552
patient|3553,3560
reports|3561,3568
the|3569,3572
pain|3573,3577
is|3578,3580
_|3581,3582
_|3582,3583
_|3583,3584
.|3584,3585
<EOL>|3585,3586
She|3586,3589
reports|3590,3597
again|3598,3603
that|3604,3608
this|3609,3613
pain|3614,3618
is|3619,3621
similar|3622,3629
to|3630,3632
the|3633,3636
pain|3637,3641
she|3642,3645
had|3646,3649
<EOL>|3649,3650
on|3650,3652
_|3653,3654
_|3654,3655
_|3655,3656
but|3657,3660
even|3661,3665
then|3666,3670
an|3671,3673
ultrasound|3674,3684
showed|3685,3691
no|3692,3694
DVT|3695,3698
.|3698,3699
She|3700,3703
is|3704,3706
able|3707,3711
<EOL>|3712,3713
to|3713,3715
<EOL>|3715,3716
move|3716,3720
her|3721,3724
toes|3725,3729
but|3730,3733
has|3734,3737
pain|3738,3742
with|3743,3747
lifting|3748,3755
her|3756,3759
leg|3760,3763
.|3763,3764
She|3765,3768
has|3769,3772
never|3773,3778
<EOL>|3778,3779
had|3779,3782
this|3783,3787
kind|3788,3792
of|3793,3795
pain|3796,3800
before|3801,3807
,|3807,3808
even|3809,3813
with|3814,3818
the|3819,3822
vein|3823,3827
stripping|3828,3837
that|3838,3842
<EOL>|3842,3843
she|3843,3846
had|3847,3850
in|3851,3853
the|3854,3857
past|3858,3862
(|3863,3864
age|3864,3867
_|3868,3869
_|3869,3870
_|3870,3871
.|3871,3872
She|3873,3876
has|3877,3880
no|3881,3883
chest|3884,3889
pain|3890,3894
or|3895,3897
shortness|3898,3907
<EOL>|3907,3908
of|3908,3910
breath|3911,3917
.|3917,3918
She|3919,3922
has|3923,3926
had|3927,3930
no|3931,3933
recent|3934,3940
travel|3941,3947
or|3948,3950
trauma|3951,3957
to|3958,3960
her|3961,3964
leg|3965,3968
.|3968,3969
<EOL>|3970,3971
<EOL>|3971,3972
<EOL>|3973,3974
Past|3974,3978
Medical|3979,3986
History|3987,3994
:|3994,3995
<EOL>|3995,3996
Dyslipidemia|3996,4008
,|4008,4009
<EOL>|4010,4011
Varicose|4011,4019
veins|4020,4025
(|4026,4027
R|4027,4028
>|4028,4029
L|4029,4030
)|4030,4031
s|4032,4033
/|4033,4034
p|4034,4035
ligation|4036,4044
,|4044,4045
<EOL>|4046,4047
COPD|4047,4051
,|4051,4052
<EOL>|4053,4054
OSA|4054,4057
(|4058,4059
+|4059,4060
CPap|4060,4064
)|4064,4065
,|4065,4066
<EOL>|4067,4068
recent|4068,4074
URI|4075,4078
(|4079,4080
received|4080,4088
course|4089,4095
of|4096,4098
Zithromax|4099,4108
)|4108,4109
,|4109,4110
<EOL>|4111,4112
bilateral|4112,4121
PEs|4122,4125
(|4126,4127
_|4127,4128
_|4128,4129
_|4129,4130
)|4130,4131
,|4131,4132
<EOL>|4133,4134
antiphospholipid|4134,4150
antibody|4151,4159
syndrome|4160,4168
(|4169,4170
on|4170,4172
lifelong|4173,4181
<EOL>|4182,4183
anticoagulation|4183,4198
)|4198,4199
,|4199,4200
<EOL>|4200,4201
<EOL>|4201,4202
T2DM|4202,4206
(|4207,4208
last|4208,4212
A1C|4213,4216
6.2|4217,4220
on|4221,4223
_|4224,4225
_|4225,4226
_|4226,4227
,|4227,4228
<EOL>|4229,4230
cerebral|4230,4238
aneurysm|4239,4247
(|4248,4249
followed|4249,4257
by|4258,4260
Dr.|4261,4264
_|4265,4266
_|4266,4267
_|4267,4268
,|4268,4269
unchanged|4270,4279
)|4279,4280
,|4280,4281
<EOL>|4282,4283
GERD|4283,4287
,|4287,4288
<EOL>|4289,4290
diverticulosis|4290,4304
,|4304,4305
<EOL>|4306,4307
h|4307,4308
/|4308,4309
o|4309,4310
colon|4311,4316
polyps|4317,4323
,|4323,4324
<EOL>|4325,4326
depression|4326,4336
,|4336,4337
<EOL>|4338,4339
s|4339,4340
/|4340,4341
p|4341,4342
right|4343,4348
CMC|4349,4352
joint|4353,4358
arthroplasty|4359,4371
,|4371,4372
<EOL>|4373,4374
b|4374,4375
/|4375,4376
l|4376,4377
rotator|4378,4385
cuff|4386,4390
repair|4391,4397
,|4397,4398
<EOL>|4399,4400
excision|4400,4408
right|4409,4414
_|4415,4416
_|4416,4417
_|4417,4418
digit|4419,4424
mass|4425,4429
,|4429,4430
<EOL>|4431,4432
CCY|4432,4435
w|4436,4437
/|4437,4438
stone|4438,4443
&|4444,4445
pancreatic|4446,4456
duct|4457,4461
exploration|4462,4473
(|4474,4475
_|4475,4476
_|4476,4477
_|4477,4478
)|4478,4479
,|4479,4480
<EOL>|4481,4482
hysterectomy|4482,4494
,|4494,4495
<EOL>|4496,4497
tonsillectomy|4497,4510
<EOL>|4511,4512
<EOL>|4512,4513
<EOL>|4514,4515
Social|4515,4521
History|4522,4529
:|4529,4530
<EOL>|4530,4531
_|4531,4532
_|4532,4533
_|4533,4534
<EOL>|4534,4535
Family|4535,4541
History|4542,4549
:|4549,4550
<EOL>|4550,4551
Mother|4551,4557
_|4558,4559
_|4559,4560
_|4560,4561
_|4562,4563
_|4563,4564
_|4564,4565
OVARIAN|4566,4573
CANCER|4574,4580
dx|4581,4583
age|4584,4587
_|4588,4589
_|4589,4590
_|4590,4591
<EOL>|4592,4593
Father|4593,4599
_|4600,4601
_|4601,4602
_|4602,4603
_|4604,4605
_|4605,4606
_|4606,4607
BRAIN|4608,4613
CANCER|4614,4620
<EOL>|4621,4622
PGM|4622,4625
OVARIAN|4626,4633
CANCER|4634,4640
<EOL>|4641,4642
Aunt|4642,4646
OVARIAN|4647,4654
CANCER|4655,4661
paternal|4662,4670
aunt|4671,4675
in|4676,4678
<EOL>|4679,4680
_|4681,4682
_|4682,4683
_|4683,4684
<EOL>|4685,4686
MGM|4686,4689
ENDOMETRIAL|4690,4701
CANCER|4702,4708
<EOL>|4709,4710
MGF|4710,4713
PROSTATE|4714,4722
CANCER|4723,4729
<EOL>|4730,4731
Brother|4731,4738
_|4739,4740
_|4740,4741
_|4741,4742
_|4743,4744
_|4744,4745
_|4745,4746
KIDNEY|4747,4753
CANCER|4754,4760
<EOL>|4761,4762
RENAL|4763,4768
FAILURE|4769,4776
<EOL>|4777,4778
CONGESTIVE|4779,4789
HEART|4790,4795
<EOL>|4796,4797
FAILURE|4798,4805
<EOL>|4806,4807
DIABETES|4808,4816
MELLITUS|4817,4825
<EOL>|4826,4827
TOBACCO|4828,4835
ABUSE|4836,4841
<EOL>|4842,4843
ALCOHOL|4844,4851
ABUSE|4852,4857
<EOL>|4858,4859
Sister|4859,4865
_|4866,4867
_|4867,4868
_|4868,4869
_|4870,4871
_|4871,4872
_|4872,4873
OVARIAN|4874,4881
CANCER|4882,4888
dx|4889,4891
age|4892,4895
_|4896,4897
_|4897,4898
_|4898,4899
<EOL>|4900,4901
Brother|4901,4908
_|4909,4910
_|4910,4911
_|4911,4912
THROAT|4913,4919
CANCER|4920,4926
dx|4927,4929
age|4930,4933
_|4934,4935
_|4935,4936
_|4936,4937
,|4937,4938
died|4939,4943
in|4944,4946
<EOL>|4947,4948
_|4949,4950
_|4950,4951
_|4951,4952
<EOL>|4953,4954
Sister|4954,4960
BRCA1|4961,4966
MUTATION|4967,4975
,|4975,4976
BREAST|4977,4983
CANCER|4984,4990
<EOL>|4991,4992
Daughter|4992,5000
Living|5001,5007
_|5008,5009
_|5009,5010
_|5010,5011
ABNORMAL|5012,5020
PAP|5021,5024
SMEAR|5025,5030
_|5031,5032
_|5032,5033
_|5033,5034
<EOL>|5034,5035
SUBSTANCE|5036,5045
ABUSE|5046,5051
<EOL>|5052,5053
Son|5053,5056
Died|5057,5061
_|5062,5063
_|5063,5064
_|5064,5065
SUBSTANCE|5066,5075
ABUSE|5076,5081
_|5082,5083
_|5083,5084
_|5084,5085
-|5086,5087
heroin|5088,5094
overdose|5095,5103
on|5104,5106
_|5107,5108
_|5108,5109
_|5109,5110
.|5110,5111
<EOL>|5111,5112
<EOL>|5113,5114
Physical|5114,5122
Exam|5123,5127
:|5127,5128
<EOL>|5128,5129
ADMISSION|5129,5138
EXAM|5139,5143
:|5143,5144
<EOL>|5144,5145
=|5145,5146
=|5146,5147
=|5147,5148
=|5148,5149
=|5149,5150
=|5150,5151
=|5151,5152
=|5152,5153
=|5153,5154
=|5154,5155
=|5155,5156
=|5156,5157
=|5157,5158
=|5158,5159
=|5159,5160
=|5160,5161
=|5161,5162
=|5162,5163
<EOL>|5163,5164
VITALS|5164,5170
:|5170,5171
T|5173,5174
97.9|5175,5179
BP|5180,5182
125|5183,5186
/|5187,5188
80|5189,5191
HR|5192,5194
82|5195,5197
RR|5198,5200
16|5201,5203
O2|5205,5207
Sat|5208,5211
94|5212,5214
RA|5215,5217
<EOL>|5218,5219
General|5219,5226
:|5226,5227
Alert|5228,5233
,|5233,5234
oriented|5235,5243
,|5243,5244
no|5245,5247
acute|5248,5253
distress|5254,5262
<EOL>|5264,5265
HEENT|5265,5270
:|5270,5271
MMM|5272,5275
,|5275,5276
oropharynx|5277,5287
clear|5288,5293
,|5293,5294
EOMI|5295,5299
,|5299,5300
PERRL|5301,5306
,|5306,5307
neck|5308,5312
supple|5313,5319
,|5319,5320
JVP|5321,5324
not|5325,5328
<EOL>|5328,5329
elevated|5329,5337
<EOL>|5337,5338
Chest|5338,5343
:|5343,5344
L|5345,5346
breast|5347,5353
incisions|5354,5363
well|5364,5368
healed|5369,5375
.|5375,5376
S|5377,5378
/|5378,5379
p|5379,5380
L|5381,5382
axilla|5383,5389
surgical|5390,5398
<EOL>|5398,5399
drain|5399,5404
removal|5405,5412
.|5412,5413
<EOL>|5413,5414
CV|5414,5416
:|5416,5417
Regular|5418,5425
rate|5426,5430
and|5431,5434
rhythm|5435,5441
,|5441,5442
normal|5443,5449
S1|5450,5452
+|5453,5454
S2|5455,5457
,|5457,5458
no|5459,5461
murmurs|5462,5469
<EOL>|5469,5470
Lungs|5470,5475
:|5475,5476
Clear|5477,5482
to|5483,5485
auscultation|5486,5498
bilaterally|5499,5510
,|5510,5511
no|5512,5514
wheezes|5515,5522
or|5523,5525
crackles|5526,5534
<EOL>|5534,5535
Abdomen|5535,5542
:|5542,5543
Soft|5544,5548
,|5548,5549
non-tender|5550,5560
,|5560,5561
non-distended|5562,5575
,|5575,5576
bowel|5577,5582
sounds|5583,5589
present|5590,5597
<EOL>|5597,5598
Ext|5598,5601
:|5601,5602
Warm|5603,5607
,|5607,5608
well|5609,5613
perfused|5614,5622
,|5622,5623
right|5624,5629
lower|5630,5635
extremity|5636,5645
is|5646,5648
tender|5649,5655
to|5656,5658
<EOL>|5658,5659
palpation|5659,5668
and|5669,5672
movement|5673,5681
limited|5682,5689
by|5690,5692
pain|5693,5697
.|5697,5698
Swelling|5699,5707
of|5708,5710
RLE|5711,5714
>|5715,5716
LLE|5717,5720
.|5720,5721
<EOL>|5721,5722
Palpable|5722,5730
2|5731,5732
+|5732,5733
_|5734,5735
_|5735,5736
_|5736,5737
pulses|5738,5744
bilaterally|5745,5756
.|5756,5757
<EOL>|5757,5758
Skin|5758,5762
:|5762,5763
Warm|5764,5768
,|5768,5769
dry|5770,5773
,|5773,5774
varicose|5775,5783
veins|5784,5789
noted|5790,5795
in|5796,5798
lower|5799,5804
extremities|5805,5816
.|5816,5817
<EOL>|5818,5819
Neuro|5819,5824
:|5824,5825
CNII|5826,5830
-|5830,5831
XII|5831,5834
intact|5835,5841
,|5841,5842
grossly|5843,5850
normal|5851,5857
strength|5858,5866
and|5867,5870
sensation|5871,5880
<EOL>|5881,5882
and|5882,5885
<EOL>|5885,5886
symmetric|5886,5895
bilaterally|5896,5907
<EOL>|5907,5908
<EOL>|5908,5909
DISCHARGE|5909,5918
EXAM|5919,5923
:|5923,5924
<EOL>|5924,5925
=|5925,5926
=|5926,5927
=|5927,5928
=|5928,5929
=|5929,5930
=|5930,5931
=|5931,5932
=|5932,5933
=|5933,5934
=|5934,5935
=|5935,5936
=|5936,5937
=|5937,5938
=|5938,5939
=|5939,5940
=|5940,5941
<EOL>|5941,5942
VITALS|5942,5948
:|5948,5949
Temp|5950,5954
:|5954,5955
98.2|5956,5960
(|5961,5962
Tm|5962,5964
98.9|5965,5969
)|5969,5970
,|5970,5971
BP|5972,5974
:|5974,5975
133|5976,5979
/|5979,5980
74|5980,5982
(|5983,5984
127|5984,5987
-|5987,5988
147|5988,5991
/|5991,5992
72|5992,5994
-|5994,5995
83|5995,5997
)|5997,5998
,|5998,5999
HR|6000,6002
:|6002,6003
76|6004,6006
<EOL>|6006,6007
(|6007,6008
76|6008,6010
-|6010,6011
91|6011,6013
)|6013,6014
,|6014,6015
RR|6016,6018
:|6018,6019
18|6020,6022
,|6022,6023
O2|6024,6026
sat|6027,6030
:|6030,6031
99|6032,6034
%|6034,6035
(|6036,6037
90|6037,6039
-|6039,6040
99|6040,6042
)|6042,6043
,|6043,6044
O2|6045,6047
delivery|6048,6056
:|6056,6057
Ra|6058,6060
<EOL>|6065,6066
General|6066,6073
:|6073,6074
Alert|6075,6080
,|6080,6081
oriented|6082,6090
,|6090,6091
no|6092,6094
acute|6095,6100
distress|6101,6109
<EOL>|6111,6112
HEENT|6112,6117
:|6117,6118
MMM|6119,6122
,|6122,6123
oropharynx|6124,6134
clear|6135,6140
,|6140,6141
EOMI|6142,6146
,|6146,6147
PERRL|6148,6153
,|6153,6154
neck|6155,6159
supple|6160,6166
,|6166,6167
JVP|6168,6171
not|6172,6175
<EOL>|6175,6176
elevated|6176,6184
<EOL>|6184,6185
Chest|6185,6190
:|6190,6191
L|6192,6193
breast|6194,6200
incisions|6201,6210
well|6211,6215
healed|6216,6222
.|6222,6223
S|6224,6225
/|6225,6226
p|6226,6227
L|6228,6229
axilla|6230,6236
surgical|6237,6245
<EOL>|6245,6246
drain|6246,6251
removal|6252,6259
.|6259,6260
<EOL>|6260,6261
CV|6261,6263
:|6263,6264
RRR|6265,6268
,|6268,6269
no|6270,6272
murmurs|6273,6280
<EOL>|6280,6281
Lungs|6281,6286
:|6286,6287
Clear|6288,6293
<EOL>|6293,6294
Abdomen|6294,6301
:|6301,6302
Soft|6303,6307
,|6307,6308
non-tender|6309,6319
,|6319,6320
non-distended|6321,6334
,|6334,6335
bowel|6336,6341
sounds|6342,6348
present|6349,6356
<EOL>|6356,6357
Ext|6357,6360
:|6360,6361
Warm|6362,6366
,|6366,6367
well|6368,6372
perfused|6373,6381
.|6381,6382
No|6383,6385
asymmetric|6386,6396
swelling|6397,6405
.|6405,6406
Minimally|6407,6416
<EOL>|6416,6417
tender|6417,6423
to|6424,6426
palpation|6427,6436
along|6437,6442
the|6443,6446
right|6447,6452
trochanteric|6453,6465
bursa|6466,6471
and|6472,6475
<EOL>|6475,6476
minimally|6476,6485
tender|6486,6492
to|6493,6495
palpation|6496,6505
along|6506,6511
the|6512,6515
right|6516,6521
tibia|6522,6527
.|6527,6528
Normal|6529,6535
ROM|6536,6539
<EOL>|6539,6540
though|6540,6546
pain|6547,6551
elicited|6552,6560
with|6561,6565
knee|6566,6570
flexion|6571,6578
;|6578,6579
improves|6580,6588
with|6589,6593
leg|6594,6597
raise|6598,6603
<EOL>|6603,6604
and|6604,6607
extension|6608,6617
.|6617,6618
Palpable|6619,6627
2|6628,6629
+|6629,6630
_|6631,6632
_|6632,6633
_|6633,6634
pulses|6635,6641
bilaterally|6642,6653
.|6653,6654
<EOL>|6654,6655
Skin|6655,6659
:|6659,6660
varicose|6661,6669
veins|6670,6675
noted|6676,6681
in|6682,6684
lower|6685,6690
extremities|6691,6702
.|6702,6703
<EOL>|6704,6705
Neuro|6705,6710
:|6710,6711
lower|6712,6717
extremity|6718,6727
sensation|6728,6737
is|6738,6740
equal|6741,6746
on|6747,6749
both|6750,6754
sides|6755,6760
to|6761,6763
light|6764,6769
<EOL>|6769,6770
touch|6770,6775
.|6775,6776
Normal|6777,6783
bilateral|6784,6793
lower|6794,6799
extremity|6800,6809
strength|6810,6818
.|6818,6819
Negative|6820,6828
<EOL>|6828,6829
babinsky|6829,6837
.|6837,6838
Ambulating|6840,6850
in|6851,6853
hallway|6854,6861
independently|6862,6875
though|6876,6882
it|6883,6885
<EOL>|6886,6887
precipitates|6887,6899
<EOL>|6900,6901
right|6901,6906
tibial|6907,6913
pain|6914,6918
<EOL>|6918,6919
<EOL>|6920,6921
Pertinent|6921,6930
Results|6931,6938
:|6938,6939
<EOL>|6939,6940
ADMISSION|6940,6949
LABS|6950,6954
:|6954,6955
<EOL>|6955,6956
=|6956,6957
=|6957,6958
=|6958,6959
=|6959,6960
=|6960,6961
=|6961,6962
=|6962,6963
=|6963,6964
=|6964,6965
=|6965,6966
=|6966,6967
=|6967,6968
=|6968,6969
=|6969,6970
=|6970,6971
=|6971,6972
<EOL>|6972,6973
_|6973,6974
_|6974,6975
_|6975,6976
12|6977,6979
:|6979,6980
00PM|6980,6984
BLOOD|6985,6990
WBC|6991,6994
-|6994,6995
5.6|6995,6998
RBC|6999,7002
-|7002,7003
3|7003,7004
.|7004,7005
48|7005,7007
*|7007,7008
Hgb|7009,7012
-|7012,7013
10|7013,7015
.|7015,7016
8|7016,7017
*|7017,7018
Hct|7019,7022
-|7022,7023
32|7023,7025
.|7025,7026
3|7026,7027
*|7027,7028
<EOL>|7029,7030
MCV|7030,7033
-|7033,7034
93|7034,7036
MCH|7037,7040
-|7040,7041
31.0|7041,7045
MCHC|7046,7050
-|7050,7051
33.4|7051,7055
RDW|7056,7059
-|7059,7060
14.7|7060,7064
RDWSD|7065,7070
-|7070,7071
48|7071,7073
.|7073,7074
6|7074,7075
*|7075,7076
Plt|7077,7080
_|7081,7082
_|7082,7083
_|7083,7084
<EOL>|7084,7085
_|7085,7086
_|7086,7087
_|7087,7088
12|7089,7091
:|7091,7092
00PM|7092,7096
BLOOD|7097,7102
Neuts|7103,7108
-|7108,7109
73|7109,7111
.|7111,7112
6|7112,7113
*|7113,7114
_|7115,7116
_|7116,7117
_|7117,7118
Monos|7119,7124
-|7124,7125
4|7125,7126
.|7126,7127
9|7127,7128
*|7128,7129
<EOL>|7130,7131
Eos|7131,7134
-|7134,7135
0|7135,7136
.|7136,7137
9|7137,7138
*|7138,7139
Baso|7140,7144
-|7144,7145
0.7|7145,7148
Im|7149,7151
_|7152,7153
_|7153,7154
_|7154,7155
AbsNeut|7156,7163
-|7163,7164
4|7164,7165
.|7165,7166
09|7166,7168
AbsLymp|7169,7176
-|7176,7177
1|7177,7178
.|7178,7179
08|7179,7181
*|7181,7182
<EOL>|7183,7184
AbsMono|7184,7191
-|7191,7192
0|7192,7193
.|7193,7194
27|7194,7196
AbsEos|7197,7203
-|7203,7204
0|7204,7205
.|7205,7206
05|7206,7208
AbsBaso|7209,7216
-|7216,7217
0.04|7217,7221
<EOL>|7221,7222
_|7222,7223
_|7223,7224
_|7224,7225
12|7226,7228
:|7228,7229
00PM|7229,7233
BLOOD|7234,7239
_|7240,7241
_|7241,7242
_|7242,7243
PTT|7244,7247
-|7247,7248
28.2|7248,7252
_|7253,7254
_|7254,7255
_|7255,7256
<EOL>|7256,7257
_|7257,7258
_|7258,7259
_|7259,7260
12|7261,7263
:|7263,7264
00PM|7264,7268
BLOOD|7269,7274
Glucose|7275,7282
-|7282,7283
107|7283,7286
*|7286,7287
UreaN|7288,7293
-|7293,7294
7|7294,7295
Creat|7296,7301
-|7301,7302
0.8|7302,7305
Na|7306,7308
-|7308,7309
139|7309,7312
<EOL>|7313,7314
K|7314,7315
-|7315,7316
4.0|7316,7319
Cl|7320,7322
-|7322,7323
100|7323,7326
HCO3|7327,7331
-|7331,7332
26|7332,7334
AnGap|7335,7340
-|7340,7341
13|7341,7343
<EOL>|7343,7344
_|7344,7345
_|7345,7346
_|7346,7347
05|7348,7350
:|7350,7351
40AM|7351,7355
BLOOD|7356,7361
Calcium|7362,7369
-|7369,7370
8.6|7370,7373
Phos|7374,7378
-|7378,7379
4|7379,7380
.|7380,7381
8|7381,7382
*|7382,7383
Mg|7384,7386
-|7386,7387
2.2|7387,7390
Iron|7391,7395
-|7395,7396
36|7396,7398
<EOL>|7398,7399
_|7399,7400
_|7400,7401
_|7401,7402
05|7403,7405
:|7405,7406
40AM|7406,7410
BLOOD|7411,7416
calTIBC|7417,7424
-|7424,7425
291|7425,7428
VitB12|7429,7435
-|7435,7436
331|7436,7439
Ferritn|7440,7447
-|7447,7448
50|7448,7450
TRF|7451,7454
-|7454,7455
224|7455,7458
<EOL>|7458,7459
_|7459,7460
_|7460,7461
_|7461,7462
07|7463,7465
:|7465,7466
15AM|7466,7470
BLOOD|7471,7476
25VitD|7477,7483
-|7483,7484
45|7484,7486
<EOL>|7486,7487
_|7487,7488
_|7488,7489
_|7489,7490
12|7491,7493
:|7493,7494
25PM|7494,7498
BLOOD|7499,7504
Lactate|7505,7512
-|7512,7513
1.1|7513,7516
<EOL>|7516,7517
<EOL>|7517,7518
DISCHARGE|7518,7527
LABS|7528,7532
:|7532,7533
<EOL>|7533,7534
=|7534,7535
=|7535,7536
=|7536,7537
=|7537,7538
=|7538,7539
=|7539,7540
=|7540,7541
=|7541,7542
=|7542,7543
=|7543,7544
=|7544,7545
=|7545,7546
=|7546,7547
=|7547,7548
=|7548,7549
=|7549,7550
<EOL>|7550,7551
_|7551,7552
_|7552,7553
_|7553,7554
04|7555,7557
:|7557,7558
41AM|7558,7562
BLOOD|7563,7568
WBC|7569,7572
-|7572,7573
5.6|7573,7576
RBC|7577,7580
-|7580,7581
3|7581,7582
.|7582,7583
36|7583,7585
*|7585,7586
Hgb|7587,7590
-|7590,7591
10|7591,7593
.|7593,7594
1|7594,7595
*|7595,7596
Hct|7597,7600
-|7600,7601
31|7601,7603
.|7603,7604
1|7604,7605
*|7605,7606
<EOL>|7607,7608
MCV|7608,7611
-|7611,7612
93|7612,7614
MCH|7615,7618
-|7618,7619
30.1|7619,7623
MCHC|7624,7628
-|7628,7629
32.5|7629,7633
RDW|7634,7637
-|7637,7638
14.5|7638,7642
RDWSD|7643,7648
-|7648,7649
48|7649,7651
.|7651,7652
7|7652,7653
*|7653,7654
Plt|7655,7658
_|7659,7660
_|7660,7661
_|7661,7662
<EOL>|7662,7663
_|7663,7664
_|7664,7665
_|7665,7666
04|7667,7669
:|7669,7670
41AM|7670,7674
BLOOD|7675,7680
_|7681,7682
_|7682,7683
_|7683,7684
<EOL>|7684,7685
_|7685,7686
_|7686,7687
_|7687,7688
04|7689,7691
:|7691,7692
41AM|7692,7696
BLOOD|7697,7702
Glucose|7703,7710
-|7710,7711
132|7711,7714
*|7714,7715
UreaN|7716,7721
-|7721,7722
15|7722,7724
Creat|7725,7730
-|7730,7731
0.7|7731,7734
Na|7735,7737
-|7737,7738
140|7738,7741
<EOL>|7742,7743
K|7743,7744
-|7744,7745
5.0|7745,7748
Cl|7749,7751
-|7751,7752
103|7752,7755
HCO3|7756,7760
-|7760,7761
26|7761,7763
AnGap|7764,7769
-|7769,7770
11|7770,7772
<EOL>|7772,7773
_|7773,7774
_|7774,7775
_|7775,7776
04|7777,7779
:|7779,7780
41AM|7780,7784
BLOOD|7785,7790
Calcium|7791,7798
-|7798,7799
9.2|7799,7802
Phos|7803,7807
-|7807,7808
4.0|7808,7811
Mg|7812,7814
-|7814,7815
2.4|7815,7818
<EOL>|7818,7819
<EOL>|7819,7820
IMAGING|7820,7827
:|7827,7828
<EOL>|7828,7829
=|7829,7830
=|7830,7831
=|7831,7832
=|7832,7833
=|7833,7834
=|7834,7835
=|7835,7836
=|7836,7837
=|7837,7838
=|7838,7839
=|7839,7840
=|7840,7841
=|7841,7842
=|7842,7843
=|7843,7844
=|7844,7845
=|7845,7846
=|7846,7847
=|7847,7848
<EOL>|7848,7849
Unilat|7849,7855
lower|7856,7861
extremity|7862,7871
vein|7872,7876
-|7876,7877
R|7878,7879
_|7880,7881
_|7881,7882
_|7882,7883
<EOL>|7883,7884
Right|7884,7889
calf|7890,7894
veins|7895,7900
not|7901,7904
visualized|7905,7915
.|7915,7916
Otherwise|7917,7926
,|7926,7927
no|7928,7930
evidence|7931,7939
of|7940,7942
deep|7943,7947
<EOL>|7947,7948
venous|7948,7954
thrombosis|7955,7965
in|7966,7968
the|7969,7972
right|7973,7978
lower|7979,7984
extremity|7985,7994
veins|7995,8000
.|8000,8001
<EOL>|8001,8002
<EOL>|8002,8003
CT|8003,8005
RLE|8006,8009
_|8010,8011
_|8011,8012
_|8012,8013
<EOL>|8013,8014
Unremarkable|8014,8026
contrast|8027,8035
enhanced|8036,8044
CT|8045,8047
of|8048,8050
the|8051,8054
right|8055,8060
calf|8061,8065
with|8066,8070
a|8071,8072
two|8073,8076
<EOL>|8077,8078
vessel|8078,8084
runoff|8085,8091
to|8092,8094
the|8095,8098
foot|8099,8103
.|8103,8104
<EOL>|8105,8106
The|8106,8109
veins|8110,8115
of|8116,8118
the|8119,8122
lower|8123,8128
extremity|8129,8138
are|8139,8142
not|8143,8146
opacified|8147,8156
therefore|8157,8166
<EOL>|8167,8168
can|8168,8171
not|8171,8174
be|8175,8177
assessed|8178,8186
for|8187,8190
patency|8191,8198
.|8198,8199
Consider|8201,8209
repeat|8210,8216
ultrasound|8217,8227
to|8228,8230
<EOL>|8231,8232
more|8232,8236
fully|8237,8242
evaluate|8243,8251
.|8251,8252
<EOL>|8253,8254
No|8254,8256
focal|8257,8262
collection|8263,8273
or|8274,8276
obvious|8277,8284
muscular|8285,8293
abnormality|8294,8305
identified|8306,8316
<EOL>|8317,8318
by|8318,8320
CT|8321,8323
<EOL>|8323,8324
<EOL>|8324,8325
_|8325,8326
_|8326,8327
_|8327,8328
:|8328,8329
<EOL>|8329,8330
1.|8330,8332
.|8332,8333
Uneventful|8335,8345
ultrasound|8346,8356
-|8356,8357
guided|8357,8363
injection|8364,8373
of|8374,8376
long|8377,8381
-|8381,8382
acting|8382,8388
<EOL>|8389,8390
anesthetic|8390,8400
and|8401,8404
<EOL>|8404,8405
steroid|8405,8412
into|8413,8417
theright|8418,8426
greater|8427,8434
trochanteric|8435,8447
bursa|8448,8453
.|8453,8454
<EOL>|8454,8455
2.|8455,8457
Prior|8459,8464
injection|8465,8474
,|8474,8475
small|8476,8481
amount|8482,8488
of|8489,8491
fluid|8492,8497
in|8498,8500
the|8501,8504
right|8505,8510
greater|8511,8518
<EOL>|8519,8520
trochanteric|8520,8532
<EOL>|8532,8533
bursa|8533,8538
and|8539,8542
dystrophic|8543,8553
calcification|8554,8567
within|8568,8574
the|8575,8578
bursal|8579,8585
space|8586,8591
.|8591,8592
<EOL>|8594,8595
Findings|8595,8603
raise|8604,8609
<EOL>|8609,8610
suspicion|8610,8619
for|8620,8623
chronic|8624,8631
trochanteric|8632,8644
bursitis|8645,8653
.|8653,8654
<EOL>|8654,8655
<EOL>|8656,8657
Brief|8657,8662
Hospital|8663,8671
Course|8672,8678
:|8678,8679
<EOL>|8679,8680
SUMMARY|8680,8687
:|8687,8688
<EOL>|8688,8689
=|8689,8690
=|8690,8691
=|8691,8692
=|8692,8693
=|8693,8694
=|8694,8695
=|8695,8696
=|8696,8697
=|8697,8698
=|8698,8699
=|8699,8700
=|8700,8701
=|8701,8702
=|8702,8703
=|8703,8704
=|8704,8705
=|8705,8706
=|8706,8707
<EOL>|8707,8708
Ms.|8708,8711
_|8712,8713
_|8713,8714
_|8714,8715
is|8716,8718
a|8719,8720
_|8721,8722
_|8722,8723
_|8723,8724
with|8725,8729
a|8730,8731
PMH|8732,8735
significant|8736,8747
for|8748,8751
<EOL>|8752,8753
antiphospholipid|8753,8769
syndrome|8770,8778
with|8779,8783
DVTs|8784,8788
and|8789,8792
PEs|8793,8796
on|8797,8799
Coumadin|8800,8808
,|8808,8809
recent|8810,8816
<EOL>|8817,8818
L|8818,8819
-|8819,8820
sided|8820,8825
breast|8826,8832
cancer|8833,8839
s|8840,8841
/|8841,8842
p|8842,8843
lumpectomy|8844,8854
,|8854,8855
who|8856,8859
presented|8860,8869
to|8870,8872
the|8873,8876
ED|8877,8879
<EOL>|8880,8881
with|8881,8885
acute|8886,8891
on|8892,8894
chronic|8895,8902
right|8903,8908
lower|8909,8914
extremity|8915,8924
and|8925,8928
right|8929,8934
hip|8935,8938
pain|8939,8943
,|8943,8944
<EOL>|8945,8946
making|8946,8952
it|8953,8955
difficult|8956,8965
to|8966,8968
ambulate|8969,8977
.|8977,8978
Right|8979,8984
lower|8985,8990
extremity|8991,9000
U|9001,9002
/|9002,9003
S|9003,9004
and|9005,9008
<EOL>|9009,9010
CT|9010,9012
did|9013,9016
not|9017,9020
reveal|9021,9027
a|9028,9029
DVT|9030,9033
though|9034,9040
calf|9041,9045
veins|9046,9051
were|9052,9056
not|9057,9060
well|9061,9065
<EOL>|9066,9067
visualized|9067,9077
.|9077,9078
<EOL>|9079,9080
<EOL>|9080,9081
ACTIVE|9081,9087
ISSUES|9088,9094
:|9094,9095
<EOL>|9095,9096
=|9096,9097
=|9097,9098
=|9098,9099
=|9099,9100
=|9100,9101
=|9101,9102
=|9102,9103
=|9103,9104
=|9104,9105
=|9105,9106
=|9106,9107
=|9107,9108
=|9108,9109
=|9109,9110
=|9110,9111
=|9111,9112
=|9112,9113
=|9113,9114
<EOL>|9114,9115
#|9115,9116
Right|9117,9122
trochanteric|9123,9135
bursitis|9136,9144
<EOL>|9144,9145
#|9145,9146
Right|9147,9152
anterior|9153,9161
lower|9162,9167
leg|9168,9171
pain|9172,9176
<EOL>|9176,9177
#|9177,9178
Right|9179,9184
sided|9185,9190
varicose|9191,9199
veins|9200,9205
<EOL>|9205,9206
Pt|9206,9208
endorsed|9209,9217
>|9218,9219
4mths|9219,9224
of|9225,9227
pain|9228,9232
in|9233,9235
RLE|9236,9239
that|9240,9244
became|9245,9251
acutely|9252,9259
worse|9260,9265
over|9266,9270
<EOL>|9271,9272
the|9272,9275
last|9276,9280
few|9281,9284
wks|9285,9288
.|9288,9289
Her|9291,9294
initial|9295,9302
exam|9303,9307
was|9308,9311
most|9312,9316
consistent|9317,9327
with|9328,9332
<EOL>|9333,9334
severe|9334,9340
trochanteric|9341,9353
bursitis|9354,9362
on|9363,9365
the|9366,9369
right|9370,9375
.|9375,9376
She|9377,9380
also|9381,9385
has|9386,9389
some|9390,9394
<EOL>|9395,9396
focal|9396,9401
pain|9402,9406
along|9407,9412
the|9413,9416
right|9417,9422
tibia|9423,9428
which|9429,9434
she|9435,9438
felt|9439,9443
was|9444,9447
most|9448,9452
<EOL>|9453,9454
consistent|9454,9464
with|9465,9469
pain|9470,9474
from|9475,9479
her|9480,9483
varicose|9484,9492
veins|9493,9498
.|9498,9499
The|9500,9503
XRs|9504,9507
of|9508,9510
her|9511,9514
<EOL>|9515,9516
tibia|9516,9521
/|9521,9522
fibula|9522,9528
and|9529,9532
right|9533,9538
hip|9539,9542
were|9543,9547
without|9548,9555
obvious|9556,9563
pathology|9564,9573
.|9573,9574
There|9575,9580
<EOL>|9581,9582
are|9582,9585
no|9586,9588
concerning|9589,9599
neurologic|9600,9610
symptoms|9611,9619
to|9620,9622
suggest|9623,9630
a|9631,9632
<EOL>|9633,9634
radiculopathy|9634,9647
,|9647,9648
no|9649,9651
weakness|9652,9660
or|9661,9663
numbness|9664,9672
though|9673,9679
she|9680,9683
may|9684,9687
have|9688,9692
some|9693,9697
<EOL>|9698,9699
degree|9699,9705
of|9706,9708
chronic|9709,9716
sciatica|9717,9725
.|9725,9726
Mildly|9728,9734
decreased|9735,9744
patellar|9745,9753
reflex|9754,9760
on|9761,9763
<EOL>|9764,9765
the|9765,9768
right|9769,9774
as|9775,9777
compared|9778,9786
to|9787,9789
left|9790,9794
may|9795,9798
have|9799,9803
been|9804,9808
in|9809,9811
the|9812,9815
setting|9816,9823
of|9824,9826
<EOL>|9827,9828
pain|9828,9832
and|9833,9836
guarding|9837,9845
;|9845,9846
strength|9847,9855
was|9856,9859
normal|9860,9866
bilaterally|9867,9878
as|9879,9881
was|9882,9885
her|9886,9889
<EOL>|9890,9891
sensation|9891,9900
.|9900,9901
<EOL>|9902,9903
She|9903,9906
underwent|9907,9916
U|9917,9918
/|9918,9919
S|9919,9920
guided|9921,9927
steroid|9928,9935
injection|9936,9945
of|9946,9948
her|9949,9952
trochanteric|9953,9965
<EOL>|9966,9967
bursa|9967,9972
w|9973,9974
/|9974,9975
significant|9976,9987
improvement|9988,9999
in|10000,10002
symptoms|10003,10011
;|10011,10012
_|10013,10014
_|10014,10015
_|10015,10016
stated|10017,10023
that|10024,10028
<EOL>|10029,10030
there|10030,10035
was|10036,10039
some|10040,10044
fluid|10045,10050
near|10051,10055
the|10056,10059
bursa|10060,10065
,|10065,10066
suggestive|10067,10077
of|10078,10080
acute|10081,10086
on|10087,10089
<EOL>|10090,10091
chronic|10091,10098
trochanteric|10099,10111
bursitis|10112,10120
.|10120,10121
Her|10122,10125
anterior|10126,10134
shin|10135,10139
pain|10140,10144
improved|10145,10153
<EOL>|10154,10155
with|10155,10159
initiation|10160,10170
of|10171,10173
gabapentin|10174,10184
and|10185,10188
lidocaine|10189,10198
patch|10199,10204
in|10205,10207
addition|10208,10216
to|10217,10219
<EOL>|10220,10221
her|10221,10224
home|10225,10229
tylenol|10230,10237
and|10238,10241
an|10242,10244
increase|10245,10253
in|10254,10256
the|10257,10260
frequency|10261,10270
of|10271,10273
her|10274,10277
home|10278,10282
<EOL>|10283,10284
tramadol|10284,10292
(|10293,10294
q8h|10294,10297
PRN|10298,10301
to|10302,10304
q4h|10305,10308
PRN|10309,10312
)|10312,10313
.|10313,10314
Pt|10316,10318
was|10319,10322
not|10323,10326
given|10327,10332
her|10333,10336
home|10337,10341
<EOL>|10342,10343
hydromorphone|10343,10356
PRN|10357,10360
,|10360,10361
though|10362,10368
she|10369,10372
did|10373,10376
require|10377,10384
one|10385,10388
dose|10389,10393
of|10394,10396
0.5|10397,10400
mg|10401,10403
IV|10404,10406
<EOL>|10407,10408
hydromorphone|10408,10421
following|10422,10431
her|10432,10435
injection|10436,10445
in|10446,10448
the|10449,10452
setting|10453,10460
of|10461,10463
an|10464,10466
acute|10467,10472
<EOL>|10473,10474
pain|10474,10478
episode|10479,10486
.|10486,10487
She|10488,10491
was|10492,10495
discharged|10496,10506
with|10507,10511
Tramadol|10512,10520
50mg|10521,10525
x15|10526,10529
tablets|10530,10537
<EOL>|10538,10539
given|10539,10544
increased|10545,10554
requirement|10555,10566
.|10566,10567
By|10568,10570
discharge|10571,10580
,|10580,10581
she|10582,10585
was|10586,10589
able|10590,10594
ambulate|10595,10603
<EOL>|10604,10605
and|10605,10608
was|10609,10612
felt|10613,10617
safe|10618,10622
for|10623,10626
discharge|10627,10636
home|10637,10641
with|10642,10646
a|10647,10648
cane|10649,10653
per|10654,10657
_|10658,10659
_|10659,10660
_|10660,10661
<EOL>|10662,10663
evaluation|10663,10673
.|10673,10674
Pt|10676,10678
was|10679,10682
eager|10683,10688
to|10689,10691
leave|10692,10697
and|10698,10701
will|10702,10706
reach|10707,10712
out|10713,10716
to|10717,10719
her|10720,10723
<EOL>|10724,10725
vascular|10725,10733
surgeon|10734,10741
for|10742,10745
an|10746,10748
appointment|10749,10760
early|10761,10766
in|10767,10769
the|10770,10773
new|10774,10777
year|10778,10782
for|10783,10786
<EOL>|10787,10788
treatment|10788,10797
of|10798,10800
her|10801,10804
painful|10805,10812
varicose|10813,10821
veins|10822,10827
.|10827,10828
<EOL>|10828,10829
<EOL>|10829,10830
#|10830,10831
Iron|10832,10836
deficiency|10837,10847
anemia|10848,10854
:|10854,10855
<EOL>|10855,10856
Anemia|10856,10862
is|10863,10865
new|10866,10869
since|10870,10875
_|10876,10877
_|10877,10878
_|10878,10879
.|10879,10880
Normocytic|10881,10891
.|10891,10892
Downtrended|10893,10904
overnight|10905,10914
to|10915,10917
<EOL>|10918,10919
8.9|10919,10922
from|10923,10927
10.8|10928,10932
.|10932,10933
No|10934,10936
concern|10937,10944
for|10945,10948
active|10949,10955
bleeding|10956,10964
.|10964,10965
Per|10966,10969
iron|10970,10974
studies|10975,10982
,|10982,10983
<EOL>|10984,10985
she|10985,10988
is|10989,10991
iron|10992,10996
deficient|10997,11006
with|11007,11011
a|11012,11013
ferritin|11014,11022
of|11023,11025
50|11026,11028
.|11028,11029
She|11030,11033
endorses|11034,11042
<EOL>|11043,11044
fatigue|11044,11051
and|11052,11055
restless|11056,11064
leg|11065,11068
syndrome|11069,11077
.|11077,11078
Etiology|11079,11087
is|11088,11090
unclear|11091,11098
,|11098,11099
though|11100,11106
<EOL>|11107,11108
it|11108,11110
may|11111,11114
be|11115,11117
related|11118,11125
to|11126,11128
the|11129,11132
recent|11133,11139
left|11140,11144
breast|11145,11151
hematoma|11152,11160
of|11161,11163
her|11164,11167
<EOL>|11168,11169
breast|11169,11175
(|11176,11177
unlikely|11177,11185
though|11186,11192
the|11193,11196
timing|11197,11203
fits|11204,11208
)|11208,11209
.|11209,11210
Prior|11211,11216
EGD|11217,11220
with|11221,11225
<EOL>|11226,11227
gastritis|11227,11236
(|11237,11238
_|11238,11239
_|11239,11240
_|11240,11241
)|11241,11242
for|11243,11246
which|11247,11252
she|11253,11256
is|11257,11259
on|11260,11262
a|11263,11264
BID|11265,11268
PPI|11269,11272
;|11272,11273
prior|11274,11279
<EOL>|11280,11281
colonoscopy|11281,11292
_|11293,11294
_|11294,11295
_|11295,11296
with|11297,11301
findings|11302,11310
that|11311,11315
may|11316,11319
be|11320,11322
suggestive|11323,11333
of|11334,11336
<EOL>|11337,11338
celiac|11338,11344
disease|11345,11352
,|11352,11353
though|11354,11360
ttg|11361,11364
at|11365,11367
that|11368,11372
time|11373,11377
was|11378,11381
normal|11382,11388
with|11389,11393
a|11394,11395
normal|11396,11402
<EOL>|11403,11404
IgA|11404,11407
.|11407,11408
She|11409,11412
also|11413,11417
had|11418,11421
two|11422,11425
polyps|11426,11432
biopsied|11433,11441
and|11442,11445
were|11446,11450
normal|11451,11457
.|11457,11458
On|11459,11461
this|11462,11466
<EOL>|11467,11468
admission|11468,11477
,|11477,11478
a|11479,11480
vitamin|11481,11488
D|11489,11490
level|11491,11496
was|11497,11500
obtained|11501,11509
to|11510,11512
assess|11513,11519
for|11520,11523
evidence|11524,11532
<EOL>|11533,11534
of|11534,11536
malabsorption|11537,11550
iso|11551,11554
daily|11555,11560
supplementation|11561,11576
:|11576,11577
level|11578,11583
was|11584,11587
45|11588,11590
.|11590,11591
She|11592,11595
<EOL>|11596,11597
was|11597,11600
given|11601,11606
ferric|11607,11613
gluconate|11614,11623
IV|11624,11626
x1|11627,11629
on|11630,11632
_|11633,11634
_|11634,11635
_|11635,11636
.|11636,11637
TTG|11638,11641
was|11642,11645
repeated|11646,11654
and|11655,11658
<EOL>|11659,11660
pending|11660,11667
at|11668,11670
discharge|11671,11680
.|11680,11681
<EOL>|11682,11683
<EOL>|11683,11684
CHRONIC|11684,11691
ISSUES|11692,11698
:|11698,11699
<EOL>|11699,11700
=|11700,11701
=|11701,11702
=|11702,11703
=|11703,11704
=|11704,11705
=|11705,11706
=|11706,11707
=|11707,11708
=|11708,11709
=|11709,11710
=|11710,11711
=|11711,11712
=|11712,11713
=|11713,11714
=|11714,11715
=|11715,11716
=|11716,11717
=|11717,11718
=|11718,11719
<EOL>|11719,11720
#|11720,11721
History|11722,11729
of|11730,11732
DVT|11733,11736
/|11736,11737
PE|11737,11739
on|11740,11742
warfarin|11743,11751
:|11751,11752
<EOL>|11752,11753
#|11753,11754
Antiphospholipid|11755,11771
antibody|11772,11780
syndrome|11781,11789
:|11789,11790
<EOL>|11790,11791
#|11791,11792
Subtherapeutic|11793,11807
INR|11808,11811
:|11811,11812
<EOL>|11812,11813
Lupus|11813,11818
anticoagulant|11819,11832
positive|11833,11841
in|11842,11844
_|11845,11846
_|11846,11847
_|11847,11848
.|11848,11849
She|11850,11853
has|11854,11857
been|11858,11862
taking|11863,11869
her|11870,11873
<EOL>|11874,11875
home|11875,11879
dose|11880,11884
of|11885,11887
warfarin|11888,11896
(|11897,11898
5|11898,11899
mg|11900,11902
_|11903,11904
_|11904,11905
_|11905,11906
and|11907,11910
7.5|11911,11914
mg|11915,11917
other|11918,11923
days|11924,11928
)|11928,11929
.|11929,11930
Her|11931,11934
<EOL>|11935,11936
warfarin|11936,11944
was|11945,11948
held|11949,11953
last|11954,11958
_|11959,11960
_|11960,11961
_|11961,11962
iso|11963,11966
hematoma|11967,11975
and|11976,11979
she|11980,11983
was|11984,11987
not|11988,11991
<EOL>|11992,11993
bridged|11993,12000
with|12001,12005
Lovenox|12006,12013
upon|12014,12018
reinitiation|12019,12031
.|12031,12032
INR|12033,12036
on|12037,12039
this|12040,12044
admission|12045,12054
<EOL>|12055,12056
was|12056,12059
subtherapeutic|12060,12074
at|12075,12077
1.4|12078,12081
.|12081,12082
Bridged|12083,12090
during|12091,12097
this|12098,12102
hospitalization|12103,12118
<EOL>|12119,12120
with|12120,12124
Lovenox|12125,12132
for|12133,12136
goal|12137,12141
INR|12142,12145
_|12146,12147
_|12147,12148
_|12148,12149
.|12149,12150
She|12151,12154
was|12155,12158
given|12159,12164
an|12165,12167
increased|12168,12177
dose|12178,12182
<EOL>|12183,12184
of|12184,12186
warfarin|12187,12195
,|12195,12196
7.5|12197,12200
mg|12201,12203
daily|12204,12209
while|12210,12215
in|12216,12218
house|12219,12224
.|12224,12225
INR|12226,12229
at|12230,12232
discharge|12233,12242
was|12243,12246
<EOL>|12247,12248
1.9|12248,12251
,|12251,12252
with|12253,12257
plan|12258,12262
to|12263,12265
continue|12266,12274
home|12275,12279
warfarin|12280,12288
regimen|12289,12296
.|12296,12297
Patient|12298,12305
will|12306,12310
<EOL>|12311,12312
get|12312,12315
repeat|12316,12322
INR|12323,12326
on|12327,12329
_|12330,12331
_|12331,12332
_|12332,12333
.|12333,12334
<EOL>|12335,12336
<EOL>|12336,12337
#|12337,12338
Vitamin|12339,12346
D|12347,12348
deficiency|12349,12359
:|12359,12360
pt|12361,12363
takes|12364,12369
2,000|12370,12375
U|12376,12377
vitamin|12378,12385
D|12386,12387
daily|12388,12393
.|12393,12394
Repeat|12395,12401
<EOL>|12402,12403
level|12403,12408
IS|12409,12411
45|12412,12414
which|12415,12420
suggests|12421,12429
against|12430,12437
malabsorption|12438,12451
to|12452,12454
account|12455,12462
for|12463,12466
<EOL>|12467,12468
her|12468,12471
iron|12472,12476
deficiency|12477,12487
.|12487,12488
<EOL>|12489,12490
<EOL>|12490,12491
TRANSITIONAL|12491,12503
ISSUES|12504,12510
:|12510,12511
<EOL>|12511,12512
=|12512,12513
=|12513,12514
=|12514,12515
=|12515,12516
=|12516,12517
=|12517,12518
=|12518,12519
=|12519,12520
=|12520,12521
=|12521,12522
=|12522,12523
=|12523,12524
=|12524,12525
=|12525,12526
=|12526,12527
=|12527,12528
=|12528,12529
=|12529,12530
=|12530,12531
=|12531,12532
<EOL>|12532,12533
Code|12533,12537
status|12538,12544
:|12544,12545
Full|12546,12550
,|12550,12551
presumed|12552,12560
<EOL>|12560,12561
HCP|12561,12564
:|12564,12565
_|12566,12567
_|12567,12568
_|12568,12569
,|12569,12570
granddaughter|12571,12584
-|12585,12586
_|12587,12588
_|12588,12589
_|12589,12590
.|12590,12591
<EOL>|12591,12592
<EOL>|12592,12593
-|12593,12594
Right|12595,12600
trochanteric|12601,12613
bursitis|12614,12622
:|12622,12623
<EOL>|12623,12624
[|12624,12625
]|12625,12626
Consider|12627,12635
repeat|12636,12642
injection|12643,12652
<EOL>|12652,12653
[|12653,12654
]|12654,12655
Consider|12656,12664
physical|12665,12673
therapy|12674,12681
<EOL>|12681,12682
<EOL>|12682,12683
-|12683,12684
Right|12685,12690
anterior|12691,12699
leg|12700,12703
pain|12704,12708
<EOL>|12708,12709
[|12709,12710
]|12710,12711
discharged|12712,12722
on|12723,12725
gabapentin|12726,12736
600|12737,12740
mg|12741,12743
three|12744,12749
times|12750,12755
daily|12756,12761
<EOL>|12761,12762
[|12762,12763
]|12763,12764
discharged|12765,12775
with|12776,12780
tramadol|12781,12789
50mg|12790,12794
,|12794,12795
home|12796,12800
regimen|12801,12808
is|12809,12811
Q8hrs|12812,12817
and|12818,12821
<EOL>|12822,12823
required|12823,12831
Q4hrs|12832,12837
during|12838,12844
hospitalization|12845,12860
.|12860,12861
Will|12862,12866
give|12867,12871
two|12872,12875
day|12876,12879
supply|12880,12886
<EOL>|12887,12888
of|12888,12890
increased|12891,12900
dose|12901,12905
.|12905,12906
Plan|12907,12911
to|12912,12914
see|12915,12918
PCP|12919,12922
next|12923,12927
week|12928,12932
.|12932,12933
<EOL>|12933,12934
[|12934,12935
]|12935,12936
Consider|12937,12945
outpatient|12946,12956
MRI|12957,12960
of|12961,12963
the|12964,12967
lumbar|12968,12974
spine|12975,12980
for|12981,12984
chronic|12985,12992
pain|12993,12997
<EOL>|12998,12999
[|12999,13000
]|13000,13001
Consider|13002,13010
EMG|13011,13014
<EOL>|13014,13015
[|13015,13016
]|13016,13017
Vascular|13018,13026
surgery|13027,13034
follow|13035,13041
up|13042,13044
as|13045,13047
outpt|13048,13053
for|13054,13057
treatment|13058,13067
of|13068,13070
painful|13071,13078
<EOL>|13079,13080
veins|13080,13085
<EOL>|13085,13086
<EOL>|13086,13087
-|13087,13088
Iron|13089,13093
deficiency|13094,13104
anemia|13105,13111
:|13111,13112
<EOL>|13112,13113
[|13113,13114
]|13114,13115
Consider|13116,13124
repeat|13125,13131
IV|13132,13134
iron|13135,13139
infusion|13140,13148
<EOL>|13148,13149
[|13149,13150
]|13150,13151
F|13152,13153
/|13153,13154
u|13154,13155
pending|13156,13163
TTG|13164,13167
<EOL>|13167,13168
[|13168,13169
]|13169,13170
Consider|13171,13179
further|13180,13187
work|13188,13192
up|13193,13195
(|13196,13197
though|13197,13203
may|13204,13207
be|13208,13210
related|13211,13218
to|13219,13221
left|13222,13226
<EOL>|13227,13228
breast|13228,13234
hematoma|13235,13243
)|13243,13244
<EOL>|13244,13245
<EOL>|13245,13246
-|13246,13247
History|13248,13255
of|13256,13258
DVT|13259,13262
/|13262,13263
PE|13263,13265
,|13265,13266
antiphospholipid|13267,13283
antibody|13284,13292
syndrome|13293,13301
,|13301,13302
<EOL>|13303,13304
subtherapeutic|13304,13318
INR|13319,13322
:|13322,13323
<EOL>|13323,13324
[|13324,13325
]|13325,13326
F|13327,13328
/|13328,13329
u|13329,13330
_|13331,13332
_|13332,13333
_|13333,13334
clinic|13335,13341
on|13342,13344
_|13345,13346
_|13346,13347
_|13347,13348
.|13348,13349
Patient|13350,13357
can|13358,13361
continue|13362,13370
home|13371,13375
<EOL>|13376,13377
Warfarin|13377,13385
regimen|13386,13393
<EOL>|13393,13394
<EOL>|13395,13396
Medications|13396,13407
on|13408,13410
Admission|13411,13420
:|13420,13421
<EOL>|13421,13422
The|13422,13425
Preadmission|13426,13438
Medication|13439,13449
list|13450,13454
is|13455,13457
accurate|13458,13466
and|13467,13470
complete|13471,13479
.|13479,13480
<EOL>|13480,13481
1.|13481,13483
Atorvastatin|13484,13496
40|13497,13499
mg|13500,13502
PO|13503,13505
QPM|13506,13509
<EOL>|13510,13511
2.|13511,13513
Docusate|13514,13522
Sodium|13523,13529
100|13530,13533
mg|13534,13536
PO|13537,13539
BID|13540,13543
<EOL>|13544,13545
3.|13545,13547
Omeprazole|13548,13558
20|13559,13561
mg|13562,13564
PO|13565,13567
BID|13568,13571
<EOL>|13572,13573
4.|13573,13575
Senna|13576,13581
8.6|13582,13585
mg|13586,13588
PO|13589,13591
HS|13592,13594
<EOL>|13595,13596
5.|13596,13598
Sertraline|13599,13609
150|13610,13613
mg|13614,13616
PO|13617,13619
DAILY|13620,13625
<EOL>|13626,13627
6.|13627,13629
TraZODone|13630,13639
50|13640,13642
mg|13643,13645
PO|13646,13648
QHS|13649,13652
:|13652,13653
PRN|13653,13656
sleep|13657,13662
<EOL>|13663,13664
7.|13664,13666
TraMADol|13667,13675
50|13676,13678
mg|13679,13681
PO|13682,13684
Q8H|13685,13688
:|13688,13689
PRN|13689,13692
Pain|13693,13697
-|13698,13699
Moderate|13700,13708
<EOL>|13709,13710
Reason|13712,13718
for|13719,13722
PRN|13723,13726
duplicate|13727,13736
override|13737,13745
:|13745,13746
Alternating|13747,13758
agents|13759,13765
for|13766,13769
<EOL>|13770,13771
similar|13771,13778
severity|13779,13787
<EOL>|13787,13788
8.|13788,13790
Polyethylene|13791,13803
Glycol|13804,13810
17|13811,13813
g|13814,13815
PO|13816,13818
DAILY|13819,13824
:|13824,13825
PRN|13825,13828
Constipation|13829,13841
-|13842,13843
First|13844,13849
<EOL>|13850,13851
Line|13851,13855
<EOL>|13856,13857
9.|13857,13859
ProAir|13860,13866
HFA|13867,13870
(|13871,13872
albuterol|13872,13881
sulfate|13882,13889
)|13889,13890
90|13891,13893
mcg|13894,13897
/|13897,13898
actuation|13898,13907
inhalation|13908,13918
<EOL>|13919,13920
Q4H|13920,13923
:|13923,13924
PRN|13924,13927
<EOL>|13928,13929
10.|13929,13932
Acetaminophen|13933,13946
1000|13947,13951
mg|13952,13954
PO|13955,13957
Q8H|13958,13961
:|13961,13962
PRN|13962,13965
Pain|13966,13970
-|13971,13972
Mild|13973,13977
/|13977,13978
Fever|13978,13983
<EOL>|13984,13985
11.|13985,13988
Albuterol|13989,13998
0.083|13999,14004
%|14004,14005
Neb|14006,14009
Soln|14010,14014
1|14015,14016
NEB|14017,14020
IH|14021,14023
Q6H|14024,14027
:|14027,14028
PRN|14028,14031
cough|14032,14037
,|14037,14038
wheeze|14039,14045
<EOL>|14046,14047
12.|14047,14050
Vitamin|14051,14058
D|14059,14060
_|14061,14062
_|14062,14063
_|14063,14064
UNIT|14065,14069
PO|14070,14072
DAILY|14073,14078
<EOL>|14079,14080
13.|14080,14083
Erythromycin|14084,14096
0.5|14097,14100
%|14100,14101
Ophth|14102,14107
Oint|14108,14112
0.5|14113,14116
in|14117,14119
BOTH|14120,14124
EYES|14125,14129
QID|14130,14133
<EOL>|14134,14135
14.|14135,14138
Furosemide|14139,14149
20|14150,14152
mg|14153,14155
PO|14156,14158
DAILY|14159,14164
:|14164,14165
PRN|14165,14168
Leg|14169,14172
swelling|14173,14181
<EOL>|14182,14183
15.|14183,14186
HYDROmorphone|14187,14200
(|14201,14202
Dilaudid|14202,14210
)|14210,14211
2|14212,14213
mg|14214,14216
PO|14217,14219
Q4H|14220,14223
:|14223,14224
PRN|14224,14227
Pain|14228,14232
-|14233,14234
Severe|14235,14241
<EOL>|14242,14243
16|14243,14245
.|14245,14246
Warfarin|14247,14255
7.5|14256,14259
mg|14260,14262
PO|14263,14265
2X|14266,14268
/|14268,14269
WEEK|14269,14273
(|14274,14275
_|14275,14276
_|14276,14277
_|14277,14278
)|14278,14279
<EOL>|14280,14281
17.|14281,14284
Warfarin|14285,14293
5|14294,14295
mg|14296,14298
PO|14299,14301
5X|14302,14304
/|14304,14305
WEEK|14305,14309
(|14310,14311
_|14311,14312
_|14312,14313
_|14313,14314
)|14314,14315
<EOL>|14316,14317
<EOL>|14317,14318
<EOL>|14319,14320
Discharge|14320,14329
Medications|14330,14341
:|14341,14342
<EOL>|14342,14343
1.|14343,14345
Gabapentin|14347,14357
600|14358,14361
mg|14362,14364
PO|14365,14367
TID|14368,14371
<EOL>|14372,14373
RX|14373,14375
*|14376,14377
gabapentin|14377,14387
600|14388,14391
mg|14392,14394
1|14395,14396
tablet|14397,14403
(|14403,14404
s|14404,14405
)|14405,14406
by|14407,14409
mouth|14410,14415
three|14416,14421
times|14422,14427
daily|14428,14433
<EOL>|14434,14435
Disp|14435,14439
#|14440,14441
*|14441,14442
90|14442,14444
Tablet|14445,14451
Refills|14452,14459
:|14459,14460
*|14460,14461
0|14461,14462
<EOL>|14463,14464
2.|14464,14466
Lidocaine|14468,14477
5|14478,14479
%|14479,14480
Patch|14481,14486
1|14487,14488
PTCH|14489,14493
TD|14494,14496
QAM|14497,14500
right|14501,14506
hip|14507,14510
<EOL>|14511,14512
RX|14512,14514
*|14515,14516
lidocaine|14516,14525
5|14526,14527
%|14528,14529
Apply|14530,14535
_|14536,14537
_|14537,14538
_|14538,14539
patches|14540,14547
daily|14548,14553
Disp|14554,14558
#|14559,14560
*|14560,14561
12|14561,14563
Patch|14564,14569
<EOL>|14570,14571
Refills|14571,14578
:|14578,14579
*|14579,14580
0|14580,14581
<EOL>|14582,14583
3.|14583,14585
TraMADol|14587,14595
50|14596,14598
mg|14599,14601
PO|14602,14604
Q6H|14605,14608
:|14608,14609
PRN|14609,14612
Pain|14613,14617
-|14618,14619
Moderate|14620,14628
<EOL>|14629,14630
RX|14630,14632
*|14633,14634
tramadol|14634,14642
50|14643,14645
mg|14646,14648
1|14649,14650
tablet|14651,14657
(|14657,14658
s|14658,14659
)|14659,14660
by|14661,14663
mouth|14664,14669
Every|14670,14675
six|14676,14679
hours|14680,14685
as|14686,14688
<EOL>|14689,14690
needed|14690,14696
Disp|14697,14701
#|14702,14703
*|14703,14704
15|14704,14706
Tablet|14707,14713
Refills|14714,14721
:|14721,14722
*|14722,14723
0|14723,14724
<EOL>|14725,14726
4.|14726,14728
Acetaminophen|14730,14743
1000|14744,14748
mg|14749,14751
PO|14752,14754
Q8H|14755,14758
:|14758,14759
PRN|14759,14762
Pain|14763,14767
-|14768,14769
Mild|14770,14774
/|14774,14775
Fever|14775,14780
<EOL>|14782,14783
5.|14783,14785
Albuterol|14787,14796
0.083|14797,14802
%|14802,14803
Neb|14804,14807
Soln|14808,14812
1|14813,14814
NEB|14815,14818
IH|14819,14821
Q6H|14822,14825
:|14825,14826
PRN|14826,14829
cough|14830,14835
,|14835,14836
wheeze|14837,14843
<EOL>|14845,14846
6.|14846,14848
Atorvastatin|14850,14862
40|14863,14865
mg|14866,14868
PO|14869,14871
QPM|14872,14875
<EOL>|14877,14878
7.|14878,14880
Docusate|14882,14890
Sodium|14891,14897
100|14898,14901
mg|14902,14904
PO|14905,14907
BID|14908,14911
<EOL>|14913,14914
8.|14914,14916
Erythromycin|14918,14930
0.5|14931,14934
%|14934,14935
Ophth|14936,14941
Oint|14942,14946
0.5|14947,14950
in|14951,14953
BOTH|14954,14958
EYES|14959,14963
QID|14964,14967
<EOL>|14969,14970
9.|14970,14972
Furosemide|14974,14984
20|14985,14987
mg|14988,14990
PO|14991,14993
DAILY|14994,14999
:|14999,15000
PRN|15000,15003
Leg|15004,15007
swelling|15008,15016
<EOL>|15018,15019
10.|15019,15022
Omeprazole|15024,15034
20|15035,15037
mg|15038,15040
PO|15041,15043
BID|15044,15047
<EOL>|15049,15050
11.|15050,15053
Polyethylene|15055,15067
Glycol|15068,15074
17|15075,15077
g|15078,15079
PO|15080,15082
DAILY|15083,15088
:|15088,15089
PRN|15089,15092
Constipation|15093,15105
-|15106,15107
First|15108,15113
<EOL>|15114,15115
Line|15115,15119
<EOL>|15121,15122
12.|15122,15125
ProAir|15127,15133
HFA|15134,15137
(|15138,15139
albuterol|15139,15148
sulfate|15149,15156
)|15156,15157
90|15158,15160
mcg|15161,15164
/|15164,15165
actuation|15165,15174
inhalation|15175,15185
<EOL>|15186,15187
Q4H|15187,15190
:|15190,15191
PRN|15191,15194
<EOL>|15196,15197
13.|15197,15200
Senna|15202,15207
8.6|15208,15211
mg|15212,15214
PO|15215,15217
HS|15218,15220
<EOL>|15222,15223
14.|15223,15226
Sertraline|15228,15238
150|15239,15242
mg|15243,15245
PO|15246,15248
DAILY|15249,15254
<EOL>|15256,15257
15.|15257,15260
TraZODone|15262,15271
50|15272,15274
mg|15275,15277
PO|15278,15280
QHS|15281,15284
:|15284,15285
PRN|15285,15288
sleep|15289,15294
<EOL>|15296,15297
16|15297,15299
.|15299,15300
Vitamin|15302,15309
D|15310,15311
_|15312,15313
_|15313,15314
_|15314,15315
UNIT|15316,15320
PO|15321,15323
DAILY|15324,15329
<EOL>|15331,15332
17.|15332,15335
Warfarin|15337,15345
5|15346,15347
mg|15348,15350
PO|15351,15353
2X|15354,15356
/|15356,15357
WEEK|15357,15361
(|15362,15363
_|15363,15364
_|15364,15365
_|15365,15366
)|15366,15367
<EOL>|15369,15370
18.|15370,15373
Warfarin|15375,15383
7.5|15384,15387
mg|15388,15390
PO|15391,15393
5X|15394,15396
/|15396,15397
WEEK|15397,15401
(|15402,15403
_|15403,15404
_|15404,15405
_|15405,15406
)|15406,15407
<EOL>|15409,15410
<EOL>|15410,15411
<EOL>|15412,15413
Discharge|15413,15422
Disposition|15423,15434
:|15434,15435
<EOL>|15435,15436
Home|15436,15440
With|15441,15445
Service|15446,15453
<EOL>|15453,15454
<EOL>|15455,15456
Facility|15456,15464
:|15464,15465
<EOL>|15465,15466
_|15466,15467
_|15467,15468
_|15468,15469
<EOL>|15469,15470
<EOL>|15471,15472
Discharge|15472,15481
Diagnosis|15482,15491
:|15491,15492
<EOL>|15492,15493
PRIMARY|15493,15500
:|15500,15501
<EOL>|15501,15502
=|15502,15503
=|15503,15504
=|15504,15505
=|15505,15506
=|15506,15507
=|15507,15508
=|15508,15509
=|15509,15510
=|15510,15511
=|15511,15512
=|15512,15513
=|15513,15514
=|15514,15515
=|15515,15516
=|15516,15517
=|15517,15518
=|15518,15519
<EOL>|15519,15520
Right|15520,15525
trochanteric|15526,15538
bursitis|15539,15547
<EOL>|15547,15548
Right|15548,15553
anterior|15554,15562
leg|15563,15566
pain|15567,15571
<EOL>|15571,15572
Right|15572,15577
sided|15578,15583
varicose|15584,15592
veins|15593,15598
<EOL>|15599,15600
<EOL>|15600,15601
SECONDARY|15601,15610
:|15610,15611
<EOL>|15611,15612
=|15612,15613
=|15613,15614
=|15614,15615
=|15615,15616
=|15616,15617
=|15617,15618
=|15618,15619
=|15619,15620
=|15620,15621
=|15621,15622
=|15622,15623
=|15623,15624
=|15624,15625
=|15625,15626
=|15626,15627
=|15627,15628
=|15628,15629
<EOL>|15629,15630
Iron|15630,15634
deficiency|15635,15645
anemia|15646,15652
<EOL>|15652,15653
History|15653,15660
of|15661,15663
DVT|15664,15667
/|15667,15668
PE|15668,15670
on|15671,15673
warfarin|15674,15682
<EOL>|15682,15683
Antiphospholipid|15683,15699
antibody|15700,15708
syndrome|15709,15717
<EOL>|15717,15718
Subtherapeutic|15718,15732
INR|15733,15736
<EOL>|15736,15737
Vitamin|15737,15744
D|15745,15746
deficiency|15747,15757
<EOL>|15757,15758
<EOL>|15758,15759
<EOL>|15760,15761
Discharge|15761,15770
Condition|15771,15780
:|15780,15781
<EOL>|15781,15782
Mental|15782,15788
Status|15789,15795
:|15795,15796
Clear|15797,15802
and|15803,15806
coherent|15807,15815
.|15815,15816
<EOL>|15816,15817
Level|15817,15822
of|15823,15825
Consciousness|15826,15839
:|15839,15840
Alert|15841,15846
and|15847,15850
interactive|15851,15862
.|15862,15863
<EOL>|15863,15864
Activity|15864,15872
Status|15873,15879
:|15879,15880
Ambulatory|15881,15891
-|15892,15893
requires|15894,15902
assistance|15903,15913
or|15914,15916
aid|15917,15920
(|15921,15922
walker|15922,15928
<EOL>|15929,15930
or|15930,15932
cane|15933,15937
)|15937,15938
.|15938,15939
<EOL>|15939,15940
<EOL>|15940,15941
<EOL>|15942,15943
Discharge|15943,15952
Instructions|15953,15965
:|15965,15966
<EOL>|15966,15967
Dear|15967,15971
_|15972,15973
_|15973,15974
_|15974,15975
,|15975,15976
<EOL>|15977,15978
<EOL>|15978,15979
You|15979,15982
were|15983,15987
admitted|15988,15996
because|15997,16004
you|16005,16008
were|16009,16013
having|16014,16020
a|16021,16022
lot|16023,16026
of|16027,16029
leg|16030,16033
pain|16034,16038
,|16038,16039
<EOL>|16040,16041
making|16041,16047
it|16048,16050
difficult|16051,16060
to|16061,16063
walk|16064,16068
.|16068,16069
<EOL>|16070,16071
<EOL>|16071,16072
In|16072,16074
the|16075,16078
hospital|16079,16087
,|16087,16088
we|16089,16091
gave|16092,16096
you|16097,16100
a|16101,16102
steroid|16103,16110
injection|16111,16120
near|16121,16125
your|16126,16130
right|16131,16136
<EOL>|16137,16138
thigh|16138,16143
for|16144,16147
a|16148,16149
condition|16150,16159
called|16160,16166
,|16166,16167
Trochanteric|16168,16180
Bursitis|16181,16189
.|16189,16190
We|16191,16193
also|16194,16198
<EOL>|16199,16200
gave|16200,16204
you|16205,16208
a|16209,16210
medication|16211,16221
called|16222,16228
Gabapentin|16229,16239
to|16240,16242
help|16243,16247
with|16248,16252
your|16253,16257
leg|16258,16261
<EOL>|16262,16263
pain|16263,16267
lower|16268,16273
down|16274,16278
.|16278,16279
<EOL>|16280,16281
<EOL>|16281,16282
We|16282,16284
also|16285,16289
started|16290,16297
you|16298,16301
on|16302,16304
a|16305,16306
medication|16307,16317
called|16318,16324
Lovenox|16325,16332
in|16333,16335
order|16336,16341
to|16342,16344
<EOL>|16345,16346
bridge|16346,16352
you|16353,16356
back|16357,16361
to|16362,16364
your|16365,16369
warfarin|16370,16378
-|16379,16380
currently|16381,16390
,|16390,16391
your|16392,16396
warfarin|16397,16405
dose|16406,16410
<EOL>|16411,16412
is|16412,16414
7.5|16415,16418
mg|16419,16421
daily|16422,16427
and|16428,16431
your|16432,16436
INR|16437,16440
was|16441,16444
1.9|16445,16448
at|16449,16451
discharge|16452,16461
(|16462,16463
goal|16463,16467
_|16468,16469
_|16469,16470
_|16470,16471
.|16471,16472
<EOL>|16473,16474
<EOL>|16474,16475
Finally|16475,16482
,|16482,16483
you|16484,16487
received|16488,16496
1|16497,16498
dose|16499,16503
of|16504,16506
intravenous|16507,16518
iron|16519,16523
because|16524,16531
you|16532,16535
are|16536,16539
<EOL>|16540,16541
iron|16541,16545
deficient|16546,16555
which|16556,16561
may|16562,16565
be|16566,16568
why|16569,16572
you|16573,16576
are|16577,16580
more|16581,16585
fatigued|16586,16594
than|16595,16599
<EOL>|16600,16601
usual|16601,16606
.|16606,16607
<EOL>|16607,16608
<EOL>|16608,16609
When|16609,16613
you|16614,16617
go|16618,16620
home|16621,16625
,|16625,16626
please|16627,16633
take|16634,16638
your|16639,16643
medications|16644,16655
as|16656,16658
prescribed|16659,16669
and|16670,16673
<EOL>|16674,16675
make|16675,16679
an|16680,16682
appointment|16683,16694
with|16695,16699
your|16700,16704
primary|16705,16712
care|16713,16717
doctor|16718,16724
.|16724,16725
We|16726,16728
do|16729,16731
not|16732,16735
<EOL>|16736,16737
know|16737,16741
what|16742,16746
exactly|16747,16754
is|16755,16757
causing|16758,16765
the|16766,16769
lower|16770,16775
leg|16776,16779
pain|16780,16784
,|16784,16785
so|16786,16788
you|16789,16792
may|16793,16796
want|16797,16801
<EOL>|16802,16803
to|16803,16805
talk|16806,16810
to|16811,16813
your|16814,16818
doctor|16819,16825
about|16826,16831
having|16832,16838
an|16839,16841
MRI|16842,16845
of|16846,16848
your|16849,16853
spine|16854,16859
.|16859,16860
You|16861,16864
<EOL>|16865,16866
can|16866,16869
also|16870,16874
ask|16875,16878
your|16879,16883
doctor|16884,16890
about|16891,16896
prescribing|16897,16908
a|16909,16910
medication|16911,16921
called|16922,16928
<EOL>|16929,16930
DICLOFENAC|16930,16940
GEL|16941,16944
,|16944,16945
also|16946,16950
called|16951,16957
VOLTAREN|16958,16966
.|16966,16967
This|16968,16972
is|16973,16975
essentially|16976,16987
Motrin|16988,16994
<EOL>|16995,16996
or|16996,16998
Advil|16999,17004
in|17005,17007
a|17008,17009
topical|17010,17017
form|17018,17022
and|17023,17026
may|17027,17030
help|17031,17035
your|17036,17040
pain|17041,17045
.|17045,17046
<EOL>|17046,17047
<EOL>|17047,17048
Additionally|17048,17060
,|17060,17061
please|17062,17068
talk|17069,17073
to|17074,17076
your|17077,17081
doctor|17082,17088
about|17089,17094
why|17095,17098
you|17099,17102
may|17103,17106
be|17107,17109
<EOL>|17110,17111
iron|17111,17115
deficient|17116,17125
.|17125,17126
<EOL>|17127,17128
<EOL>|17128,17129
It|17129,17131
was|17132,17135
a|17136,17137
pleasure|17138,17146
taking|17147,17153
part|17154,17158
in|17159,17161
your|17162,17166
care|17167,17171
.|17171,17172
We|17173,17175
wish|17176,17180
you|17181,17184
all|17185,17188
the|17189,17192
<EOL>|17193,17194
best|17194,17198
with|17199,17203
your|17204,17208
health|17209,17215
.|17215,17216
<EOL>|17216,17217
<EOL>|17217,17218
Sincerely|17218,17227
,|17227,17228
<EOL>|17228,17229
The|17229,17232
team|17233,17237
at|17238,17240
_|17241,17242
_|17242,17243
_|17243,17244
<EOL>|17244,17245
<EOL>|17245,17246
<EOL>|17247,17248
Followup|17248,17256
Instructions|17257,17269
:|17269,17270
<EOL>|17270,17271
_|17271,17272
_|17272,17273
_|17273,17274
<EOL>|17274,17275

