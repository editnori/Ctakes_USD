CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Morbid obesity|Disorder|false|false||Morbid obesitynull|Obesity|Disorder|false|false||obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|false|false||obesitynull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Laparoscopy|Procedure|false|false||Laparoscopicnull|Laparoscopic approach|Modifier|false|false||Laparoscopicnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Paraesophageal hernia|Disorder|false|false||paraesophageal hernianull|Paraesophageal|Modifier|false|false||paraesophagealnull|Hernia|Disorder|false|false||hernianull|Laparoscopic adjustable gastric banding|Procedure|false|false|C0038351|Laparoscopic adjustable gastric bandnull|Laparoscopy|Procedure|false|false||Laparoscopicnull|Laparoscopic approach|Modifier|false|false||Laparoscopicnull|Partitioning of stomach using band|Procedure|false|false|C0038351|gastric bandnull|Gastric band (physical object)|Device|false|false||gastric bandnull|Stomach|Anatomy|false|false|C1532765;C1960832|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Bands|Device|false|false||bandnull|Band form|Modifier|false|false||bandnull|Canadian Cardiovascular Society Grading of Angina Pectoris CCSGA101 Standardized Character Result Grade III|Finding|false|false||class III
null|Class 3|Finding|false|false||class IIInull|LOINC class types|Finding|false|false||class
null|Class|Finding|false|false||class
null|Classification|Finding|false|false||class
null|Taxonomic|Finding|false|false||class
null|Taxonomic Class|Finding|false|false||classnull|Kind of quantity - Class|LabModifier|false|false||classnull|Morbid obesity|Disorder|false|false||morbid obesitynull|Obesity|Disorder|false|false||obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|false|false||obesitynull|Pounds|LabModifier|false|false||poundsnull|Initial screening|Procedure|false|false||initial screennull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Toxicology screen, general (procedure)|Procedure|false|false||screen
null|Disease Screening|Procedure|false|false||screen
null|Screening for cancer|Procedure|false|false||screen
null|Screening procedure|Procedure|false|false||screennull|Screen Device|Device|false|false||screennull|Pounds|LabModifier|false|false||poundsnull|Height|LabModifier|false|false||heightnull|Inch Unit of Length|LabModifier|false|false||inchesnull|Finding of body mass index|Finding|false|false||BMInull|null|Attribute|false|false||BMI
null|Body mass index|Attribute|false|false||BMInull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Loss (adaptation)|Finding|false|false||Lossnull|Loss (quantitative)|LabModifier|false|false||Lossnull|PDLIM2 wt Allele|Finding|false|false||Slim
null|KLHDC10 gene|Finding|false|false||Slim
null|PDLIM2 gene|Finding|false|false||Slimnull|Fas-activated serine/threonine kinase activity|Finding|false|false||Fast
null|FASTK Gene|Finding|false|false||Fast
null|FOXD3-AS1 gene|Finding|false|false||Fast
null|FASTK wt Allele|Finding|false|false||Fast
null|Fasting|Finding|false|false||Fastnull|Rapid|Modifier|false|false||Fastnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|pancreatic lipase|Drug|false|false|C0030274|pancreatic lipase
null|pancreatic lipase|Drug|false|false|C0030274|pancreatic lipase
null|pancreatic lipase|Drug|false|false|C0030274|pancreatic lipase
null|PNLIP protein, human|Drug|false|false|C0030274|pancreatic lipase
null|PNLIP protein, human|Drug|false|false|C0030274|pancreatic lipasenull|PNLIP gene|Finding|false|false|C0030274|pancreatic lipasenull|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreaticnull|Pancreas|Anatomy|false|false|C1872737;C0443469;C0373670;C1418708;C0030292|pancreaticnull|lipase|Drug|false|false||lipase
null|lipase|Drug|false|false||lipase
null|lipase|Drug|false|false||lipasenull|Lipase measurement|Procedure|false|false|C0030274|lipasenull|Inhibitor|Drug|false|false||inhibitornull|Visit|Finding|false|false||visitsnull|Patient Visit|Procedure|false|false||visitsnull|20 pounds|Finding|false|false||20 poundsnull|Pounds|LabModifier|false|false||poundsnull|Unable|Finding|false|false||unablenull|Lowest|Modifier|false|false||lowestnull|Legal Adult|Subject|false|false||adult
null|Adult|Subject|false|false||adultnull|Pounds|LabModifier|false|false||poundsnull|Highest|Modifier|false|false||highestnull|Initial screening|Procedure|false|false||initial screennull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Toxicology screen, general (procedure)|Procedure|false|false||screen
null|Disease Screening|Procedure|false|false||screen
null|Screening for cancer|Procedure|false|false||screen
null|Screening procedure|Procedure|false|false||screennull|Screen Device|Device|false|false||screennull|Pounds|LabModifier|false|false||poundsnull|Pounds|LabModifier|false|false||poundsnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Pounds|LabModifier|false|false||poundsnull|One Year Ago|Modifier|false|false||one year agonull|One year|Time|false|false||one yearnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|year|Time|false|false||yearsnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|genetic aspects|Finding|false|false||genetics
null|Genetic|Finding|false|false||geneticsnull|genetics (procedure)|Procedure|false|false||geneticsnull|Science of genetics|Title|false|false||geneticsnull|Inconsistent|Modifier|false|false||inconsistentnull|Eating routine|Finding|false|false||meal patternnull|Meal (occasion for eating)|Finding|false|false||mealnull|Patterns|Modifier|false|false||patternnull|Late|Time|false|false||latenull|Night time|Time|false|false||nightnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Carbohydrates|Drug|false|false||carbohydrates
null|Carbohydrate nutrients|Drug|false|false||carbohydratesnull|Superficial abrasion|Disorder|false|false||grazingnull|Emotional Eating|Finding|false|false||emotional eatingnull|Emotional|Finding|false|false||emotional
null|Emotions|Finding|false|false||emotionalnull|Eating|Finding|false|false||eatingnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Hour|Time|false|false||hournull|times/week|LabModifier|false|false||times per weeknull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Weekly|Time|false|false||per weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Ellipse (shape)|Modifier|false|false||ellipticalnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|times/week|LabModifier|false|false||times per weeknull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Weekly|Time|false|false||per weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Bell Device|Device|false|false||bellnull|Processing ID - Training|Finding|false|false||trainingnull|Training Programs|Procedure|false|false||training
null|Training|Procedure|false|false||trainingnull|training aspects|Modifier|false|false||trainingnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Disease|Disorder|false|false||disordersnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|therapist|Subject|false|false||therapistnull|mental health|Finding|false|false||mental healthnull|null|Attribute|false|false||mental healthnull|Mental Health Specialty|Title|false|false||mental healthnull|Psyche structure|Finding|false|false||mentalnull|Health|Finding|false|false||healthnull|Psychotropic Drugs|Drug|true|false||psychotropicnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Triglycerides|Drug|false|false||triglyceride
null|Triglycerides|Drug|false|false||triglyceridenull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Deficiency anemias|Disorder|false|false||deficiency anemianull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Irritable Bowel Syndrome|Disorder|false|false|C0021853|irritable bowel syndromenull|Irritable Bowel Syndrome|Disorder|false|false|C0021853|irritable bowelnull|Irritable Mood|Finding|false|false||irritable
null|Irritability - emotion|Finding|false|false||irritablenull|Intestines|Anatomy|false|false|C0022104;C0022104|bowelnull|Syndrome|Disorder|false|false||syndromenull|Allergic rhinitis (disorder)|Disorder|false|false||allergic rhinitisnull|IL13 gene|Finding|false|false||allergic rhinitisnull|Allergic|Finding|false|false||allergicnull|Rhinitis|Disorder|false|false||rhinitisnull|Dysmenorrhea|Disorder|false|false||dysmenorrheanull|Vitamin D Deficiency|Disorder|false|false||vitamin D deficiencynull|Decreased circulating vitamin D concentration|Finding|false|false||vitamin D deficiencynull|Vitamin D Drug Class|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|D Vitamin|Drug|false|false||vitamin D
null|Vitamin D [EPC]|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|Vitamin D Drug Class|Drug|false|false||vitamin Dnull|Vitamin D measurement|Procedure|false|false||vitamin Dnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Suspected diagnosis|Modifier|false|false||question ofnull|Question (inquiry)|Finding|false|false||questionnull|Hypothyroidism|Disorder|false|false||hypothyroidismnull|Raised TSH level|Finding|false|false||elevated TSHnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Thyroid stimulating hormone measurement|Procedure|false|false||TSH levelnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Thalassemia trait|Disorder|false|false||thalassemia traitnull|Thalassemia|Disorder|false|false||thalassemianull|Trait|Subject|false|false||traitnull|Fatty Liver|Disorder|false|false|C4037986;C1278929;C0023884|fatty liver
null|Steatohepatitis|Disorder|false|false|C4037986;C1278929;C0023884|fatty livernull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0872387;C2711227;C0015695;C0023895;C0496870;C0577060;C0721399;C0023899|liver
null|null|Anatomy|false|false|C0872387;C2711227;C0015695;C0023895;C0496870;C0577060;C0721399;C0023899|liver
null|Liver|Anatomy|false|false|C0872387;C2711227;C0015695;C0023895;C0496870;C0577060;C0721399;C0023899|livernull|Cholelithiasis|Disorder|false|false||cholelithiasisnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Medical History|Finding|false|false|C0040421;C0836921|history ofnull|History of present illness (finding)|Finding|false|false|C0040421;C0836921|history
null|History of previous events|Finding|false|false|C0040421;C0836921|history
null|Historical aspects qualifier|Finding|false|false|C0040421;C0836921|history
null|Medical History|Finding|false|false|C0040421;C0836921|history
null|Concept History|Finding|false|false|C0040421;C0836921|historynull|History|Subject|false|false||historynull|examination of tonsils|Procedure|false|false|C0040421;C0836921|tonsilsnull|Palatine Tonsil|Anatomy|false|false|C2239123;C0262926;C0262926;C1705255;C0019665;C0262512;C2004062|tonsils
null|Tonsil|Anatomy|false|false|C2239123;C0262926;C0262926;C1705255;C0019665;C0262512;C2004062|tonsilsnull|Sleep Apnea, Obstructive|Disorder|false|false||obstructive sleep apneanull|Obstructed|Finding|false|false||obstructivenull|Sleep Apnea Syndromes|Disorder|false|false||sleep apneanull|SLEEP APNEA (device)|Device|false|false||sleep apneanull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Apnea|Finding|false|false||apneanull|Gastroesophageal reflux disease|Disorder|false|false|C0744316|gastroesophageal refluxnull|Infantile Gastroesophageal Reflux|Finding|false|false|C0744316|gastroesophageal reflux
null|Acid reflux|Finding|false|false|C0744316|gastroesophageal refluxnull|gastroesophageal|Anatomy|false|false|C3813607;C4317146;C0232483;C0017168|gastroesophagealnull|Reflux|Finding|false|false|C0744316|refluxnull|Completely Resolved|Finding|false|false||resolved completelynull|physiologic resolution|Finding|false|false||resolved
null|Resolution|Finding|false|false||resolvednull|Resolved|Modifier|false|false||resolvednull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Medical History|Finding|false|false|C4266530;C0029939;C0227898|History ofnull|History of present illness (finding)|Finding|false|false|C4266530;C0029939;C0227898|History
null|History of previous events|Finding|false|false|C4266530;C0029939;C0227898|History
null|Historical aspects qualifier|Finding|false|false|C4266530;C0029939;C0227898|History
null|Medical History|Finding|false|false|C4266530;C0029939;C0227898|History
null|Concept History|Finding|false|false|C4266530;C0029939;C0227898|Historynull|History|Subject|false|false||Historynull|Polycystic Ovary Syndrome|Disorder|false|false|C4266530;C0029939;C0227898|polycystic ovarynull|Polycystic|Modifier|false|false||polycysticnull|Neoplasm of uncertain or unknown behavior of ovary|Disorder|false|false|C4266530;C0029939;C0227898|ovary
null|Ovarian Diseases|Disorder|false|false|C4266530;C0029939;C0227898|ovarynull|Pelvis>Ovary|Anatomy|false|false|C0032460;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926;C0496920;C0029928|ovary
null|Ovary|Anatomy|false|false|C0032460;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926;C0496920;C0029928|ovary
null|Both ovaries|Anatomy|false|false|C0032460;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926;C0496920;C0029928|ovarynull|Syndrome|Disorder|false|false||syndromenull|Malignant neoplasm of urinary bladder|Disorder|false|false|C0005682|bladder CAnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0005684;C0872388|bladdernull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0567499;C0191838;C0007102;C0496956;C1882062;C0027651|breastnull|Neoplastic disease|Disorder|false|false|C0006141|neoplasia
null|Neoplasms|Disorder|false|false|C0006141|neoplasianull|Malignant tumor of colon|Disorder|false|false|C0006141;C0009368;C4071907|colon CAnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0007102|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0007102|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Ovarian|Anatomy|false|false||ovariannull|Sarcoma|Disorder|false|false||sarcoma
null|Malignant neoplasm of soft tissue|Disorder|false|false||sarcomanull|CONSTITUTIONAL PROBLEM|Finding|false|false||Constitutional
null|Constitutional|Finding|false|false||Constitutionalnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Lung|Anatomy|false|false||Lungsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Obesity|Disorder|false|false||Obesenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Appropriate|Modifier|false|false||appropriatenull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Traumatic Wound|Disorder|false|false||Woundsnull|Wounds - qualifier|Modifier|false|false||Woundsnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Site|Modifier|false|false||sitesnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|gusperimus|Drug|false|false||dsg
null|gusperimus|Drug|false|false||dsgnull|DSG1 wt Allele|Finding|false|false||dsg
null|DSG1 gene|Finding|false|false||dsgnull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|Serosanguineous|Modifier|false|false||serosanguinousnull|Staining (finding)|Finding|false|false||stainingnull|Staining method|Procedure|false|false||stainingnull|Periwound|Anatomy|false|false|C0041834|periwoundnull|Erythema|Disorder|true|false|C3534099|erythemanull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|uGy|LabModifier|false|false||UGInull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Slightly (qualifier value)|Modifier|false|false||Slightly
null|Slight (qualifier value)|Modifier|false|false||Slightlynull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Bands|Device|false|false||bandnull|Band form|Modifier|false|false||bandnull|Legal patent|Finding|false|false|C1955856|patentnull|Open|Modifier|false|false||patentnull|Surgical Stoma|Anatomy|false|false|C3887511;C0030650;C0332120;C0332234|stomanull|Evidence of (contextual qualifier)|Finding|true|false|C1955856|evidence ofnull|Evidence|Finding|true|false|C1955856|evidencenull|Leaking|Finding|true|false|C1955856|leaknull|Absence of sensation|Finding|false|false||anaesthesianull|Anesthesia procedures|Procedure|false|false||anaesthesianull|Anesthesiology|Title|false|false||anaesthesianull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Laparoscopic adjustable gastric banding|Procedure|false|false|C0038351|laparoscopic adjustable gastric bandnull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Partitioning of stomach using band|Procedure|false|false|C0038351|gastric bandnull|Gastric band (physical object)|Device|false|false||gastric bandnull|Stomach|Anatomy|false|false|C1960832;C1532765|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Bands|Device|false|false||bandnull|Band form|Modifier|false|false||bandnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Paraesophageal hernia|Disorder|false|false||paraesophageal hernianull|Paraesophageal|Modifier|false|false||paraesophagealnull|Hernia|Disorder|false|false||hernianull|Event|Event|false|false||eventsnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|null|Attribute|false|false||operative notenull|Operative|Time|false|false||operativenull|Details|Modifier|false|false||detailsnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Ward (environment)|Device|false|false||wardnull|Ward (person)|Subject|false|false||wardnull|Ward (environment)|Entity|false|false||wardnull|Examination and observation for unspecified reason|Finding|false|false||observation
null|null|Finding|false|false||observation
null|null|Finding|false|false||observation
null|Observation (finding)|Finding|false|false||observationnull|Observation - diagnostic procedure|Procedure|false|false||observation
null|Observation in research|Procedure|false|false||observation
null|Patient observation|Procedure|false|false||observationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Roxicet|Drug|false|false||Roxicet
null|Roxicet|Drug|false|false||Roxicetnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Cardiovascular and Pulmonary|Title|false|false||cardiovascular and pulmonarynull|Cardiovascular system|Anatomy|false|false||cardiovascular
null|Cardiovascular|Anatomy|false|false||cardiovascularnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|CENPJ gene|Finding|false|false||CPAPnull|Continuous Positive Airway Pressure|Procedure|false|false||CPAPnull|Overnight|Time|false|false||overnightnull|Known|Modifier|false|false||knownnull|Sleep Apnea Syndromes|Disorder|false|false||sleep apneanull|SLEEP APNEA (device)|Device|false|false||sleep apneanull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Apnea|Finding|false|false||apneanull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Initially|Time|false|false||initiallynull|Stage level 1|Finding|false|false||stage 1
null|Stage 1|Finding|false|false||stage 1null|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|TCF21 wt Allele|Finding|false|false||POD1
null|CORO7 gene|Finding|false|false||POD1
null|TCF21 gene|Finding|false|false||POD1null|uGy|LabModifier|false|false||UGInull|Series|LabModifier|false|false||seriesnull|uGy|LabModifier|false|false||UGInull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Leaking|Finding|true|false||leaknull|Obstruction|Finding|true|false||obstructionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Stage level 3|Finding|false|false||stage 3null|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Measuring intake and output|Procedure|false|false||intake and outputnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|monitoring of urine output for fluid balance|Procedure|false|false||Urine outputnull|null|Attribute|false|false||Urine output
null|null|Attribute|false|false||Urine outputnull|Urine volume finding|LabModifier|false|false||Urine outputnull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Hospitalization|Procedure|false|false||hospitalizationnull|subcutaneous heparin|Drug|false|false||subcutaneous heparin
null|subcutaneous heparin|Drug|false|false||subcutaneous heparinnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Boots|Device|false|false||bootsnull|Boots pharmaceutical company|Entity|false|false||bootsnull|During admission|Time|false|false||during admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Early|Time|false|false||earlynull|Frequently|Time|false|false||frequentnull|Ambulation|Finding|false|false||ambulation
null|Walking (function)|Finding|false|false||ambulationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|TCF21 wt Allele|Finding|false|false||POD1
null|CORO7 gene|Finding|false|false||POD1
null|TCF21 gene|Finding|false|false||POD1null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Teaching|Finding|false|false||teachingnull|Teaching aspects|Procedure|false|false||teaching
null|Education (procedure)|Procedure|false|false||teachingnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Comprehension|Finding|false|false||understandingnull|Agreement (document)|Finding|false|false||agreement
null|Agreement|Finding|false|false||agreementnull|null|Attribute|false|false||agreementnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Dietitian|Subject|false|false||dietitiannull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acidnull|Ascorbic acid measurement|Procedure|false|false||Ascorbic Acidnull|Daily|Time|false|false||DAILYnull|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferolnull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|Oralnull|Oral|Modifier|false|false||Oralnull|Daily|Time|false|false||dailynull|cyclobenzaprine|Drug|false|false||Cyclobenzaprine
null|cyclobenzaprine|Drug|false|false||Cyclobenzaprinenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false|C4083049;C0026845|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Spasm|Finding|false|false|C4083049;C0026845|muscle spasmsnull|Muscle (organ)|Anatomy|false|false|C1422467;C0037763|muscle
null|Muscle Tissue|Anatomy|false|false|C1422467;C0037763|musclenull|Spasm|Finding|false|false||spasmsnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|acetaminophen / oxycodone|Drug|false|false||OxycoDONE-Acetaminophennull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Elixir|Drug|false|false||Elixirnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|acetaminophen / oxycodone|Drug|false|false||oxycodone-acetaminophennull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Roxicet|Drug|false|false||Roxicet
null|Roxicet|Drug|false|false||Roxicetnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|milliliter|LabModifier|false|false||Milliliternull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|milliliter|LabModifier|false|false||Milliliternull|refill|Finding|false|false||Refillsnull|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acidnull|Ascorbic acid measurement|Procedure|false|false||Ascorbic Acidnull|Daily|Time|false|false||DAILYnull|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferolnull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|Oralnull|Oral|Modifier|false|false||Oralnull|Daily|Time|false|false||dailynull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Morbid obesity|Disorder|false|false||Morbid obesitynull|Obesity|Disorder|false|false||obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|false|false||obesitynull|Sleep Apnea, Obstructive|Disorder|false|false||Obstructive sleep apneanull|Obstructed|Finding|false|false||Obstructivenull|Sleep Apnea Syndromes|Disorder|false|false||sleep apneanull|SLEEP APNEA (device)|Device|false|false||sleep apneanull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Apnea|Finding|false|false||apneanull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||return tonull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Accident and Emergency department|Device|false|false||emergency departmentnull|interventional services emergency department|Entity|false|false||emergency department
null|Accident and Emergency department|Entity|false|false||emergency departmentnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Department - No suggested values defined|Finding|false|false||department
null|Organization Unit Type - Department|Finding|false|false||department
null|Department - Charge type|Finding|false|false||departmentnull|Department|Entity|false|false||departmentnull|Patient location type - Department|Modifier|false|false||department
null|Department - Person location type|Modifier|false|false||departmentnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Severe nausea|Finding|false|false||severe nauseanull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Abdominal bloating|Finding|false|false|C0000726|abdominal bloating
null|Abdomen distended|Finding|false|false|C0000726|abdominal bloatingnull|Abdomen|Anatomy|false|false|C1291077;C0000731|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Abdominal bloating|Finding|false|false||bloating
null|Abdomen distended|Finding|false|false||bloatingnull|Smell Perception|Finding|false|false||smellingnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical incisions|Procedure|false|false||incisionsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Surgical incisions|Procedure|false|false||incisionsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Advance [medical device]|Device|false|false||advancenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Cereal plant straw|Drug|false|false||strawnull|Straw package type|Device|false|false||strawnull|Straw Color|Modifier|false|false||strawnull|Straw (unit of presentation)|LabModifier|false|false||strawnull|Chew (administration method)|Finding|false|false||chew
null|Does chew (finding)|Finding|false|false||chew
null|Chewing|Finding|false|false||chewnull|Gum as an ingredient|Drug|false|false|C0017562|gum
null|Gum Dose Form|Drug|false|false|C0017562|gumnull|OTULIN wt Allele|Finding|false|false|C0017562|gum
null|OTULIN gene|Finding|false|false|C0017562|gumnull|Gingiva|Anatomy|false|false|C5444202;C1825233;C0812395;C1378701|gumnull|Gum - unit of product usage|LabModifier|false|false||gum
null|Gum Dosing Unit|LabModifier|false|false||gumnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|cyclobenzaprine|Drug|false|false||cyclobenzaprine
null|cyclobenzaprine|Drug|false|false||cyclobenzaprinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Crushing (procedure)|Procedure|false|false||CRUSHnull|Pills|Drug|false|false||PILLSnull|New medications|Drug|false|false||new medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Drowsiness|Finding|false|false||drowsynull|Ability Question|Finding|false|false||ability tonull|Oral Intake Ability|Finding|false|false||abilitynull|Ability|Subject|false|false||abilitynull|Motor Vehicles|Device|false|false||motor vehiclenull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Drug vehicle|Drug|false|false||vehiclenull|Vehicle (transportation)|Device|false|false||vehiclenull|operate|Finding|false|false||operatenull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Minerals|Drug|false|false||mineralsnull|Chewable Gel Dosing Unit|LabModifier|false|false||gummynull|VITAMINS [VA Class]|Drug|true|false||vitamins
null|Vitamin IV solution additives|Drug|true|false||vitamins
null|Vitamins|Drug|true|false||vitamins
null|Vitamins|Drug|true|false||vitamins
null|Vitamins|Drug|true|false||vitaminsnull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Constipation|Finding|false|false||constipationnull|Intestines|Anatomy|false|false||bowelnull|Patterns|Modifier|false|false||patternnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|false|false||NSAIDS
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDSnull|Anti-Inflammatory Agents|Drug|false|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|false|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|false|false||drugsnull|Drugs - dental services|Procedure|false|false||drugsnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|Aleve|Drug|false|false||Aleve
null|Aleve|Drug|false|false||Alevenull|Nuprin|Drug|false|false||Nuprin
null|Nuprin|Drug|false|false||Nuprinnull|naproxen|Drug|false|false||Naproxen
null|naproxen|Drug|false|false||Naproxennull|Hemorrhage|Finding|false|false||bleedingnull|Ulcer|Finding|false|false||ulcersnull|Gastrointestinal system|Anatomy|false|false|C0012238;C5671121;C0449913;C5441654|digestive systemnull|Digestion|Finding|false|false|C0012240;C0012240|digestivenull|Gastrointestinal system|Anatomy|false|false|C0012238;C0449913;C5441654|digestivenull|System (basic dose form)|Drug|false|false|C0012240|systemnull|System, LOINC Axis 4|Finding|false|false|C0012240;C0012240|system
null|System|Finding|false|false|C0012240;C0012240|systemnull|Device system|Device|false|false||system
null|System - kit|Device|false|false||systemnull|System (unit of presentation)|LabModifier|false|false||systemnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|true|false||liftingnull|Pounds|LabModifier|false|false||poundsnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Moderate Exercise|Finding|false|false||moderate exercisenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Discretion|Finding|false|false||discretionnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Exercise|Finding|false|false||exercisesnull|Physical therapy exercises|Procedure|false|false||exercisesnull|Wound care management|Procedure|false|false||Wound Care
null|wound care|Procedure|false|false||Wound Carenull|Wound Care kit|Device|false|false||Wound Carenull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|TUB gene|Finding|true|false||tubnull|Tub - container|Device|true|false||tubnull|Tub Dosing Unit|LabModifier|false|false||tubnull|Bathing|Procedure|true|false||bathsnull|Baths (medical device)|Device|true|false||bathsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical incisions|Procedure|false|false||incisionsnull|null|Finding|false|false||covernull|Cover (physical object)|Device|false|false||cover
null|Cover Device|Device|false|false||covernull|Cleaning (activity)|Event|false|false||cleannull|Gauzes|Device|false|false||gauzenull|Steri-Strip|Device|false|false||steri-stripsnull|Silene|Entity|false|false||sterinull|strip medical device|Device|false|false||stripsnull|Own|Finding|false|false||ownnull|strip medical device|Device|false|false||stripsnull|day|Time|false|false||daysnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Site of incision|Modifier|false|false||incision sitesnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Site|Modifier|false|false||sitesnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions