 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|165,174|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|165,174|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|165,174|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|177,182|false|false|false|C0749139|sulfa|Sulfa
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|184,196|false|false|false|C0161497;C2876788|Poisoning by sulfonamide;Poisoning by, adverse effect of and underdosing of sulfonamides|Sulfonamides
Drug|Antibiotic|SIMPLE_SEGMENT|184,196|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Drug|Organic Chemical|SIMPLE_SEGMENT|184,196|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|184,196|false|false|false|C0038760;C0599503;C3539179;C3539184;C3541962;C3541963|Sulfonamide Anti-Infective Agents;Sulfonamides;Sulfonamides, Gynecological;Sulfonamides, intestinal antiinfectives;Sulfonamides, ophthalmologic antiinfectives;Sulfonamides, topical|Sulfonamides
Event|Event|SIMPLE_SEGMENT|184,196|false|false|false|||Sulfonamides
Finding|Pathologic Function|SIMPLE_SEGMENT|184,196|false|false|false|C0261773|Adverse reaction to sulfonamides|Sulfonamides
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|200,211|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|200,211|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|200,211|false|false|false|C0030842|penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|200,211|false|false|false|||Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|200,211|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|214,223|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|214,223|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|231,246|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|237,246|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|237,246|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|237,246|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|248,254|false|false|false|C0015450|Face|Facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|248,263|false|false|false|C0427055|Facial Paresis|Facial weakness
Event|Event|SIMPLE_SEGMENT|255,263|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|255,263|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Classification|SIMPLE_SEGMENT|266,271|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|272,280|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|272,280|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|284,302|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|293,302|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|293,302|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|293,302|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|293,302|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|293,302|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|311,318|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|311,318|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|311,318|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|311,318|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|311,321|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|311,337|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|311,337|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|322,329|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|322,329|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|322,337|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|330,337|true|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|339,342|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|339,342|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|339,342|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|339,342|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|348,351|false|false|false|C0228528|Rhomboid fossa structure|RHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|358,362|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|358,362|false|false|false|||GERD
Finding|Intellectual Product|SIMPLE_SEGMENT|364,368|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|364,379|false|false|false|C0588006|Mild depression|mild depression
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|369,379|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|369,379|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|369,379|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|369,379|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|391,400|false|false|false|C0149931|Migraine Disorders|migraines
Event|Event|SIMPLE_SEGMENT|391,400|false|false|false|||migraines
Event|Event|SIMPLE_SEGMENT|402,410|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|420,427|false|false|false|||episode
Anatomy|Body Location or Region|SIMPLE_SEGMENT|431,437|false|false|false|C0015450|Face|facial
Finding|Sign or Symptom|SIMPLE_SEGMENT|431,446|false|false|false|C0239511|Numbness of face|facial numbness
Event|Event|SIMPLE_SEGMENT|438,446|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|438,446|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|438,446|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|461,466|false|false|false|||lying
Finding|Functional Concept|SIMPLE_SEGMENT|474,478|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|479,483|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|479,483|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|479,483|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|479,483|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|485,493|false|false|false|||watching
Finding|Mental Process|SIMPLE_SEGMENT|485,493|false|false|false|C2371283|Watching|watching
Finding|Intellectual Product|SIMPLE_SEGMENT|485,496|false|false|false|C3827501|Watching TV|watching TV
Event|Event|SIMPLE_SEGMENT|494,496|false|false|false|||TV
Event|Event|SIMPLE_SEGMENT|502,509|false|false|false|||noticed
Finding|Functional Concept|SIMPLE_SEGMENT|535,539|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|540,544|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|540,544|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|540,544|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|540,544|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|549,553|false|false|false|||numb
Finding|Gene or Genome|SIMPLE_SEGMENT|549,553|false|false|false|C1417890;C1709287|NUMB gene;Numb (emotional response)|numb
Finding|Individual Behavior|SIMPLE_SEGMENT|549,553|false|false|false|C1417890;C1709287|NUMB gene;Numb (emotional response)|numb
Event|Event|SIMPLE_SEGMENT|569,577|false|false|false|||injected
Event|Event|SIMPLE_SEGMENT|600,612|false|false|false|||distribution
Finding|Cell Function|SIMPLE_SEGMENT|600,612|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|SIMPLE_SEGMENT|600,612|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Event|Event|SIMPLE_SEGMENT|622,628|false|false|false|||traces
Event|Event|SIMPLE_SEGMENT|635,641|false|false|false|||mid-V2
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|654,657|false|false|false|C0022359|Jaw|jaw
Drug|Biologically Active Substance|SIMPLE_SEGMENT|659,663|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|659,663|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|659,663|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|659,663|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|659,663|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|679,686|false|false|false|||thought
Event|Event|SIMPLE_SEGMENT|714,719|false|false|false|||lying
Event|Event|SIMPLE_SEGMENT|732,741|false|false|false|||concerned
Event|Event|SIMPLE_SEGMENT|750,759|false|false|false|||persisted
Event|Event|SIMPLE_SEGMENT|765,773|false|false|false|||endorsed
Finding|Intellectual Product|SIMPLE_SEGMENT|776,780|true|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|781,788|true|false|false|||diffuse
Finding|Sign or Symptom|SIMPLE_SEGMENT|789,793|true|false|false|C0278144|Dull pain|dull
Event|Event|SIMPLE_SEGMENT|809,816|true|false|false|||unusual
Event|Event|SIMPLE_SEGMENT|830,836|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|854,858|false|false|false|||felt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|871,879|false|false|false|C0149931|Migraine Disorders|migraine
Event|Event|SIMPLE_SEGMENT|871,879|false|false|false|||migraine
Event|Event|SIMPLE_SEGMENT|885,891|false|false|false|||coming
Event|Event|SIMPLE_SEGMENT|926,933|true|false|false|||typical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|946,955|true|false|false|C0149931|Migraine Disorders|migraines
Event|Event|SIMPLE_SEGMENT|946,955|true|false|false|||migraines
Event|Event|SIMPLE_SEGMENT|961,969|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|961,969|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|961,969|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|970,976|false|false|false|||lasted
Event|Event|SIMPLE_SEGMENT|980,987|false|false|false|||minutes
Event|Event|SIMPLE_SEGMENT|1001,1009|false|false|false|||resolved
Finding|Intellectual Product|SIMPLE_SEGMENT|1010,1020|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|1047,1055|true|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1047,1055|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|1068,1075|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1068,1075|true|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1091,1095|true|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1091,1095|true|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|1091,1095|true|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|1091,1095|true|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1105,1112|true|false|false|C1135208|Vertigo as late effect of cerebrovascular disease|vertigo
Event|Event|SIMPLE_SEGMENT|1105,1112|true|false|false|||vertigo
Finding|Sign or Symptom|SIMPLE_SEGMENT|1105,1112|true|false|false|C0042571|Vertigo|vertigo
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1117,1125|false|false|false|C2706915||language
Finding|Intellectual Product|SIMPLE_SEGMENT|1117,1125|false|false|false|C0033348|Programming Languages|language
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1117,1136|false|false|false|C0023015|Language Disorders|language impairment
Event|Event|SIMPLE_SEGMENT|1126,1136|false|false|false|||impairment
Finding|Finding|SIMPLE_SEGMENT|1126,1136|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|SIMPLE_SEGMENT|1126,1136|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Event|Event|SIMPLE_SEGMENT|1149,1155|true|false|false|||recall
Event|Event|SIMPLE_SEGMENT|1176,1185|true|false|false|||happening
Event|Event|SIMPLE_SEGMENT|1198,1204|false|false|false|||states
Finding|Idea or Concept|SIMPLE_SEGMENT|1214,1217|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1214,1217|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1232,1239|false|false|false|||routine
Finding|Idea or Concept|SIMPLE_SEGMENT|1232,1239|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|SIMPLE_SEGMENT|1232,1239|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1232,1239|false|false|false|C1979801|Routine coag|routine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1244,1247|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1244,1247|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1244,1247|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|SIMPLE_SEGMENT|1244,1247|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1244,1247|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|SIMPLE_SEGMENT|1244,1247|false|false|false|||ROS
Finding|Gene or Genome|SIMPLE_SEGMENT|1244,1247|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|SIMPLE_SEGMENT|1244,1247|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|SIMPLE_SEGMENT|1253,1258|false|false|false|||notes
Finding|Gene or Genome|SIMPLE_SEGMENT|1278,1281|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|1290,1298|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1290,1298|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1290,1298|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Intellectual Product|SIMPLE_SEGMENT|1305,1309|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|1316,1324|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|1349,1357|false|false|false|||endorses
Event|Event|SIMPLE_SEGMENT|1358,1365|false|false|false|||feeling
Finding|Mental Process|SIMPLE_SEGMENT|1358,1365|false|false|false|C1527305|Feelings|feeling
Finding|Gene or Genome|SIMPLE_SEGMENT|1381,1384|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|1401,1407|false|false|false|||health
Finding|Idea or Concept|SIMPLE_SEGMENT|1401,1407|false|false|false|C0018684|Health|health
Event|Event|SIMPLE_SEGMENT|1417,1423|false|false|false|||normal
Finding|Finding|SIMPLE_SEGMENT|1429,1449|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1434,1441|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1434,1441|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1434,1441|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1434,1441|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1434,1441|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1434,1449|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1442,1449|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1442,1449|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1442,1449|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1451,1455|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|1451,1455|false|false|false|||GERD
Finding|Intellectual Product|SIMPLE_SEGMENT|1457,1461|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1457,1472|false|false|false|C0588006|Mild depression|mild depression
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1462,1472|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|1462,1472|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|1462,1472|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|1462,1472|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1473,1482|false|false|false|C0149931|Migraine Disorders|migraines
Event|Event|SIMPLE_SEGMENT|1473,1482|false|false|false|||migraines
Finding|Mental Process|SIMPLE_SEGMENT|1498,1503|false|false|false|C0004083|Mental association|assoc
Finding|Functional Concept|SIMPLE_SEGMENT|1509,1515|false|false|false|C0234621|Visual|visual
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1509,1523|false|false|false|C0085635|Photopsia|visual flashes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1516,1523|false|false|false|C0085635|Photopsia|flashes
Event|Event|SIMPLE_SEGMENT|1516,1523|false|false|false|||flashes
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1516,1523|false|false|false|C0542555|Natural flashes|flashes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1516,1532|false|false|false|C0085635|Photopsia|flashes of light
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1527,1532|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1527,1532|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|1527,1532|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|1527,1532|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|1527,1532|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|1527,1532|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1527,1532|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1527,1532|false|false|false|C0031765|Phototherapy|light
Finding|Gene or Genome|SIMPLE_SEGMENT|1550,1553|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|1555,1562|false|false|false|C0006386|Bunion|bunions
Event|Event|SIMPLE_SEGMENT|1555,1562|false|false|false|||bunions
Finding|Functional Concept|SIMPLE_SEGMENT|1565,1571|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1565,1579|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1572,1579|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1572,1579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1572,1579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1572,1579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1585,1591|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1585,1591|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1585,1591|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1585,1591|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1585,1599|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1592,1599|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1592,1599|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1592,1599|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1592,1599|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1601,1607|false|false|false|||Father
Finding|Conceptual Entity|SIMPLE_SEGMENT|1601,1607|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1601,1607|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|1617,1626|false|false|false|||sustained
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1629,1635|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1629,1635|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1629,1635|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1644,1651|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|1644,1651|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1644,1656|false|false|false|C0018795|Cardiac Catheterization Procedures|cardiac cath
Event|Event|SIMPLE_SEGMENT|1652,1656|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1652,1656|false|false|false|C0007430|Catheterization|cath
Finding|Idea or Concept|SIMPLE_SEGMENT|1668,1672|false|false|false|C0376558|Life|life
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1668,1672|false|false|false|C1522684|Laser-Induced Fluorescence Endoscopy|life
Event|Event|SIMPLE_SEGMENT|1673,1679|false|false|false|||father
Finding|Conceptual Entity|SIMPLE_SEGMENT|1673,1679|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|1673,1679|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|SIMPLE_SEGMENT|1680,1689|false|false|false|||developed
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1692,1702|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|SIMPLE_SEGMENT|1692,1702|false|false|false|||meningioma
Event|Event|SIMPLE_SEGMENT|1718,1726|false|false|false|||seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|1718,1726|false|false|false|C0036572|Seizures|seizures
Event|Event|SIMPLE_SEGMENT|1732,1740|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1732,1740|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1732,1740|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1732,1740|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1732,1745|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1732,1745|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1741,1745|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1741,1745|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1741,1745|false|false|false|C0582103|Medical Examination|Exam
Finding|Classification|SIMPLE_SEGMENT|1775,1778|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|1775,1778|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|1780,1785|false|false|false|||Lying
Finding|Individual Behavior|SIMPLE_SEGMENT|1780,1785|false|false|false|C0600261|Telling untruths|Lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1789,1792|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|1789,1792|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|1789,1792|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1794,1797|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1794,1797|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1794,1797|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1794,1797|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1794,1797|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1794,1797|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1794,1797|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1798,1803|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|1812,1829|false|false|false|C0455900|Moist oral mucosa|moist oral mucosa
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1818,1822|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1818,1822|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|1818,1822|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|1818,1822|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1818,1829|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|1823,1829|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|1823,1829|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1833,1837|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|1833,1837|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|1833,1837|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|1842,1852|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|1842,1852|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1842,1852|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|1856,1865|true|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1856,1865|true|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|1874,1877|true|false|false|||ROM
Finding|Finding|SIMPLE_SEGMENT|1874,1877|true|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|SIMPLE_SEGMENT|1874,1877|true|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1874,1877|true|false|false|C1562926|Range of motion technique (procedure)|ROM
Event|Event|SIMPLE_SEGMENT|1879,1885|true|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|1879,1885|true|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1890,1897|true|false|false|C0007272|Carotid Arteries|carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1901,1910|true|false|false|C0549207|Bone structure of spine|vertebral
Event|Event|SIMPLE_SEGMENT|1911,1916|true|false|false|||bruit
Finding|Finding|SIMPLE_SEGMENT|1911,1916|true|false|false|C0006318|Bruit|bruit
Event|Event|SIMPLE_SEGMENT|1921,1924|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1943,1950|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|1943,1950|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|1959,1963|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|1959,1963|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1965,1969|true|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1965,1969|true|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1965,1969|true|false|false|C0024115|Lung diseases|Lung
Event|Event|SIMPLE_SEGMENT|1965,1969|true|false|false|||Lung
Finding|Finding|SIMPLE_SEGMENT|1965,1969|true|false|false|C0740941|Lung Problem|Lung
Event|Event|SIMPLE_SEGMENT|1971,1976|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|1971,1976|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|1980,1992|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1980,1992|false|false|false|C0004339|Auscultation|auscultation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2006,2009|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|aBd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2006,2009|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|aBd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2015,2019|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2015,2019|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2021,2030|false|false|false|||nontender
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2032,2035|false|false|false|C0015306|Hereditary Multiple Exostoses|ext
Event|Event|SIMPLE_SEGMENT|2032,2035|false|false|false|||ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2032,2035|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|ext
Finding|Intellectual Product|SIMPLE_SEGMENT|2047,2052|false|false|false|C1549782|Relational Operator - Equal|equal
Event|Event|SIMPLE_SEGMENT|2053,2059|false|false|false|||radial
Finding|Conceptual Entity|SIMPLE_SEGMENT|2053,2059|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2064,2069|false|false|false|C0016504;C0687080|Foot;Paw|pedal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2064,2076|false|false|false|C0232157|Pedal pulse|pedal pulses
Drug|Food|SIMPLE_SEGMENT|2070,2076|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2070,2076|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2070,2076|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2070,2076|false|false|false|C0034107|Pulse taking|pulses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2086,2108|false|false|false|C0027853|Neurologic Examination|Neurologic examination
Event|Activity|SIMPLE_SEGMENT|2097,2108|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|2097,2108|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|2097,2108|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Finding|Mental Process|SIMPLE_SEGMENT|2111,2117|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2111,2124|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|SIMPLE_SEGMENT|2111,2124|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2118,2124|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|2118,2124|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|2118,2124|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|2126,2131|false|false|false|||Awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2136,2141|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2136,2141|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2136,2141|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2136,2141|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2136,2141|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2136,2141|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2136,2141|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|2143,2154|false|false|false|||cooperative
Event|Event|SIMPLE_SEGMENT|2160,2164|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2160,2164|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2160,2164|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|2166,2172|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|2174,2180|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|2174,2180|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|2174,2180|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|2183,2191|false|false|false|||Oriented
Finding|Finding|SIMPLE_SEGMENT|2183,2191|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|SIMPLE_SEGMENT|2183,2201|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2195,2201|false|false|false|C5890614||person
Event|Event|SIMPLE_SEGMENT|2195,2201|false|false|false|||person
Finding|Intellectual Product|SIMPLE_SEGMENT|2195,2201|false|false|false|C1522390|Person Info|person
Event|Activity|SIMPLE_SEGMENT|2203,2208|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|2203,2208|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|2203,2208|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|2203,2208|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|2241,2250|false|false|false|||backwards
Event|Event|SIMPLE_SEGMENT|2253,2259|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|2253,2259|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2253,2259|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|2263,2269|false|false|false|||fluent
Event|Event|SIMPLE_SEGMENT|2282,2295|false|false|false|||comprehension
Finding|Mental Process|SIMPLE_SEGMENT|2282,2295|false|false|false|C0162340|Comprehension|comprehension
Event|Event|SIMPLE_SEGMENT|2300,2310|false|false|false|||repetition
Finding|Finding|SIMPLE_SEGMENT|2300,2310|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|SIMPLE_SEGMENT|2300,2310|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|SIMPLE_SEGMENT|2312,2318|false|false|false|||naming
Event|Event|SIMPLE_SEGMENT|2319,2325|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2319,2325|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2330,2340|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|SIMPLE_SEGMENT|2330,2340|true|false|false|||dysarthria
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2342,2349|false|false|false|C5890786||Reading
Finding|Conceptual Entity|SIMPLE_SEGMENT|2342,2349|false|false|false|C0034754;C1705179;C4284139|Reading (activity);Reading (datum presentation);Reading Ability question|Reading
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|2342,2349|false|false|false|C0034754;C1705179;C4284139|Reading (activity);Reading (datum presentation);Reading Ability question|Reading
Finding|Intellectual Product|SIMPLE_SEGMENT|2342,2349|false|false|false|C0034754;C1705179;C4284139|Reading (activity);Reading (datum presentation);Reading Ability question|Reading
Event|Event|SIMPLE_SEGMENT|2350,2356|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2350,2356|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|SIMPLE_SEGMENT|2361,2366|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|SIMPLE_SEGMENT|2367,2371|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2372,2381|true|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|2372,2381|true|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|2372,2381|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|2386,2394|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|2386,2394|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|2386,2397|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2398,2405|true|false|false|C0003635|Apraxias|apraxia
Event|Event|SIMPLE_SEGMENT|2398,2405|true|false|false|||apraxia
Event|Event|SIMPLE_SEGMENT|2409,2416|true|false|false|||neglect
Event|Event|SIMPLE_SEGMENT|2409,2416|true|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|SIMPLE_SEGMENT|2409,2416|true|false|false|C0521874|Victim of neglect (finding)|neglect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2420,2427|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2420,2434|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2420,2434|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2428,2434|false|false|false|C0027740|Nerve|Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2438,2444|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|2453,2458|false|false|false|||round
Event|Event|SIMPLE_SEGMENT|2463,2471|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2463,2471|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|SIMPLE_SEGMENT|2463,2480|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2475,2480|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2475,2480|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|2475,2480|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|2475,2480|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|2475,2480|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|2475,2480|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2475,2480|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2475,2480|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|SIMPLE_SEGMENT|2505,2511|false|false|false|C0234621|Visual|Visual
Event|Event|SIMPLE_SEGMENT|2512,2518|false|false|false|||fields
Event|Event|SIMPLE_SEGMENT|2523,2527|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|2531,2544|false|false|false|||confrontation
Finding|Finding|SIMPLE_SEGMENT|2531,2544|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2531,2544|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2531,2544|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2546,2553|false|false|false|C0035298|Retina|Retinas
Finding|Finding|SIMPLE_SEGMENT|2559,2564|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|SIMPLE_SEGMENT|2559,2564|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2565,2569|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|SIMPLE_SEGMENT|2565,2569|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2565,2569|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|SIMPLE_SEGMENT|2565,2569|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|SIMPLE_SEGMENT|2565,2569|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Event|Event|SIMPLE_SEGMENT|2570,2577|false|false|false|||margins
Finding|Functional Concept|SIMPLE_SEGMENT|2583,2594|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2583,2604|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|SIMPLE_SEGMENT|2595,2604|true|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2595,2604|true|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2605,2611|true|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2605,2611|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2628,2637|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|SIMPLE_SEGMENT|2628,2637|true|false|false|||nystagmus
Event|Event|SIMPLE_SEGMENT|2639,2648|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|2639,2648|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2639,2648|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2639,2648|false|false|false|C2229507|sensory exam|Sensation
Finding|Finding|SIMPLE_SEGMENT|2649,2655|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2682,2688|false|false|false|C0015450|Face|Facial
Event|Event|SIMPLE_SEGMENT|2689,2697|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2689,2697|false|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|2698,2707|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|2698,2707|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|2698,2707|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|2710,2717|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|2710,2717|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|SIMPLE_SEGMENT|2718,2724|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2718,2724|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2728,2734|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2753,2759|false|false|false|C0700374|Palate|Palate
Event|Event|SIMPLE_SEGMENT|2760,2769|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2760,2769|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|SIMPLE_SEGMENT|2770,2781|false|false|false|||symmetrical
Finding|Finding|SIMPLE_SEGMENT|2770,2781|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2784,2803|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2808,2817|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|SIMPLE_SEGMENT|2818,2824|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2838,2844|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2838,2844|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Event|Event|SIMPLE_SEGMENT|2838,2844|false|false|false|||Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|2838,2844|false|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|SIMPLE_SEGMENT|2838,2852|false|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|SIMPLE_SEGMENT|2845,2852|false|false|false|C1660780|midline cell component|midline
Event|Event|SIMPLE_SEGMENT|2854,2863|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2854,2863|false|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2864,2870|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2864,2870|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|2873,2878|false|false|false|||Motor
Finding|Functional Concept|SIMPLE_SEGMENT|2873,2878|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2888,2892|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|2888,2892|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|SIMPLE_SEGMENT|2888,2892|false|false|false|||bulk
Event|Event|SIMPLE_SEGMENT|2911,2917|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|2922,2930|true|false|false|||observed
Event|Event|SIMPLE_SEGMENT|2931,2940|true|false|false|||myoclonus
Finding|Finding|SIMPLE_SEGMENT|2931,2940|true|false|false|C0027066|Myoclonus|myoclonus
Event|Event|SIMPLE_SEGMENT|2944,2950|true|false|false|||tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|2944,2950|true|false|false|C0040822|Tremor|tremor
Finding|Pathologic Function|SIMPLE_SEGMENT|2954,2968|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|SIMPLE_SEGMENT|2963,2968|true|false|false|||drift
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2971,2974|true|false|false|C0008628;C1511760;C4524186|Chromosome Deletion;Deletion Mutation;Double-Expressor Lymphoma|Del
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2971,2974|true|false|false|C0008628;C1511760;C4524186|Chromosome Deletion;Deletion Mutation;Double-Expressor Lymphoma|Del
Finding|Gene or Genome|SIMPLE_SEGMENT|2975,2978|true|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|SIMPLE_SEGMENT|2975,2978|true|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Drug|Organic Chemical|SIMPLE_SEGMENT|2975,2981|true|false|false|C0053809|Bistris|Tri Bi
Event|Event|SIMPLE_SEGMENT|3076,3085|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|3076,3085|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3076,3085|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3076,3085|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|3087,3093|false|false|false|||Intact
Finding|Finding|SIMPLE_SEGMENT|3087,3093|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3097,3102|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3097,3102|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|3097,3102|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|3097,3102|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|3097,3102|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|3097,3102|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3097,3102|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3097,3102|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|3097,3108|false|false|false|C0423553|Light touch|light touch
Event|Event|SIMPLE_SEGMENT|3103,3108|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|3103,3108|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3103,3108|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3103,3108|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|3110,3118|false|false|false|||pinprick
Event|Event|SIMPLE_SEGMENT|3124,3138|false|false|false|||proprioception
Finding|Mental Process|SIMPLE_SEGMENT|3124,3138|false|false|false|C0033499|Proprioception|proprioception
Event|Event|SIMPLE_SEGMENT|3153,3161|false|false|false|||Reflexes
Finding|Finding|SIMPLE_SEGMENT|3153,3161|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3153,3161|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3153,3161|false|false|false|C0436145|Examination of reflexes|Reflexes
Finding|Conceptual Entity|SIMPLE_SEGMENT|3171,3180|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3171,3180|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3195,3199|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|SIMPLE_SEGMENT|3200,3209|false|false|false|||downgoing
Event|Event|SIMPLE_SEGMENT|3225,3237|false|false|false|||Coordination
Finding|Functional Concept|SIMPLE_SEGMENT|3225,3237|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|3225,3237|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|3225,3237|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3239,3245|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3251,3257|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Event|Event|SIMPLE_SEGMENT|3258,3264|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3266,3270|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3274,3278|false|false|false|C0230444|Shin|shin
Event|Event|SIMPLE_SEGMENT|3279,3285|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|3294,3298|false|false|false|||RAMs
Event|Event|SIMPLE_SEGMENT|3299,3305|false|false|false|||normal
Finding|Finding|SIMPLE_SEGMENT|3310,3314|false|false|false|C0016928|Gait|Gait
Finding|Finding|SIMPLE_SEGMENT|3316,3322|false|false|false|C1837463|Narrow face|Narrow
Finding|Finding|SIMPLE_SEGMENT|3338,3342|true|false|false|C1299581|Able (qualifier value)|Able
Event|Event|SIMPLE_SEGMENT|3353,3357|true|false|false|||walk
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3353,3357|true|false|false|C0080331|Walking (function)|walk
Event|Event|SIMPLE_SEGMENT|3366,3376|true|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|3366,3376|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3378,3385|true|false|false|C0015458|Facial Hemiatrophy|Romberg
Event|Event|SIMPLE_SEGMENT|3378,3385|true|false|false|||Romberg
Event|Event|SIMPLE_SEGMENT|3387,3395|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|3387,3395|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|3387,3395|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3387,3395|false|false|false|C5237010|Expression Negative|Negative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3430,3435|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3430,3435|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3430,3435|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3436,3439|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3444,3447|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3444,3447|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3444,3447|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3453,3456|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3453,3456|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3453,3456|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3453,3456|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3463,3466|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3463,3466|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3473,3476|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3473,3476|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3473,3476|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3473,3476|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3473,3476|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3480,3483|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3480,3483|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3480,3483|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3480,3483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3480,3483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3480,3483|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3490,3494|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3509,3512|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3529,3534|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3529,3534|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3529,3534|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|3550,3555|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3550,3555|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3550,3555|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3560,3563|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3560,3563|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3560,3563|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3590,3595|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3590,3595|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3590,3595|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3600,3603|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3600,3603|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3600,3603|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3625,3630|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3625,3630|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3625,3630|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3625,3638|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3625,3638|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3625,3638|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3631,3638|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3631,3638|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3631,3638|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3631,3638|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3631,3638|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3631,3638|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3682,3686|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3682,3686|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3682,3686|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3711,3716|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3711,3716|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3711,3716|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3717,3720|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3717,3720|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3717,3720|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3717,3720|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3717,3720|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3717,3720|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3717,3720|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3717,3720|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3724,3727|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3724,3727|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3724,3727|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3724,3727|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3724,3727|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3724,3727|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3724,3727|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3734,3737|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|3734,3737|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|3734,3737|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|3734,3737|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3734,3737|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3742,3749|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|3742,3749|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3778,3783|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3778,3783|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3778,3783|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3784,3789|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3784,3789|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3784,3789|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3784,3789|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3824,3829|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3824,3829|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3824,3829|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3842,3849|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3842,3849|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3842,3849|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|3842,3849|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|3842,3849|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|3842,3849|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3842,3849|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3867,3874|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3867,3874|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3867,3874|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3867,3874|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3867,3874|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3867,3874|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3867,3874|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3867,3874|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3907,3912|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3907,3912|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3907,3912|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3914,3919|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3914,3919|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|SIMPLE_SEGMENT|3914,3919|false|false|false|||HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3914,3919|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3936,3941|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3936,3941|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3936,3941|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3942,3945|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|3942,3945|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|3942,3945|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3942,3945|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|3942,3945|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|3942,3945|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|3946,3949|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3946,3949|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3950,3957|false|false|false|C0161679|Toxic effect of ethyl alcohol|Ethanol
Drug|Organic Chemical|SIMPLE_SEGMENT|3950,3957|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3950,3957|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Event|Event|SIMPLE_SEGMENT|3950,3957|false|false|false|||Ethanol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3950,3957|false|false|false|C0202304|Ethanol measurement|Ethanol
Event|Event|SIMPLE_SEGMENT|3958,3961|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3958,3961|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3970,3973|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3970,3973|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3983,3986|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3983,3986|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3995,3998|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3995,3998|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|4007,4010|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4007,4010|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|4012,4021|false|false|false|||Radiology
Finding|Finding|SIMPLE_SEGMENT|4012,4021|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Idea or Concept|SIMPLE_SEGMENT|4012,4021|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Intellectual Product|SIMPLE_SEGMENT|4012,4021|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4012,4021|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|Radiology
Finding|Intellectual Product|SIMPLE_SEGMENT|4012,4028|false|false|false|C1299496|Radiology report|Radiology Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4022,4028|false|false|false|C4255046||Report
Event|Event|SIMPLE_SEGMENT|4022,4028|false|false|false|||Report
Finding|Intellectual Product|SIMPLE_SEGMENT|4022,4028|false|false|false|C0684224|Report (document)|Report
Procedure|Health Care Activity|SIMPLE_SEGMENT|4022,4028|false|false|false|C0700287|Reporting|Report
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4029,4032|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|4029,4032|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4029,4032|false|false|false|C1609165|tocilizumab|MRA
Event|Event|SIMPLE_SEGMENT|4029,4032|false|false|false|||MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4029,4032|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4029,4032|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4033,4038|false|false|false|C0006104;C4266577|Brain;Head>Brain|BRAIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4033,4038|false|false|false|C0006111|Brain Diseases|BRAIN
Event|Event|SIMPLE_SEGMENT|4033,4038|false|false|false|||BRAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4043,4051|false|true|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|4052,4057|false|false|false|||Study
Finding|Intellectual Product|SIMPLE_SEGMENT|4052,4057|false|true|false|C1705923|Study Object|Study
Procedure|Research Activity|SIMPLE_SEGMENT|4052,4057|false|true|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|Study
Finding|Intellectual Product|SIMPLE_SEGMENT|4086,4091|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4092,4104|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|4092,4104|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4105,4116|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4105,4116|true|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|4105,4116|true|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4145,4153|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4145,4153|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4145,4156|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|4165,4170|true|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|4165,4170|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Functional Concept|SIMPLE_SEGMENT|4183,4191|false|false|false|C0475224|Ischemic|ischemic
Event|Event|SIMPLE_SEGMENT|4192,4197|false|true|false|C0441471|Event|event
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4210,4217|true|false|false|C0037303|Bone structure of cranium|cranial
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4222,4230|true|false|false|C0027530|Neck|cervical
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4231,4234|true|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|4231,4234|true|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4231,4234|true|false|false|C1609165|tocilizumab|MRA
Event|Event|SIMPLE_SEGMENT|4231,4234|true|false|false|||MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4231,4234|true|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4231,4234|true|false|false|C0243032|Magnetic Resonance Angiography|MRA
Finding|Idea or Concept|SIMPLE_SEGMENT|4244,4255|true|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|4263,4275|true|false|false|||irregularity
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4280,4284|true|false|false|C0806140|Flow|flow
Event|Event|SIMPLE_SEGMENT|4294,4302|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|4294,4302|false|false|false|C1261287|Stenosis|stenosis
Finding|Intellectual Product|SIMPLE_SEGMENT|4308,4313|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4314,4322|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4314,4329|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4314,4329|false|false|false|C0489547|Hospital course|Hospital Course
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4370,4380|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|4370,4380|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|4370,4380|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|4370,4380|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4382,4386|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|4382,4386|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4392,4401|false|false|false|C0149931|Migraine Disorders|migraines
Event|Event|SIMPLE_SEGMENT|4392,4401|false|false|false|||migraines
Event|Event|SIMPLE_SEGMENT|4403,4413|false|false|false|||presenting
Event|Event|SIMPLE_SEGMENT|4422,4429|false|false|false|||episode
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4433,4439|false|false|false|C0015450|Face|facial
Finding|Sign or Symptom|SIMPLE_SEGMENT|4433,4448|false|false|false|C0239511|Numbness of face|facial numbness
Event|Event|SIMPLE_SEGMENT|4440,4448|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|4440,4448|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4440,4448|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4454,4460|false|false|false|C0015450|Face|Facial
Finding|Sign or Symptom|SIMPLE_SEGMENT|4454,4469|false|false|false|C0239511|Numbness of face|Facial numbness
Event|Event|SIMPLE_SEGMENT|4461,4469|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|4461,4469|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4461,4469|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|4480,4487|false|false|false|||episode
Event|Event|SIMPLE_SEGMENT|4488,4497|false|false|false|||preceeded
Event|Event|SIMPLE_SEGMENT|4500,4508|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|4500,4508|false|false|false|C0018681|Headache|headache
Finding|Finding|SIMPLE_SEGMENT|4519,4525|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4519,4525|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4535,4543|false|false|false|C0149931|Migraine Disorders|migraine
Event|Event|SIMPLE_SEGMENT|4544,4554|false|false|false|||equivalent
Event|Event|SIMPLE_SEGMENT|4564,4571|false|false|false|||episode
Event|Event|SIMPLE_SEGMENT|4587,4590|false|false|false|||due
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4596,4599|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|SIMPLE_SEGMENT|4596,4599|false|false|false|||TIA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4607,4615|false|false|false|C0039729|Thalamic structure|thalamus
Finding|Body Substance|SIMPLE_SEGMENT|4622,4629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4622,4629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4622,4629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|4634,4636|false|false|false|||an
Event|Event|SIMPLE_SEGMENT|4638,4641|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|4638,4641|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4638,4641|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|4638,4641|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|4649,4655|true|false|false|||showed
Event|Event|SIMPLE_SEGMENT|4659,4664|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|4659,4664|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|4659,4664|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|4668,4676|true|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|4668,4676|true|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4668,4676|true|false|false|C4321499|Ischemia Procedure|ischemia
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4689,4700|true|false|false|C3714653|Vasculature|vasculature
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4710,4718|false|false|false|C0149931|Migraine Disorders|migraine
Event|Event|SIMPLE_SEGMENT|4710,4718|false|false|false|||migraine
Event|Event|SIMPLE_SEGMENT|4719,4729|false|false|false|||equivalent
Finding|Finding|SIMPLE_SEGMENT|4732,4736|false|false|false|C4281574|Much|much
Finding|Finding|SIMPLE_SEGMENT|4742,4748|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4742,4748|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4749,4758|false|true|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|4749,4758|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|4749,4758|false|true|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4749,4758|false|true|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4749,4758|false|true|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4796,4799|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|SIMPLE_SEGMENT|4796,4799|false|false|false|||TIA
Event|Event|SIMPLE_SEGMENT|4814,4821|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|4834,4841|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4834,4841|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|4834,4841|false|false|false|||aspirin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4853,4859|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|4853,4859|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|4853,4859|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|SIMPLE_SEGMENT|4860,4871|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4860,4871|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|4874,4878|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|4874,4878|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4874,4878|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|4882,4891|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4882,4891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4882,4891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4882,4891|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4882,4891|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|4897,4904|false|false|false|||notable
Finding|Intellectual Product|SIMPLE_SEGMENT|4909,4913|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Conceptual Entity|SIMPLE_SEGMENT|4914,4923|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|4914,4923|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|4924,4937|false|false|false|||hyperreflexia
Finding|Finding|SIMPLE_SEGMENT|4924,4937|false|false|false|C0151889|Hyperreflexia|hyperreflexia
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4945,4950|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4945,4950|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4952,4963|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4986,5003|true|false|false|C0027853|Neurologic Examination|neurological exam
Event|Event|SIMPLE_SEGMENT|4999,5003|true|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|4999,5003|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4999,5003|true|false|false|C0582103|Medical Examination|exam
Finding|Finding|SIMPLE_SEGMENT|5023,5039|true|false|false|C0748618|Sensory deficit|sensory deficits
Event|Event|SIMPLE_SEGMENT|5031,5039|true|false|false|||deficits
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5043,5054|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5043,5054|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5043,5054|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5043,5054|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|5043,5067|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|5058,5067|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5058,5067|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|5069,5075|false|false|false|C0939400|Nexium|NEXIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5069,5075|false|false|false|C0939400|Nexium|NEXIUM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5085,5092|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5085,5092|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5085,5092|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|5096,5104|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5099,5104|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5099,5104|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|5105,5109|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5105,5115|false|false|false|C3537736|Once A Day|once a day
Event|Event|SIMPLE_SEGMENT|5112,5115|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|5112,5115|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5112,5115|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|5116,5122|false|false|false|C0162373|Prozac|PROZAC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5116,5122|false|false|false|C0162373|Prozac|PROZAC
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5132,5139|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5132,5139|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5132,5139|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|5143,5151|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5146,5151|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5146,5151|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|5152,5156|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5152,5162|false|false|false|C3537736|Once A Day|once a day
Event|Event|SIMPLE_SEGMENT|5159,5162|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|5159,5162|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5159,5162|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5166,5175|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5166,5175|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5166,5175|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5166,5175|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5166,5175|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5166,5187|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5176,5187|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5176,5187|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5176,5187|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5176,5187|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|5192,5204|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5192,5204|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5211,5217|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5211,5217|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5219,5226|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5219,5234|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5227,5234|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5227,5234|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5227,5234|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5227,5234|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|5242,5245|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5256,5262|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5256,5262|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5264,5271|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5264,5279|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5272,5279|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5272,5279|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5272,5279|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5272,5279|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|5318,5328|false|false|false|C0016365|fluoxetine|Fluoxetine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5318,5328|false|false|false|C0016365|fluoxetine|Fluoxetine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5335,5342|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5335,5342|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5335,5342|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5356,5363|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5356,5363|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5356,5363|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|SIMPLE_SEGMENT|5388,5395|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5388,5395|false|false|false|C0004057|aspirin|Aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5402,5408|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5402,5408|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5410,5417|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5410,5425|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5418,5425|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5418,5425|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5418,5425|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5418,5425|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|5433,5436|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5447,5453|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5447,5453|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5455,5462|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5455,5470|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5463,5470|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5463,5470|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5463,5470|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5463,5470|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|5501,5510|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5501,5510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5501,5510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5501,5510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5501,5510|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5501,5522|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|5501,5522|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5511,5522|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|5511,5522|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|5511,5522|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|5524,5528|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|5524,5528|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|5524,5528|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5524,5528|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|5531,5540|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5531,5540|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5531,5540|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5531,5540|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5531,5540|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5531,5550|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5541,5550|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|5541,5550|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|5541,5550|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|5541,5550|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5541,5550|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5552,5560|false|false|false|C0149931|Migraine Disorders|Migraine
Event|Event|SIMPLE_SEGMENT|5552,5560|false|false|false|||Migraine
Event|Event|SIMPLE_SEGMENT|5564,5573|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5564,5573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5564,5573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5564,5573|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5564,5573|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5574,5583|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5574,5583|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|5574,5583|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|5574,5583|false|false|false|C1705253|Logical Condition|Condition
Finding|Intellectual Product|SIMPLE_SEGMENT|5585,5589|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Conceptual Entity|SIMPLE_SEGMENT|5590,5599|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|5590,5599|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|5600,5613|false|false|false|||hyperreflexia
Finding|Finding|SIMPLE_SEGMENT|5600,5613|false|false|false|C0151889|Hyperreflexia|hyperreflexia
Finding|Finding|SIMPLE_SEGMENT|5600,5638|false|false|false|C4015304|Hyperreflexia in the lower extremities|hyperreflexia in the lower extremities
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5621,5626|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5621,5626|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5621,5638|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5627,5638|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5658,5675|false|false|false|C0027853|Neurologic Examination|neurological exam
Event|Event|SIMPLE_SEGMENT|5671,5675|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|5671,5675|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5671,5675|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|5680,5689|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5680,5689|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5680,5689|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5680,5689|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5680,5689|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5680,5702|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5680,5702|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|5680,5702|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5690,5702|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|5690,5702|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5690,5702|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|5713,5721|false|false|false|||admitted
Finding|Functional Concept|SIMPLE_SEGMENT|5726,5730|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5737,5743|false|false|false|C0015450|Face|facial
Finding|Sign or Symptom|SIMPLE_SEGMENT|5737,5752|false|false|false|C0239511|Numbness of face|facial numbness
Event|Event|SIMPLE_SEGMENT|5744,5752|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|5744,5752|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|5744,5752|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|5767,5770|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|5767,5770|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5767,5770|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|5767,5770|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|5777,5783|true|false|false|||showed
Event|Event|SIMPLE_SEGMENT|5787,5792|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|5787,5792|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|5787,5792|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|5796,5804|true|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|5796,5804|true|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5796,5804|true|false|false|C4321499|Ischemia Procedure|ischemia
Event|Event|SIMPLE_SEGMENT|5813,5822|false|false|false|||suspected
Drug|Organic Chemical|SIMPLE_SEGMENT|5838,5845|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|5838,5845|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|5838,5845|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|5838,5845|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5849,5857|false|false|false|C0149931|Migraine Disorders|migraine
Event|Event|SIMPLE_SEGMENT|5849,5857|false|false|false|||migraine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5849,5867|false|false|false|C0149931|Migraine Disorders|migraine headaches
Event|Event|SIMPLE_SEGMENT|5858,5867|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|5858,5867|false|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|5876,5885|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|5896,5901|false|false|false|||start
Event|Event|SIMPLE_SEGMENT|5916,5920|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|5924,5931|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5924,5931|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|5924,5931|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|5941,5947|false|false|false|||notice
Finding|Finding|SIMPLE_SEGMENT|5948,5951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5948,5951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|5952,5960|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|5952,5960|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|5952,5960|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|5962,5970|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|5962,5970|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|5982,5991|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|5982,5991|false|false|false|C0018681|Headache|headaches
Finding|Finding|SIMPLE_SEGMENT|6003,6006|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6003,6006|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|6018,6026|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6018,6026|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6018,6026|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6035,6041|false|false|false|||return
Event|Event|SIMPLE_SEGMENT|6073,6083|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|6073,6083|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6073,6083|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6087,6095|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6096,6108|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6096,6108|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6096,6108|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

