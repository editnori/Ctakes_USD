 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Chief|210,215
Complaint|216,225
:|225,226
<EOL>|226,227
chest|227,232
pain|233,237
<EOL>|237,238
<EOL>|239,240
Major|240,245
Surgical|246,254
or|255,257
Invasive|258,266
Procedure|267,276
:|276,277
<EOL>|277,278
cardiac|278,285
catheterization|286,301
<EOL>|301,302
<EOL>|302,303
<EOL>|304,305
History|305,312
of|313,315
Present|316,323
Illness|324,331
:|331,332
<EOL>|332,333
_|333,334
_|334,335
_|335,336
w|337,338
/|338,339
PMH|340,343
of|344,346
CAD|347,350
s|351,352
/|352,353
p|353,354
PCI|355,358
x3|359,361
,|361,362
s|363,364
/|364,365
p|365,366
off|367,370
-|370,371
pump|371,375
CABG|376,380
x3|381,383
_|384,385
_|385,386
_|386,387
<EOL>|388,389
(|389,390
_|390,391
_|391,392
_|392,393
-|393,394
-|394,395
>|395,396
LAD|396,399
,|399,400
SVG|401,404
-|405,406
-|406,407
>|407,408
diag|408,412
,|412,413
OM|414,416
)|416,417
,|417,418
type|419,423
2|424,425
DM|426,428
on|429,431
insulin|432,439
,|439,440
HTN|441,444
,|444,445
<EOL>|446,447
hyperlipidemia|447,461
presents|462,470
with|471,475
a|476,477
3|478,479
day|480,483
history|484,491
of|492,494
_|495,496
_|496,497
_|497,498
sharp|499,504
,|504,505
<EOL>|506,507
left|507,511
-|511,512
sided|512,517
chest|518,523
pain|524,528
and|529,532
SOB|533,536
.|536,537
She|538,541
describes|542,551
the|552,555
chest|556,561
pain|562,566
as|567,569
<EOL>|570,571
"|571,572
pinching|572,580
all|581,584
the|585,588
way|589,592
down|593,597
to|598,600
the|601,604
bone|605,609
.|609,610
"|610,611
She|612,615
endorses|616,624
_|625,626
_|626,627
_|627,628
<EOL>|629,630
episodes|630,638
of|639,641
pain|642,646
/|646,647
day|647,650
,|650,651
always|652,658
at|659,661
rest|662,666
.|666,667
The|668,671
episodes|672,680
of|681,683
pain|684,688
last|689,693
<EOL>|694,695
approximately|695,708
5|709,710
minutes|711,718
and|719,722
are|723,726
relieved|727,735
by|736,738
nitroglycerin|739,752
.|752,753
Her|754,757
<EOL>|758,759
pain|759,763
is|764,766
not|767,770
worsened|771,779
by|780,782
exertion|783,791
or|792,794
eating|795,801
.|801,802
She|803,806
described|807,816
her|817,820
<EOL>|821,822
symptoms|822,830
to|831,833
her|834,837
PCP|838,841
over|842,846
the|847,850
phone|851,856
,|856,857
who|858,861
told|862,866
her|867,870
to|871,873
come|874,878
to|879,881
the|882,885
<EOL>|886,887
ED|887,889
.|889,890
She|891,894
says|895,899
they|900,904
feel|905,909
similar|910,917
to|918,920
her|921,924
MI|925,927
in|928,930
the|931,934
past|935,939
.|939,940
She|941,944
also|945,949
<EOL>|950,951
endorsed|951,959
vomiting|960,968
last|969,973
night|974,979
.|979,980
She|981,984
denies|985,991
any|992,995
diaphoresis|996,1007
.|1007,1008
She|1009,1012
<EOL>|1013,1014
also|1014,1018
endorses|1019,1027
a|1028,1029
cough|1030,1035
.|1035,1036
<EOL>|1038,1039
The|1039,1042
patient|1043,1050
has|1051,1054
developed|1055,1064
increased|1065,1074
shortness|1075,1084
of|1085,1087
breath|1088,1094
over|1095,1099
the|1100,1103
<EOL>|1104,1105
past|1105,1109
few|1110,1113
days|1114,1118
.|1118,1119
She|1120,1123
has|1124,1127
experienced|1128,1139
orthopnea|1140,1149
for|1150,1153
the|1154,1157
past|1158,1162
few|1163,1166
<EOL>|1167,1168
years|1168,1173
,|1173,1174
but|1175,1178
denies|1179,1185
PND|1186,1189
and|1190,1193
lower|1194,1199
extremity|1200,1209
edema|1210,1215
.|1215,1216
On|1217,1219
exam|1220,1224
in|1225,1227
the|1228,1231
<EOL>|1232,1233
ED|1233,1235
she|1236,1239
was|1240,1243
tachycardic|1244,1255
,|1255,1256
in|1257,1259
a|1260,1261
regular|1262,1269
rhythm|1270,1276
.|1276,1277
Lungs|1278,1283
were|1284,1288
CTAB|1289,1293
.|1293,1294
<EOL>|1295,1296
She|1296,1299
had|1300,1303
trace|1304,1309
edema|1310,1315
in|1316,1318
her|1319,1322
left|1323,1327
lower|1328,1333
extremity|1334,1343
,|1343,1344
none|1345,1349
in|1350,1352
her|1353,1356
<EOL>|1357,1358
right|1358,1363
leg|1364,1367
.|1367,1368
<EOL>|1370,1371
<EOL>|1372,1373
In|1373,1375
the|1376,1379
ED|1380,1382
,|1382,1383
initial|1384,1391
vitals|1392,1398
were|1399,1403
96.8|1404,1408
111|1409,1412
177|1413,1416
/|1416,1417
86|1417,1419
18|1420,1422
97|1423,1425
%|1425,1426
.|1426,1427
Labs|1428,1432
and|1433,1436
<EOL>|1437,1438
imaging|1438,1445
significant|1446,1457
for|1458,1461
a|1462,1463
CXR|1464,1467
with|1468,1472
new|1473,1476
moderate|1477,1485
left|1486,1490
pleural|1491,1498
<EOL>|1499,1500
effusion|1500,1508
with|1509,1513
adjacent|1514,1522
atelectasis|1523,1534
in|1535,1537
the|1538,1541
left|1542,1546
lung|1547,1551
base|1552,1556
,|1556,1557
CBC|1558,1561
<EOL>|1562,1563
within|1563,1569
normal|1570,1576
limits|1577,1583
,|1583,1584
electrolytes|1585,1597
within|1598,1604
normal|1605,1611
limits|1612,1618
,|1618,1619
Cr|1620,1622
.|1622,1623
<EOL>|1624,1625
1.2|1625,1628
,|1628,1629
troponin|1630,1638
0.08|1639,1643
and|1644,1647
D|1648,1649
-|1649,1650
dimer|1650,1655
2350|1656,1660
.|1660,1661
A|1662,1663
CT|1664,1666
of|1667,1669
the|1670,1673
chest|1674,1679
was|1680,1683
<EOL>|1684,1685
performed|1685,1694
,|1694,1695
which|1696,1701
showed|1702,1708
no|1709,1711
CT|1712,1714
evidence|1715,1723
for|1724,1727
pulmonary|1728,1737
embolus|1738,1745
,|1745,1746
<EOL>|1747,1748
but|1748,1751
small|1752,1757
left|1758,1762
pleural|1763,1770
effusion|1771,1779
with|1780,1784
adjacent|1785,1793
atelectasis|1794,1805
.|1805,1806
<EOL>|1808,1809
Patient|1809,1816
given|1817,1822
aspirin|1823,1830
81mg|1831,1835
x|1836,1837
4|1838,1839
,|1839,1840
SL|1841,1843
nitroglycerin|1844,1857
x|1858,1859
1|1860,1861
and|1862,1865
heparin|1866,1873
<EOL>|1874,1875
bolus|1875,1880
.|1880,1881
<EOL>|1883,1884
Vitals|1884,1890
on|1891,1893
transfer|1894,1902
were|1903,1907
99.2|1908,1912
112|1913,1916
162|1917,1920
/|1920,1921
82|1921,1923
22|1924,1926
98|1927,1929
%|1929,1930
RA|1931,1933
<EOL>|1935,1936
On|1936,1938
arrival|1939,1946
to|1947,1949
the|1950,1953
floor|1954,1959
,|1959,1960
patient|1961,1968
is|1969,1971
AAOx3|1972,1977
,|1977,1978
and|1979,1982
comfortable|1983,1994
.|1994,1995
<EOL>|1997,1998
<EOL>|1999,2000
REVIEW|2000,2006
OF|2007,2009
SYSTEMS|2010,2017
<EOL>|2019,2020
On|2020,2022
review|2023,2029
of|2030,2032
systems|2033,2040
,|2040,2041
she|2042,2045
denies|2046,2052
any|2053,2056
prior|2057,2062
history|2063,2070
of|2071,2073
stroke|2074,2080
,|2080,2081
<EOL>|2082,2083
TIA|2083,2086
,|2086,2087
deep|2088,2092
venous|2093,2099
thrombosis|2100,2110
,|2110,2111
pulmonary|2112,2121
embolism|2122,2130
,|2130,2131
bleeding|2132,2140
at|2141,2143
the|2144,2147
<EOL>|2148,2149
time|2149,2153
of|2154,2156
surgery|2157,2164
,|2164,2165
myalgias|2166,2174
,|2174,2175
joint|2176,2181
pains|2182,2187
,|2187,2188
cough|2189,2194
,|2194,2195
hemoptysis|2196,2206
,|2206,2207
black|2208,2213
<EOL>|2214,2215
stools|2215,2221
or|2222,2224
red|2225,2228
stools|2229,2235
.|2235,2236
She|2237,2240
denies|2241,2247
recent|2248,2254
fevers|2255,2261
,|2261,2262
chills|2263,2269
or|2270,2272
<EOL>|2273,2274
rigors|2274,2280
.|2280,2281
She|2282,2285
denies|2286,2292
exertional|2293,2303
buttock|2304,2311
or|2312,2314
calf|2315,2319
pain|2320,2324
.|2324,2325
All|2326,2329
of|2330,2332
the|2333,2336
<EOL>|2337,2338
other|2338,2343
review|2344,2350
of|2351,2353
systems|2354,2361
were|2362,2366
negative|2367,2375
.|2375,2376
<EOL>|2378,2379
<EOL>|2379,2380
<EOL>|2381,2382
Past|2382,2386
Medical|2387,2394
History|2395,2402
:|2402,2403
<EOL>|2403,2404
1.|2404,2406
CARDIAC|2407,2414
RISK|2415,2419
FACTORS|2420,2427
:|2427,2428
(|2429,2430
-|2430,2431
)|2431,2432
Diabetes|2432,2440
,|2440,2441
(|2442,2443
+|2443,2444
)|2444,2445
Dyslipidemia|2445,2457
,|2457,2458
(|2459,2460
+|2460,2461
)|2461,2462
HTN|2462,2465
<EOL>|2467,2468
2.|2468,2470
CARDIAC|2471,2478
HISTORY|2479,2486
:|2486,2487
<EOL>|2489,2490
-|2490,2491
Coronary|2491,2499
artery|2500,2506
disease|2507,2514
<EOL>|2516,2517
-|2517,2518
Diastolic|2518,2527
congestive|2528,2538
heart|2539,2544
failure|2545,2552
<EOL>|2554,2555
-|2555,2556
CABG|2556,2560
:|2560,2561
CABG|2562,2566
x|2567,2568
3|2569,2570
(|2571,2572
Off|2572,2575
pump|2576,2580
coronary|2581,2589
artery|2590,2596
bypass|2597,2603
graft|2604,2609
x3|2610,2612
,|2612,2613
left|2614,2618
<EOL>|2620,2621
<EOL>|2621,2622
internal|2622,2630
mammary|2631,2638
artery|2639,2645
to|2646,2648
left|2649,2653
anterior|2654,2662
descending|2663,2673
artery|2674,2680
and|2681,2684
<EOL>|2686,2687
saphenous|2687,2696
vein|2697,2701
grafts|2702,2708
to|2709,2711
diagonal|2712,2720
,|2720,2721
and|2722,2725
obtuse|2726,2732
marginal|2733,2741
arteries|2742,2750
)|2750,2751
<EOL>|2752,2753
<EOL>|2754,2755
-|2755,2756
PERCUTANEOUS|2756,2768
CORONARY|2769,2777
INTERVENTIONS|2778,2791
:|2791,2792
BMS|2793,2796
to|2797,2799
proximal|2800,2808
LAD|2809,2812
<EOL>|2814,2815
_|2815,2816
_|2816,2817
_|2817,2818
,|2818,2819
DES|2820,2823
to|2824,2826
mid|2827,2830
LAD|2831,2834
_|2835,2836
_|2836,2837
_|2837,2838
,|2838,2839
DES|2840,2843
to|2844,2846
edge|2847,2851
ISR|2852,2855
of|2856,2858
mid|2859,2862
LAD|2863,2866
DES|2867,2870
and|2871,2874
<EOL>|2876,2877
stenosis|2877,2885
distal|2886,2892
to|2893,2895
stent|2896,2901
_|2902,2903
_|2903,2904
_|2904,2905
,|2905,2906
DES|2907,2910
to|2911,2913
OM1|2914,2917
,|2917,2918
_|2919,2920
_|2920,2921
_|2921,2922
<EOL>|2924,2925
-|2925,2926
PACING|2926,2932
/|2932,2933
ICD|2933,2936
:|2936,2937
none|2937,2941
<EOL>|2943,2944
Morbid|2944,2950
obesity|2951,2958
.|2958,2959
<EOL>|2961,2962
COPD|2962,2966
<EOL>|2968,2969
GERD|2969,2973
<EOL>|2975,2976
Right|2976,2981
rotator|2982,2989
cuff|2990,2994
injury|2995,3001
/|3001,3002
bursitis|3002,3010
<EOL>|3012,3013
Migraines|3013,3022
<EOL>|3024,3025
Depression|3025,3035
<EOL>|3037,3038
DJD|3038,3041
<EOL>|3043,3044
Hemorrhoids|3044,3055
<EOL>|3057,3058
Rosacea|3058,3065
<EOL>|3067,3068
<EOL>|3068,3069
<EOL>|3070,3071
Social|3071,3077
History|3078,3085
:|3085,3086
<EOL>|3086,3087
_|3087,3088
_|3088,3089
_|3089,3090
<EOL>|3090,3091
Family|3091,3097
History|3098,3105
:|3105,3106
<EOL>|3106,3107
She|3107,3110
was|3111,3114
a|3115,3116
ward|3117,3121
of|3122,3124
the|3125,3128
_|3129,3130
_|3130,3131
_|3131,3132
and|3133,3136
does|3137,3141
not|3142,3145
know|3146,3150
her|3151,3154
family|3155,3161
.|3161,3162
<EOL>|3164,3165
<EOL>|3165,3166
<EOL>|3167,3168
Physical|3168,3176
Exam|3177,3181
:|3181,3182
<EOL>|3182,3183
Admission|3183,3192
:|3192,3193
<EOL>|3193,3194
VS|3194,3196
-|3196,3197
T|3198,3199
99.4|3200,3204
BP|3205,3207
157|3208,3211
/|3211,3212
88|3212,3214
HR|3215,3217
118|3218,3221
RR|3222,3224
24|3225,3227
96|3228,3230
%|3230,3231
RA|3232,3234
<EOL>|3236,3237
GENERAL|3237,3244
-|3244,3245
WDWN|3246,3250
F|3251,3252
in|3253,3255
NAD|3256,3259
.|3259,3260
Oriented|3261,3269
x3|3270,3272
.|3272,3273
Mood|3274,3278
,|3278,3279
affect|3280,3286
appropriate|3287,3298
.|3298,3299
<EOL>|3301,3302
HEENT|3302,3307
-|3307,3308
NCAT|3309,3313
.|3313,3314
Sclera|3315,3321
anicteric|3322,3331
.|3331,3332
PERRL|3333,3338
,|3338,3339
EOMI|3340,3344
.|3344,3345
Conjunctiva|3346,3357
were|3358,3362
<EOL>|3363,3364
pink|3364,3368
,|3368,3369
no|3370,3372
pallor|3373,3379
or|3380,3382
cyanosis|3383,3391
of|3392,3394
the|3395,3398
oral|3399,3403
mucosa|3404,3410
.|3410,3411
No|3412,3414
xanthalesma|3415,3426
.|3426,3427
<EOL>|3429,3430
<EOL>|3430,3431
NECK|3431,3435
-|3435,3436
Supple|3437,3443
without|3444,3451
JVP|3452,3455
<EOL>|3457,3458
CARDIAC|3458,3465
-|3465,3466
PMI|3467,3470
located|3471,3478
in|3479,3481
_|3482,3483
_|3483,3484
_|3484,3485
intercostal|3486,3497
space|3498,3503
,|3503,3504
midclavicular|3505,3518
<EOL>|3519,3520
line|3520,3524
.|3524,3525
RRR|3526,3529
Nl|3530,3532
S1|3533,3535
/|3535,3536
S2|3536,3538
.|3538,3539
Midline|3540,3547
scar|3548,3552
from|3553,3557
recent|3558,3564
surgery|3565,3572
C|3573,3574
/|3574,3575
D|3575,3576
/|3576,3577
I|3577,3578
<EOL>|3580,3581
LUNGS|3581,3586
-|3587,3588
No|3589,3591
chest|3592,3597
wall|3598,3602
deformities|3603,3614
,|3614,3615
scoliosis|3616,3625
or|3626,3628
kyphosis|3629,3637
.|3637,3638
Resp|3639,3643
<EOL>|3644,3645
were|3645,3649
unlabored|3650,3659
,|3659,3660
no|3661,3663
accessory|3664,3673
muscle|3674,3680
use|3681,3684
.|3684,3685
CTAB|3686,3690
,|3690,3691
no|3692,3694
crackles|3695,3703
,|3703,3704
<EOL>|3705,3706
wheezes|3706,3713
or|3714,3716
rhonchi|3717,3724
.|3724,3725
<EOL>|3727,3728
ABDOMEN|3728,3735
-|3735,3736
Soft|3737,3741
,|3741,3742
NTND|3743,3747
.|3747,3748
No|3749,3751
HSM|3752,3755
or|3756,3758
tenderness|3759,3769
.|3769,3770
<EOL>|3772,3773
EXTREMITIES|3773,3784
-|3784,3785
No|3786,3788
c|3789,3790
/|3790,3791
c|3791,3792
/|3792,3793
e|3793,3794
.|3794,3795
<EOL>|3796,3797
<EOL>|3797,3798
Discharge|3798,3807
:|3807,3808
<EOL>|3808,3809
Vitals|3809,3815
:|3815,3816
T|3817,3818
:|3818,3819
98.4|3819,3823
BP|3824,3826
:|3826,3827
151|3827,3830
/|3830,3831
90|3831,3833
P|3834,3835
:|3835,3836
86|3836,3838
R|3839,3840
:|3840,3841
20|3841,3843
O2|3844,3846
:|3846,3847
97|3847,3849
RA|3850,3852
<EOL>|3854,3855
I|3855,3856
/|3856,3857
O|3857,3858
:|3858,3859
Intake|3860,3866
:|3866,3867
840|3868,3871
mL|3872,3874
;|3874,3875
Output|3876,3882
:|3882,3883
Voided|3884,3890
x2|3891,3893
(|3894,3895
not|3895,3898
recorded|3899,3907
)|3907,3908
<EOL>|3909,3910
GENERAL|3910,3917
-|3918,3919
Alert|3920,3925
,|3925,3926
interactive|3927,3938
,|3938,3939
well|3940,3944
-|3944,3945
appearing|3945,3954
in|3955,3957
NAD|3958,3961
<EOL>|3963,3964
HEENT|3964,3969
-|3970,3971
PERRLA|3972,3978
,|3978,3979
EOMI|3980,3984
,|3984,3985
sclerae|3986,3993
anicteric|3994,4003
,|4003,4004
dry|4005,4008
mucous|4009,4015
membranes|4016,4025
,|4025,4026
<EOL>|4027,4028
OP|4028,4030
clear|4031,4036
,|4036,4037
no|4038,4040
JVP|4041,4044
visualized|4045,4055
<EOL>|4058,4059
HEART|4059,4064
-|4065,4066
RRR|4067,4070
,|4070,4071
nl|4072,4074
S1|4075,4077
-|4077,4078
S2|4078,4080
,|4080,4081
no|4082,4084
MRG|4085,4088
.|4088,4089
Scar|4090,4094
from|4095,4099
recent|4100,4106
surgery|4107,4114
present|4115,4122
<EOL>|4123,4124
at|4124,4126
midline|4127,4134
.|4134,4135
Wound|4136,4141
is|4142,4144
healing|4145,4152
well|4153,4157
,|4157,4158
no|4159,4161
tenderness|4162,4172
along|4173,4178
scar|4179,4183
.|4183,4184
<EOL>|4185,4186
Slight|4186,4192
erythema|4193,4201
at|4202,4204
base|4205,4209
.|4209,4210
A|4211,4212
2|4213,4214
cm|4215,4217
area|4218,4222
of|4223,4225
newer|4226,4231
scar|4232,4236
is|4237,4239
present|4240,4247
<EOL>|4248,4249
from|4249,4253
previous|4254,4262
debridement|4263,4274
as|4275,4277
reported|4278,4286
per|4287,4290
patinent|4291,4299
.|4299,4300
<EOL>|4304,4305
LUNGS|4305,4310
-|4311,4312
Bibasilar|4313,4322
crackles|4323,4331
present|4332,4339
at|4340,4342
bases|4343,4348
.|4348,4349
No|4350,4352
wheezes|4353,4360
or|4361,4363
<EOL>|4364,4365
rhonci|4365,4371
.|4371,4372
Respirations|4373,4385
unlabored|4386,4395
.|4395,4396
<EOL>|4398,4399
ABDOMEN|4399,4406
-|4407,4408
NABS|4409,4413
,|4413,4414
soft|4415,4419
/|4419,4420
NT|4420,4422
/|4422,4423
ND|4423,4425
,|4425,4426
no|4427,4429
masses|4430,4436
or|4437,4439
HSM|4440,4443
<EOL>|4445,4446
EXTREMITIES|4446,4457
-|4458,4459
WWP|4460,4463
,|4463,4464
no|4465,4467
c|4468,4469
/|4469,4470
c|4470,4471
/|4471,4472
e|4472,4473
,|4473,4474
2|4475,4476
+|4476,4477
peripheral|4478,4488
pulses|4489,4495
<EOL>|4497,4498
NEURO|4498,4503
-|4504,4505
awake|4506,4511
,|4511,4512
A|4513,4514
&|4514,4515
Ox3|4515,4518
,|4518,4519
CNs|4520,4523
II|4524,4526
-|4526,4527
XII|4527,4530
grossly|4531,4538
intact|4539,4545
<EOL>|4547,4548
<EOL>|4549,4550
Pertinent|4550,4559
Results|4560,4567
:|4567,4568
<EOL>|4568,4569
Admission|4569,4578
labs|4579,4583
:|4583,4584
<EOL>|4584,4585
_|4585,4586
_|4586,4587
_|4587,4588
03|4589,4591
:|4591,4592
45PM|4592,4596
WBC|4599,4602
-|4602,4603
8.9|4603,4606
RBC|4607,4610
-|4610,4611
3|4611,4612
.|4612,4613
69|4613,4615
*|4615,4616
HGB|4617,4620
-|4620,4621
12.3|4621,4625
HCT|4626,4629
-|4629,4630
34|4630,4632
.|4632,4633
9|4633,4634
*|4634,4635
MCV|4636,4639
-|4639,4640
95|4640,4642
<EOL>|4643,4644
MCH|4644,4647
-|4647,4648
33|4648,4650
.|4650,4651
2|4651,4652
*|4652,4653
MCHC|4654,4658
-|4658,4659
35|4659,4661
.|4661,4662
1|4662,4663
*|4663,4664
RDW|4665,4668
-|4668,4669
13.1|4669,4673
<EOL>|4673,4674
_|4674,4675
_|4675,4676
_|4676,4677
03|4678,4680
:|4680,4681
45PM|4681,4685
NEUTS|4688,4693
-|4693,4694
67.9|4694,4698
_|4699,4700
_|4700,4701
_|4701,4702
MONOS|4703,4708
-|4708,4709
5.5|4709,4712
EOS|4713,4716
-|4716,4717
2.6|4717,4720
<EOL>|4721,4722
BASOS|4722,4727
-|4727,4728
0.9|4728,4731
<EOL>|4731,4732
_|4732,4733
_|4733,4734
_|4734,4735
03|4736,4738
:|4738,4739
45PM|4739,4743
GLUCOSE|4746,4753
-|4753,4754
484|4754,4757
*|4757,4758
UREA|4759,4763
N|4764,4765
-|4765,4766
16|4766,4768
CREAT|4769,4774
-|4774,4775
1|4775,4776
.|4776,4777
2|4777,4778
*|4778,4779
SODIUM|4780,4786
-|4786,4787
135|4787,4790
<EOL>|4791,4792
POTASSIUM|4792,4801
-|4801,4802
3.7|4802,4805
CHLORIDE|4806,4814
-|4814,4815
95|4815,4817
*|4817,4818
TOTAL|4819,4824
CO2|4825,4828
-|4828,4829
26|4829,4831
ANION|4832,4837
GAP|4838,4841
-|4841,4842
18|4842,4844
<EOL>|4844,4845
_|4845,4846
_|4846,4847
_|4847,4848
04|4849,4851
:|4851,4852
25PM|4852,4856
_|4859,4860
_|4860,4861
_|4861,4862
PTT|4863,4866
-|4866,4867
27.8|4867,4871
_|4872,4873
_|4873,4874
_|4874,4875
<EOL>|4875,4876
_|4876,4877
_|4877,4878
_|4878,4879
03|4880,4882
:|4882,4883
45PM|4883,4887
cTropnT|4890,4897
-|4897,4898
0|4898,4899
.|4899,4900
08|4900,4902
*|4902,4903
<EOL>|4903,4904
_|4904,4905
_|4905,4906
_|4906,4907
03|4908,4910
:|4910,4911
45PM|4911,4915
CK|4918,4920
(|4920,4921
CPK|4921,4924
)|4924,4925
-|4925,4926
51|4926,4928
<EOL>|4928,4929
_|4929,4930
_|4930,4931
_|4931,4932
03|4933,4935
:|4935,4936
45PM|4936,4940
D|4943,4944
-|4944,4945
DIMER|4945,4950
-|4950,4951
2350|4951,4955
*|4955,4956
<EOL>|4956,4957
<EOL>|4957,4958
Pertinent|4958,4967
labs|4968,4972
:|4972,4973
<EOL>|4973,4974
_|4974,4975
_|4975,4976
_|4976,4977
03|4978,4980
:|4980,4981
45PM|4981,4985
BLOOD|4986,4991
cTropnT|4992,4999
-|4999,5000
0|5000,5001
.|5001,5002
08|5002,5004
*|5004,5005
<EOL>|5005,5006
_|5006,5007
_|5007,5008
_|5008,5009
12|5010,5012
:|5012,5013
09AM|5013,5017
BLOOD|5018,5023
CK|5024,5026
-|5026,5027
MB|5027,5029
-|5029,5030
3|5030,5031
cTropnT|5032,5039
-|5039,5040
0|5040,5041
.|5041,5042
12|5042,5044
*|5044,5045
<EOL>|5045,5046
_|5046,5047
_|5047,5048
_|5048,5049
07|5050,5052
:|5052,5053
15AM|5053,5057
BLOOD|5058,5063
CK|5064,5066
-|5066,5067
MB|5067,5069
-|5069,5070
3|5070,5071
cTropnT|5072,5079
-|5079,5080
0|5080,5081
.|5081,5082
13|5082,5084
*|5084,5085
<EOL>|5085,5086
<EOL>|5086,5087
Imaging|5087,5094
/|5094,5095
studies|5095,5102
:|5102,5103
<EOL>|5103,5104
EKG|5104,5107
on|5108,5110
admission|5111,5120
-|5120,5121
Sinus|5122,5127
tachycardia|5128,5139
.|5139,5140
Extensive|5141,5150
ST|5151,5153
segment|5154,5161
<EOL>|5162,5163
changes|5163,5170
may|5171,5174
be|5175,5177
due|5178,5181
to|5182,5184
ischemia|5185,5193
.|5193,5194
Compared|5195,5203
to|5204,5206
the|5207,5210
previous|5211,5219
tracing|5220,5227
<EOL>|5228,5229
no|5229,5231
change|5232,5238
.|5238,5239
<EOL>|5241,5242
<EOL>|5242,5243
CXR|5243,5246
_|5247,5248
_|5248,5249
_|5249,5250
-|5250,5251
New|5252,5255
moderate|5256,5264
left|5265,5269
pleural|5270,5277
effusion|5278,5286
with|5287,5291
adjacent|5292,5300
<EOL>|5301,5302
atelectasis|5302,5313
in|5314,5316
the|5317,5320
left|5321,5325
lung|5326,5330
base|5331,5335
.|5335,5336
<EOL>|5337,5338
<EOL>|5340,5341
CTA|5341,5344
Chest|5345,5350
_|5351,5352
_|5352,5353
_|5353,5354
.|5354,5355
No|5357,5359
CT|5360,5362
evidence|5363,5371
for|5372,5375
pulmonary|5376,5385
embolus|5386,5393
.|5393,5394
<EOL>|5395,5396
2.|5396,5398
Small|5400,5405
left|5406,5410
pleural|5411,5418
effusion|5419,5427
with|5428,5432
adjacent|5433,5441
atelectasis|5442,5453
.|5453,5454
<EOL>|5456,5457
3|5457,5458
.|5458,5459
Possible|5461,5469
calcified|5470,5479
splenic|5480,5487
artery|5488,5494
aneurysm|5495,5503
in|5504,5506
the|5507,5510
region|5511,5517
of|5518,5520
<EOL>|5521,5522
the|5522,5525
hilum|5526,5531
.|5531,5532
<EOL>|5533,5534
<EOL>|5534,5535
Cardiac|5535,5542
catheterization|5543,5558
_|5559,5560
_|5560,5561
_|5561,5562
.|5562,5563
Selective|5564,5573
coronary|5574,5582
angiography|5583,5594
of|5595,5597
this|5598,5602
right|5603,5608
dominant|5609,5617
system|5618,5624
<EOL>|5625,5626
demonstrated|5626,5638
2|5639,5640
vessel|5641,5647
coronary|5648,5656
disease|5657,5664
in|5665,5667
the|5668,5671
native|5672,5678
vessels|5679,5686
.|5686,5687
<EOL>|5689,5690
The|5690,5693
_|5694,5695
_|5695,5696
_|5696,5697
<EOL>|5698,5699
had|5699,5702
no|5703,5705
angiographically|5706,5722
apparent|5723,5731
disease|5732,5739
.|5739,5740
The|5742,5745
LAD|5746,5749
had|5750,5753
a|5754,5755
70|5756,5758
%|5758,5759
<EOL>|5760,5761
lesion|5761,5767
in|5768,5770
a|5771,5772
<EOL>|5773,5774
prior|5774,5779
stent|5780,5785
,|5785,5786
and|5787,5790
a|5791,5792
jailed|5793,5799
diagnoal|5800,5808
which|5809,5814
was|5815,5818
small|5819,5824
and|5825,5828
had|5829,5832
poor|5833,5837
<EOL>|5838,5839
flow|5839,5843
.|5843,5844
<EOL>|5845,5846
The|5846,5849
LCx|5850,5853
had|5854,5857
a|5858,5859
70|5860,5862
-|5862,5863
80|5863,5865
%|5865,5866
stenosis|5867,5875
at|5876,5878
its|5879,5882
origin|5883,5889
.|5889,5890
The|5892,5895
RCA|5896,5899
had|5900,5903
no|5904,5906
<EOL>|5907,5908
angiographically|5908,5924
apparent|5925,5933
disease|5934,5941
.|5941,5942
<EOL>|5943,5944
2.|5944,5946
Arterial|5947,5955
conduit|5956,5963
angiography|5964,5975
demonstrated|5976,5988
the|5989,5992
LIMA|5993,5997
graft|5998,6003
to|6004,6006
<EOL>|6007,6008
be|6008,6010
<EOL>|6011,6012
patent|6012,6018
.|6018,6019
<EOL>|6020,6021
3.|6021,6023
Venous|6024,6030
conduit|6031,6038
angiography|6039,6050
demonstrated|6051,6063
a|6064,6065
patent|6066,6072
SVG|6073,6076
to|6077,6079
OM|6080,6082
<EOL>|6083,6084
with|6084,6088
<EOL>|6089,6090
retrograde|6090,6100
stenosis|6101,6109
involving|6110,6119
a|6120,6121
small|6122,6127
sub-branch|6128,6138
of|6139,6141
the|6142,6145
OM|6146,6148
.|6148,6149
The|6151,6154
<EOL>|6155,6156
SVG|6156,6159
to|6160,6162
<EOL>|6163,6164
small|6164,6169
diagonal|6170,6178
was|6179,6182
presumed|6183,6191
occluded|6192,6200
and|6201,6204
unable|6205,6211
to|6212,6214
be|6215,6217
<EOL>|6218,6219
identified|6219,6229
.|6229,6230
<EOL>|6231,6232
4.|6232,6234
Limited|6235,6242
resting|6243,6250
hemodynamics|6251,6263
revealed|6264,6272
systemic|6273,6281
hypertension|6282,6294
<EOL>|6295,6296
with|6296,6300
<EOL>|6301,6302
aortic|6302,6308
pressure|6309,6317
of|6318,6320
184|6321,6324
/|6324,6325
105|6325,6328
mm|6329,6331
Hg|6332,6334
.|6334,6335
<EOL>|6336,6337
FINAL|6339,6344
DIAGNOSIS|6345,6354
:|6354,6355
<EOL>|6360,6361
1|6361,6362
.|6362,6363
Two|6364,6367
vessel|6368,6374
coronary|6375,6383
artery|6384,6390
disease|6391,6398
in|6399,6401
the|6402,6405
native|6406,6412
arteries|6413,6421
<EOL>|6422,6423
2.|6423,6425
Patent|6426,6432
LIMA|6433,6437
to|6438,6440
LAD|6441,6444
,|6444,6445
patent|6446,6452
SVG|6453,6456
to|6457,6459
OM|6460,6462
,|6462,6463
occluded|6464,6472
SVG|6473,6476
to|6477,6479
small|6480,6485
<EOL>|6486,6487
diagonal|6487,6495
<EOL>|6496,6497
branch|6497,6503
.|6503,6504
<EOL>|6505,6506
<EOL>|6506,6507
<EOL>|6508,6509
Brief|6509,6514
Hospital|6515,6523
Course|6524,6530
:|6530,6531
<EOL>|6531,6532
_|6532,6533
_|6533,6534
_|6534,6535
year|6536,6540
old|6541,6544
female|6545,6551
with|6552,6556
a|6557,6558
history|6559,6566
of|6567,6569
CAD|6570,6573
s|6574,6575
/|6575,6576
p|6576,6577
PCI|6578,6581
x3|6582,6584
,|6584,6585
s|6586,6587
/|6587,6588
p|6588,6589
CABG|6590,6594
x3|6595,6597
<EOL>|6598,6599
(|6599,6600
_|6600,6601
_|6601,6602
_|6602,6603
)|6603,6604
,|6604,6605
type|6606,6610
2|6611,6612
DM|6613,6615
on|6616,6618
insulin|6619,6626
,|6626,6627
HTN|6628,6631
,|6631,6632
and|6633,6636
HLD|6637,6640
who|6641,6644
presented|6645,6654
with|6655,6659
<EOL>|6660,6661
a|6661,6662
3|6663,6664
day|6665,6668
history|6669,6676
of|6677,6679
left|6680,6684
sided|6685,6690
chest|6691,6696
pain|6697,6701
and|6702,6705
SOB|6706,6709
.|6709,6710
<EOL>|6712,6713
<EOL>|6713,6714
#|6714,6715
Chest|6716,6721
Pain|6722,6726
-|6726,6727
Patient|6728,6735
with|6736,6740
significant|6741,6752
CAD|6753,6756
history|6757,6764
,|6764,6765
s|6766,6767
/|6767,6768
p|6768,6769
recent|6770,6776
<EOL>|6777,6778
CABG|6778,6782
,|6782,6783
presenting|6784,6794
with|6795,6799
chest|6800,6805
pain|6806,6810
and|6811,6814
rising|6815,6821
troponins|6822,6831
,|6831,6832
with|6833,6837
new|6838,6841
<EOL>|6842,6843
ST|6843,6845
depressions|6846,6857
inferiorly|6858,6868
in|6869,6871
V4|6872,6874
-|6874,6875
V6|6875,6877
,|6877,6878
consistent|6879,6889
with|6890,6894
NSTEMI|6895,6901
.|6901,6902
<EOL>|6904,6905
Patient|6905,6912
's|6912,6914
troponins|6915,6924
plateaued|6925,6934
at|6935,6937
0.13|6938,6942
.|6942,6943
She|6945,6948
has|6949,6952
initiated|6953,6962
on|6963,6965
a|6966,6967
<EOL>|6968,6969
heparin|6969,6976
gtt|6977,6980
in|6981,6983
the|6984,6987
ED|6988,6990
,|6990,6991
and|6992,6995
was|6996,6999
taken|7000,7005
to|7006,7008
cardiac|7009,7016
cath|7017,7021
the|7022,7025
<EOL>|7026,7027
following|7027,7036
morning|7037,7044
.|7044,7045
Catheterization|7047,7062
showed|7063,7069
occlusion|7070,7079
of|7080,7082
the|7083,7086
SVG|7087,7090
<EOL>|7091,7092
to|7092,7094
the|7095,7098
diagonal|7099,7107
,|7107,7108
possibly|7109,7117
causing|7118,7125
her|7126,7129
current|7130,7137
symptoms|7138,7146
.|7146,7147
No|7149,7151
<EOL>|7152,7153
intervention|7153,7165
was|7166,7169
performed|7170,7179
.|7179,7180
Patient|7182,7189
was|7190,7193
medically|7194,7203
optimized|7204,7213
<EOL>|7214,7215
with|7215,7219
increased|7220,7229
metoprolol|7230,7240
,|7240,7241
initiation|7242,7252
of|7253,7255
losartan|7256,7264
,|7264,7265
and|7266,7269
<EOL>|7270,7271
initiation|7271,7281
of|7282,7284
imdur|7285,7290
.|7290,7291
Other|7293,7298
potential|7299,7308
causes|7309,7315
of|7316,7318
her|7319,7322
chest|7323,7328
pain|7329,7333
<EOL>|7334,7335
were|7335,7339
considered|7340,7350
including|7351,7360
PE|7361,7363
(|7364,7365
ruled|7365,7370
out|7371,7374
with|7375,7379
negative|7380,7388
CTA|7389,7392
)|7392,7393
,|7393,7394
<EOL>|7395,7396
pericarditis|7396,7408
(|7409,7410
symptoms|7410,7418
consistent|7419,7429
,|7429,7430
but|7431,7434
exam|7435,7439
and|7440,7443
EKG|7444,7447
not|7448,7451
<EOL>|7452,7453
consistent|7453,7463
,|7463,7464
also|7465,7469
patient|7470,7477
has|7478,7481
been|7482,7486
essentially|7487,7498
treated|7499,7506
as|7507,7509
she|7510,7513
has|7514,7517
<EOL>|7518,7519
been|7519,7523
taking|7524,7530
consistent|7531,7541
NSAIDs|7542,7548
)|7548,7549
,|7549,7550
costochondritis|7551,7566
(|7567,7568
symptoms|7568,7576
<EOL>|7577,7578
intermittently|7578,7592
reproducible|7593,7605
on|7606,7608
exam|7609,7613
)|7613,7614
,|7614,7615
or|7616,7618
pleuritis|7619,7628
secondary|7629,7638
to|7639,7641
<EOL>|7642,7643
pleural|7643,7650
effusion|7651,7659
(|7660,7661
very|7661,7665
small|7666,7671
effusion|7672,7680
,|7680,7681
stable|7682,7688
since|7689,7694
CABG|7695,7699
)|7699,7700
.|7700,7701
<EOL>|7703,7704
If|7707,7709
pain|7710,7714
persists|7715,7723
,|7723,7724
patient|7725,7732
was|7733,7736
instructed|7737,7747
to|7748,7750
speak|7751,7756
with|7757,7761
her|7762,7765
<EOL>|7766,7767
cardiologist|7767,7779
about|7780,7785
increasing|7786,7796
imdur|7797,7802
should|7803,7809
her|7810,7813
blood|7814,7819
pressure|7820,7828
<EOL>|7829,7830
tolerate|7830,7838
.|7838,7839
<EOL>|7841,7842
<EOL>|7844,7845
#|7845,7846
Acute|7847,7852
renal|7853,7858
insufficiency|7859,7872
-|7872,7873
On|7874,7876
admission|7877,7886
,|7886,7887
creatinine|7888,7898
elevated|7899,7907
<EOL>|7908,7909
to|7909,7911
1.2|7912,7915
,|7915,7916
likely|7917,7923
due|7924,7927
to|7928,7930
dehydration|7931,7942
,|7942,7943
as|7944,7946
creatinine|7947,7957
improved|7958,7966
<EOL>|7967,7968
overnight|7968,7977
with|7978,7982
gentle|7983,7989
fluids|7990,7996
and|7997,8000
remained|8001,8009
stable|8010,8016
.|8016,8017
<EOL>|8018,8019
<EOL>|8019,8020
#|8020,8021
COPD|8022,8026
-|8026,8027
Continued|8028,8037
on|8038,8040
home|8041,8045
inhalers|8046,8054
(|8055,8056
albuterol|8056,8065
,|8065,8066
fluticasone|8067,8078
)|8078,8079
<EOL>|8079,8080
<EOL>|8080,8081
#|8081,8082
DM|8083,8085
-|8085,8086
Continued|8087,8096
with|8097,8101
glargine|8102,8110
50|8111,8113
units|8114,8119
Q6|8120,8122
and|8123,8126
ISS|8127,8130
<EOL>|8132,8133
<EOL>|8133,8134
#|8134,8135
HLD|8136,8139
-|8139,8140
Continued|8141,8150
on|8151,8153
home|8154,8158
atorvastatin|8159,8171
<EOL>|8172,8173
<EOL>|8173,8174
#|8174,8175
GERD|8176,8180
-|8180,8181
Continued|8182,8191
on|8192,8194
home|8195,8199
pantoprazole|8200,8212
<EOL>|8212,8213
<EOL>|8213,8214
#|8214,8215
Transitional|8216,8228
issues|8229,8235
-|8235,8236
<EOL>|8236,8237
-|8237,8238
NEW|8239,8242
MEDICATIONS|8243,8254
-|8254,8255
losartan|8256,8264
and|8265,8268
imdur|8269,8274
<EOL>|8274,8275
-|8275,8276
MEDICATION|8277,8287
CHANGES|8288,8295
-|8295,8296
metoprolol|8297,8307
increased|8308,8317
to|8318,8320
50mg|8321,8325
po|8326,8328
TID|8329,8332
(|8333,8334
from|8334,8338
<EOL>|8339,8340
25|8340,8342
TID|8343,8346
)|8346,8347
<EOL>|8347,8348
-|8348,8349
if|8350,8352
ongoing|8353,8360
chest|8361,8366
pain|8367,8371
,|8371,8372
consider|8373,8381
titrating|8382,8391
up|8392,8394
on|8395,8397
imdur|8398,8403
if|8404,8406
c|8407,8408
/|8408,8409
w|8409,8410
<EOL>|8411,8412
anginal|8412,8419
pain|8420,8424
.|8424,8425
Also|8428,8432
may|8433,8436
consider|8437,8445
treating|8446,8454
for|8455,8458
costochondritis|8459,8474
<EOL>|8475,8476
and|8476,8479
pericarditis|8480,8492
<EOL>|8492,8493
<EOL>|8494,8495
Medications|8495,8506
on|8507,8509
Admission|8510,8519
:|8519,8520
<EOL>|8520,8521
The|8521,8524
Preadmission|8525,8537
Medication|8538,8548
list|8549,8553
is|8554,8556
accurate|8557,8565
and|8566,8569
complete|8570,8578
.|8578,8579
<EOL>|8579,8580
1.|8580,8582
Albuterol|8583,8592
Inhaler|8593,8600
2|8601,8602
PUFF|8603,8607
IH|8608,8610
Q6H|8611,8614
:|8614,8615
PRN|8615,8618
SOB|8619,8622
<EOL>|8623,8624
2.|8624,8626
Atorvastatin|8627,8639
40|8640,8642
mg|8643,8645
PO|8646,8648
DAILY|8649,8654
<EOL>|8655,8656
3.|8656,8658
Clopidogrel|8659,8670
75|8671,8673
mg|8674,8676
PO|8677,8679
DAILY|8680,8685
<EOL>|8686,8687
4.|8687,8689
Fluticasone|8690,8701
Propionate|8702,8712
110mcg|8713,8719
2|8720,8721
PUFF|8722,8726
IH|8727,8729
BID|8730,8733
<EOL>|8734,8735
5.|8735,8737
Glargine|8738,8746
50|8747,8749
Units|8750,8755
Bedtime|8756,8763
<EOL>|8763,8764
Insulin|8764,8771
SC|8772,8774
Sliding|8775,8782
Scale|8783,8788
using|8789,8794
HUM|8795,8798
Insulin|8799,8806
<EOL>|8806,8807
6.|8807,8809
Metoprolol|8810,8820
Tartrate|8821,8829
25|8830,8832
mg|8833,8835
PO|8836,8838
TID|8839,8842
<EOL>|8843,8844
Hold|8844,8848
for|8849,8852
SBP|8853,8856
<|8857,8858
100|8858,8861
,|8861,8862
HR|8863,8865
<|8865,8866
60|8866,8868
<EOL>|8869,8870
7.|8870,8872
Metrogel|8873,8881
*|8882,8883
NF|8883,8885
*|8885,8886
(|8887,8888
metroNIDAZOLE|8888,8901
)|8901,8902
0.75|8903,8907
%|8907,8908
Topical|8910,8917
Daily|8918,8923
<EOL>|8924,8925
8.|8925,8927
Oxycodone|8928,8937
-|8937,8938
Acetaminophen|8938,8951
(|8952,8953
5mg|8953,8956
-|8956,8957
325mg|8957,8962
)|8962,8963
1|8964,8965
TAB|8966,8969
PO|8970,8972
Q8H|8973,8976
:|8976,8977
PRN|8977,8980
severe|8981,8987
<EOL>|8988,8989
pain|8989,8993
<EOL>|8994,8995
9.|8995,8997
Pantoprazole|8998,9010
80|9011,9013
mg|9014,9016
PO|9017,9019
Q24H|9020,9024
<EOL>|9025,9026
10.|9026,9029
Ropinirole|9030,9040
0.25|9041,9045
mg|9046,9048
PO|9049,9051
QPM|9052,9055
<EOL>|9056,9057
11.|9057,9060
Aspirin|9061,9068
325|9069,9072
mg|9073,9075
PO|9076,9078
DAILY|9079,9084
<EOL>|9085,9086
12.|9086,9089
Vitamin|9090,9097
D|9098,9099
1000|9100,9104
UNIT|9105,9109
PO|9110,9112
DAILY|9113,9118
<EOL>|9119,9120
13.|9120,9123
Ibuprofen|9124,9133
600|9134,9137
mg|9138,9140
PO|9141,9143
Q6H|9144,9147
:|9147,9148
PRN|9148,9151
pain|9152,9156
<EOL>|9157,9158
<EOL>|9158,9159
<EOL>|9160,9161
Discharge|9161,9170
Medications|9171,9182
:|9182,9183
<EOL>|9183,9184
1.|9184,9186
Albuterol|9187,9196
Inhaler|9197,9204
2|9205,9206
PUFF|9207,9211
IH|9212,9214
Q6H|9215,9218
:|9218,9219
PRN|9219,9222
SOB|9223,9226
<EOL>|9227,9228
2.|9228,9230
Aspirin|9231,9238
81|9239,9241
mg|9242,9244
PO|9245,9247
DAILY|9248,9253
<EOL>|9254,9255
RX|9255,9257
*|9258,9259
aspirin|9259,9266
81|9267,9269
mg|9270,9272
1|9273,9274
tablet|9275,9281
(|9281,9282
s|9282,9283
)|9283,9284
by|9285,9287
mouth|9288,9293
daily|9294,9299
Disp|9300,9304
#|9305,9306
*|9306,9307
30|9307,9309
Tablet|9310,9316
<EOL>|9317,9318
Refills|9318,9325
:|9325,9326
*|9326,9327
0|9327,9328
<EOL>|9328,9329
3.|9329,9331
Atorvastatin|9332,9344
80|9345,9347
mg|9348,9350
PO|9351,9353
DAILY|9354,9359
<EOL>|9360,9361
RX|9361,9363
*|9364,9365
atorvastatin|9365,9377
80|9378,9380
mg|9381,9383
1|9384,9385
tablet|9386,9392
(|9392,9393
s|9393,9394
)|9394,9395
by|9396,9398
mouth|9399,9404
daily|9405,9410
Disp|9411,9415
#|9416,9417
*|9417,9418
30|9418,9420
<EOL>|9421,9422
Tablet|9422,9428
Refills|9429,9436
:|9436,9437
*|9437,9438
0|9438,9439
<EOL>|9439,9440
4.|9440,9442
Glargine|9443,9451
50|9452,9454
Units|9455,9460
Bedtime|9461,9468
<EOL>|9468,9469
Insulin|9469,9476
SC|9477,9479
Sliding|9480,9487
Scale|9488,9493
using|9494,9499
HUM|9500,9503
Insulin|9504,9511
<EOL>|9511,9512
5.|9512,9514
Metoprolol|9515,9525
Tartrate|9526,9534
50|9535,9537
mg|9538,9540
PO|9541,9543
TID|9544,9547
<EOL>|9548,9549
RX|9549,9551
*|9552,9553
metoprolol|9553,9563
tartrate|9564,9572
50|9573,9575
mg|9576,9578
1|9579,9580
tablet|9581,9587
(|9587,9588
s|9588,9589
)|9589,9590
by|9591,9593
mouth|9594,9599
three|9600,9605
times|9606,9611
a|9612,9613
<EOL>|9614,9615
day|9615,9618
Disp|9619,9623
#|9624,9625
*|9625,9626
90|9626,9628
Tablet|9629,9635
Refills|9636,9643
:|9643,9644
*|9644,9645
0|9645,9646
<EOL>|9646,9647
6.|9647,9649
Pantoprazole|9650,9662
40|9663,9665
mg|9666,9668
PO|9669,9671
Q24H|9672,9676
<EOL>|9677,9678
RX|9678,9680
*|9681,9682
pantoprazole|9682,9694
40|9695,9697
mg|9698,9700
1|9701,9702
tablet|9703,9709
(|9709,9710
s|9710,9711
)|9711,9712
by|9713,9715
mouth|9716,9721
daily|9722,9727
Disp|9728,9732
#|9733,9734
*|9734,9735
30|9735,9737
<EOL>|9738,9739
Tablet|9739,9745
Refills|9746,9753
:|9753,9754
*|9754,9755
0|9755,9756
<EOL>|9756,9757
7.|9757,9759
Ropinirole|9760,9770
0.25|9771,9775
mg|9776,9778
PO|9779,9781
QPM|9782,9785
<EOL>|9786,9787
8.|9787,9789
Vitamin|9790,9797
D|9798,9799
1000|9800,9804
UNIT|9805,9809
PO|9810,9812
DAILY|9813,9818
<EOL>|9819,9820
9.|9820,9822
Isosorbide|9823,9833
Mononitrate|9834,9845
(|9846,9847
Extended|9847,9855
Release|9856,9863
)|9863,9864
30|9865,9867
mg|9868,9870
PO|9871,9873
DAILY|9874,9879
<EOL>|9880,9881
RX|9881,9883
*|9884,9885
isosorbide|9885,9895
mononitrate|9896,9907
30|9908,9910
mg|9911,9913
1|9914,9915
tablet|9916,9922
(|9922,9923
s|9923,9924
)|9924,9925
by|9926,9928
mouth|9929,9934
daily|9935,9940
Disp|9941,9945
<EOL>|9946,9947
#|9947,9948
*|9948,9949
30|9949,9951
Tablet|9952,9958
Refills|9959,9966
:|9966,9967
*|9967,9968
0|9968,9969
<EOL>|9969,9970
10.|9970,9973
Metrogel|9974,9982
*|9983,9984
NF|9984,9986
*|9986,9987
(|9988,9989
metroNIDAZOLE|9989,10002
)|10002,10003
0.75|10004,10008
%|10008,10009
Topical|10011,10018
Daily|10019,10024
<EOL>|10025,10026
11|10026,10028
.|10028,10029
Oxycodone|10030,10039
-|10039,10040
Acetaminophen|10040,10053
(|10054,10055
5mg|10055,10058
-|10058,10059
325mg|10059,10064
)|10064,10065
1|10066,10067
TAB|10068,10071
PO|10072,10074
Q8H|10075,10078
:|10078,10079
PRN|10079,10082
severe|10083,10089
<EOL>|10090,10091
pain|10091,10095
<EOL>|10096,10097
12.|10097,10100
Losartan|10101,10109
Potassium|10110,10119
25|10120,10122
mg|10123,10125
PO|10126,10128
DAILY|10129,10134
<EOL>|10135,10136
RX|10136,10138
*|10139,10140
losartan|10140,10148
25|10149,10151
mg|10152,10154
1|10155,10156
tablet|10157,10163
(|10163,10164
s|10164,10165
)|10165,10166
by|10167,10169
mouth|10170,10175
daily|10176,10181
Disp|10182,10186
#|10187,10188
*|10188,10189
30|10189,10191
Tablet|10192,10198
<EOL>|10199,10200
Refills|10200,10207
:|10207,10208
*|10208,10209
0|10209,10210
<EOL>|10210,10211
13.|10211,10214
Clopidogrel|10215,10226
75|10227,10229
mg|10230,10232
PO|10233,10235
DAILY|10236,10241
<EOL>|10242,10243
14.|10243,10246
Fluticasone|10247,10258
Propionate|10259,10269
110mcg|10270,10276
2|10277,10278
PUFF|10279,10283
IH|10284,10286
BID|10287,10290
<EOL>|10291,10292
<EOL>|10292,10293
<EOL>|10294,10295
Discharge|10295,10304
Disposition|10305,10316
:|10316,10317
<EOL>|10317,10318
Home|10318,10322
<EOL>|10322,10323
<EOL>|10324,10325
Discharge|10325,10334
Diagnosis|10335,10344
:|10344,10345
<EOL>|10345,10346
Primary|10346,10353
:|10353,10354
<EOL>|10354,10355
non-ST|10355,10361
elevation|10362,10371
MI|10372,10374
<EOL>|10374,10375
coronary|10375,10383
artery|10384,10390
disease|10391,10398
<EOL>|10398,10399
<EOL>|10399,10400
Secondary|10400,10409
:|10409,10410
<EOL>|10410,10411
diabetes|10411,10419
mellitus|10420,10428
type|10429,10433
2|10434,10435
<EOL>|10435,10436
hypertension|10436,10448
<EOL>|10448,10449
hyperlipidemia|10449,10463
<EOL>|10463,10464
<EOL>|10464,10465
<EOL>|10466,10467
Discharge|10467,10476
Condition|10477,10486
:|10486,10487
<EOL>|10487,10488
Mental|10488,10494
Status|10495,10501
:|10501,10502
Clear|10503,10508
and|10509,10512
coherent|10513,10521
.|10521,10522
<EOL>|10522,10523
Level|10523,10528
of|10529,10531
Consciousness|10532,10545
:|10545,10546
Alert|10547,10552
and|10553,10556
interactive|10557,10568
.|10568,10569
<EOL>|10569,10570
Activity|10570,10578
Status|10579,10585
:|10585,10586
Ambulatory|10587,10597
-|10598,10599
Independent|10600,10611
.|10611,10612
<EOL>|10612,10613
<EOL>|10613,10614
<EOL>|10615,10616
Discharge|10616,10625
Instructions|10626,10638
:|10638,10639
<EOL>|10639,10640
It|10640,10642
was|10643,10646
a|10647,10648
pleasure|10649,10657
taking|10658,10664
care|10665,10669
of|10670,10672
you|10673,10676
during|10677,10683
your|10684,10688
recent|10689,10695
<EOL>|10696,10697
admission|10697,10706
to|10707,10709
_|10710,10711
_|10711,10712
_|10712,10713
.|10713,10714
<EOL>|10714,10715
<EOL>|10715,10716
You|10716,10719
were|10720,10724
admitted|10725,10733
with|10734,10738
chest|10739,10744
pain|10745,10749
/|10749,10750
pressure|10750,10758
concerning|10759,10769
for|10770,10773
a|10774,10775
<EOL>|10776,10777
heart|10777,10782
attack|10783,10789
.|10789,10790
A|10792,10793
cardiac|10794,10801
catheterization|10802,10817
showed|10818,10824
that|10825,10829
one|10830,10833
of|10834,10836
your|10837,10841
<EOL>|10842,10843
grafts|10843,10849
from|10850,10854
your|10855,10859
recent|10860,10866
cardiac|10867,10874
bypass|10875,10881
surgery|10882,10889
is|10890,10892
clotted|10893,10900
and|10901,10904
no|10905,10907
<EOL>|10908,10909
longer|10909,10915
working|10916,10923
,|10923,10924
potentially|10925,10936
causing|10937,10944
your|10945,10949
symptoms|10950,10958
.|10958,10959
<EOL>|10961,10962
<EOL>|10962,10963
We|10963,10965
have|10966,10970
increased|10971,10980
and|10981,10984
added|10985,10990
medications|10991,11002
to|11003,11005
control|11006,11013
your|11014,11018
<EOL>|11019,11020
symptoms|11020,11028
.|11028,11029
The|11031,11034
changes|11035,11042
are|11043,11046
below|11047,11052
:|11052,11053
<EOL>|11053,11054
START|11054,11059
losartan|11060,11068
<EOL>|11068,11069
START|11069,11074
isosorbide|11075,11085
mononitrate|11086,11097
<EOL>|11097,11098
INCREASE|11098,11106
atorvastatin|11107,11119
<EOL>|11119,11120
INCREASE|11120,11128
metoprolol|11129,11139
<EOL>|11139,11140
DECREASE|11140,11148
aspirin|11149,11156
<EOL>|11156,11157
DECREASE|11157,11165
pantoprazole|11166,11178
<EOL>|11178,11179
STOP|11179,11183
ibuprofen|11184,11193
(|11194,11195
you|11195,11198
were|11199,11203
taking|11204,11210
too|11211,11214
much|11215,11219
.|11219,11220
take|11221,11225
tylenol|11226,11233
_|11234,11235
_|11235,11236
_|11236,11237
for|11238,11241
<EOL>|11242,11243
pain|11243,11247
)|11247,11248
<EOL>|11248,11249
<EOL>|11249,11250
Once|11250,11254
you|11255,11258
leave|11259,11264
the|11265,11268
hospital|11269,11277
,|11277,11278
we|11279,11281
recommend|11282,11291
further|11292,11299
workup|11300,11306
of|11307,11309
a|11310,11311
<EOL>|11312,11313
fluid|11313,11318
collection|11319,11329
seen|11330,11334
around|11335,11341
your|11342,11346
left|11347,11351
lung|11352,11356
and|11357,11360
better|11361,11367
<EOL>|11368,11369
management|11369,11379
of|11380,11382
your|11383,11387
diabetes|11388,11396
with|11397,11401
the|11402,11405
help|11406,11410
of|11411,11413
your|11414,11418
PCP|11419,11422
.|11422,11423
<EOL>|11423,11424
<EOL>|11425,11426
Followup|11426,11434
Instructions|11435,11447
:|11447,11448
<EOL>|11448,11449
_|11449,11450
_|11450,11451
_|11451,11452
<EOL>|11452,11453

