 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|158,166|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|169,178|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|169,178|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|169,178|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|190,199|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|190,199|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|190,199|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|202,224|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|210,214|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|210,214|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|210,224|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|215,224|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|227,236|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|227,236|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|245,260|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|251,260|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|251,260|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|251,260|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|262,267|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|262,267|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|262,267|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Classification|SIMPLE_SEGMENT|270,275|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|276,284|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|276,284|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|288,306|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|297,306|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|297,306|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|297,306|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|297,306|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|297,306|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|316,323|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|316,326|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|316,342|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|316,342|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|327,334|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|327,334|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|327,342|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|335,342|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|353,360|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|353,360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|353,360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|353,360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|353,363|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|364,378|false|false|false|C0028756|Morbid obesity|morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|371,378|false|false|false|C0028754|Obesity|obesity
Event|Event|SIMPLE_SEGMENT|371,378|false|false|false|||obesity
Finding|Finding|SIMPLE_SEGMENT|371,378|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|380,388|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|380,395|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|380,403|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|389,395|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|389,395|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|389,403|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|396,403|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|396,403|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|406,416|false|false|false|||presenting
Drug|Organic Chemical|SIMPLE_SEGMENT|428,433|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|428,433|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|428,433|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|428,433|false|false|false|C0010200|Coughing|cough
Finding|Finding|SIMPLE_SEGMENT|428,444|false|false|false|C0239134|Productive Cough|cough productive
Event|Event|SIMPLE_SEGMENT|434,444|false|false|false|||productive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|448,453|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Finding|Finding|SIMPLE_SEGMENT|448,460|false|false|false|C0457099|Brown sputum|brown sputum
Event|Event|SIMPLE_SEGMENT|454,460|false|false|false|||sputum
Finding|Body Substance|SIMPLE_SEGMENT|454,460|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|454,460|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|466,472|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|466,472|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|507,515|false|false|false|||endorses
Event|Event|SIMPLE_SEGMENT|516,522|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|516,522|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|525,532|false|false|false|||Husband
Event|Event|SIMPLE_SEGMENT|546,554|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|546,554|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|546,554|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|569,578|false|false|false|||improving
Drug|Antibiotic|SIMPLE_SEGMENT|588,599|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|588,599|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|601,607|false|false|false|||Denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|612,617|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|612,617|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|612,622|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|612,622|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|618,622|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|618,622|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|618,622|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|618,622|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|627,633|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|661,666|false|false|false|||short
Finding|Sign or Symptom|SIMPLE_SEGMENT|661,676|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|670,676|false|false|false|C0225386|Breath|breath
Finding|Idea or Concept|SIMPLE_SEGMENT|693,700|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|732,735|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|732,735|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|736,742|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|758,768|false|false|false|||prominence
Event|Event|SIMPLE_SEGMENT|776,784|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|776,784|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|776,787|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|788,791|true|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|788,791|true|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|795,804|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|795,804|false|false|false|||pneumonia
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|806,810|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Drug|Enzyme|SIMPLE_SEGMENT|806,810|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Event|Event|SIMPLE_SEGMENT|809,810|false|false|false|||A
Event|Event|SIMPLE_SEGMENT|814,820|false|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|824,829|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|830,839|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|840,847|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|840,847|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|840,847|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|840,847|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|840,847|false|false|false|C1522240|Process|process
Event|Event|SIMPLE_SEGMENT|849,853|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|849,853|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|854,861|false|false|false|||notable
Anatomy|Cell|SIMPLE_SEGMENT|866,869|false|false|false|C0023516|Leukocytes|WBC
Drug|Organic Chemical|SIMPLE_SEGMENT|900,907|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|900,907|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|900,907|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|900,907|false|false|false|C0202115|Lactic acid measurement|lactate
Finding|Functional Concept|SIMPLE_SEGMENT|919,924|false|false|false|C1883002|Sequence Chromatogram|trace
Event|Event|SIMPLE_SEGMENT|925,930|false|false|false|||leuks
Finding|Intellectual Product|SIMPLE_SEGMENT|939,947|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|SIMPLE_SEGMENT|948,955|false|false|false|||picture
Event|Event|SIMPLE_SEGMENT|960,965|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|960,965|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|960,965|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Body Substance|SIMPLE_SEGMENT|967,974|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|967,974|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|967,974|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|979,986|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|991,1002|false|false|false|||presumptive
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1004,1007|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|1004,1007|false|false|false|||PNA
Drug|Antibiotic|SIMPLE_SEGMENT|1013,1025|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|1013,1025|false|false|false|C0282386|levofloxacin|Levofloxacin
Event|Event|SIMPLE_SEGMENT|1013,1025|false|false|false|||Levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|1055,1061|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1055,1061|false|false|false|C0699194|Ativan|Ativan
Drug|Organic Chemical|SIMPLE_SEGMENT|1071,1078|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1071,1078|false|false|false|C0699142|Tylenol|Tylenol
Drug|Organic Chemical|SIMPLE_SEGMENT|1083,1089|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1083,1089|false|false|false|C0206046|Zofran|Zofran
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1095,1099|false|false|false|C2317096|Saturation of Peripheral Oxygen|SpO2
Event|Event|SIMPLE_SEGMENT|1100,1107|false|false|false|||dropped
Event|Event|SIMPLE_SEGMENT|1120,1130|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1120,1130|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|1120,1130|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|SIMPLE_SEGMENT|1147,1153|false|false|false|||wanted
Event|Event|SIMPLE_SEGMENT|1157,1162|false|false|false|||leave
Event|Event|SIMPLE_SEGMENT|1172,1181|false|false|false|||convinced
Event|Event|SIMPLE_SEGMENT|1185,1189|false|false|false|||stay
Event|Event|SIMPLE_SEGMENT|1198,1206|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1198,1206|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1198,1206|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1198,1206|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1258,1263|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|1258,1263|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|1258,1263|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|1258,1263|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|1268,1274|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1279,1282|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1279,1282|true|false|false|C0013404|Dyspnea|SOB
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1290,1293|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1290,1293|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1290,1293|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|SIMPLE_SEGMENT|1290,1293|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1290,1293|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|SIMPLE_SEGMENT|1290,1293|false|false|false|||ROS
Finding|Gene or Genome|SIMPLE_SEGMENT|1290,1293|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|SIMPLE_SEGMENT|1290,1293|false|false|false|C0489633|Review of systems (procedure)|ROS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1302,1305|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|1302,1305|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|1302,1305|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|1302,1305|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Finding|SIMPLE_SEGMENT|1311,1331|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1316,1323|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1316,1323|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1316,1323|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1316,1323|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1316,1323|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1316,1331|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1324,1331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1324,1331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1324,1331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Tissue|SIMPLE_SEGMENT|1333,1343|false|false|false|C0027061|Myocardium|MYOCARDIAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1333,1351|false|false|false|C0027051|Myocardial Infarction|MYOCARDIAL INFARCT
Event|Event|SIMPLE_SEGMENT|1344,1351|false|false|false|||INFARCT
Finding|Pathologic Function|SIMPLE_SEGMENT|1344,1351|false|false|false|C0021308|Infarction|INFARCT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1372,1392|false|false|false|C0020443|Hypercholesterolemia|HYPERCHOLESTEROLEMIA
Event|Event|SIMPLE_SEGMENT|1372,1392|false|false|false|||HYPERCHOLESTEROLEMIA
Finding|Finding|SIMPLE_SEGMENT|1372,1392|false|false|false|C1522133|Hypercholesterolemia result|HYPERCHOLESTEROLEMIA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1399,1407|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1399,1416|false|false|false|C0011849|Diabetes Mellitus|diabetes mellitus
Event|Event|SIMPLE_SEGMENT|1419,1423|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|1419,1423|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|1419,1423|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|1419,1425|false|false|false|C0441730|Type 2|type 2
Event|Event|SIMPLE_SEGMENT|1427,1439|false|false|false|||uncontrolled
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1442,1454|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|SIMPLE_SEGMENT|1468,1474|false|false|false|||UNSPEC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1477,1483|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|1477,1483|false|false|false|||Anemia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040132|Thyroid Gland|Thyroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040128|Thyroid Diseases|Thyroid
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Hormone|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Organic Chemical|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1486,1493|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Procedure|Health Care Activity|SIMPLE_SEGMENT|1486,1493|false|false|false|C2228489|examination of thyroid|Thyroid
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1486,1500|false|false|false|C0040137|Thyroid Nodule|Thyroid nodule
Finding|Finding|SIMPLE_SEGMENT|1486,1500|false|false|false|C2116082||Thyroid nodule
Event|Event|SIMPLE_SEGMENT|1494,1500|false|false|false|||nodule
Finding|Finding|SIMPLE_SEGMENT|1503,1515|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|Asymptomatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1503,1539|false|false|false|C3494609|Asymptomatic carotid artery stenosis|Asymptomatic carotid artery stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1516,1523|false|false|false|C0007272|Carotid Arteries|carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1516,1530|false|false|false|C0007272;C0162859;C1305384;C4071877|Carotid Arteries;Common carotid artery;Head+Neck>Carotid artery|carotid artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1516,1539|false|false|false|C0007282|Carotid Stenosis|carotid artery stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1524,1530|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|1524,1530|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Pathologic Function|SIMPLE_SEGMENT|1524,1539|false|false|false|C0038449|Stricture of artery|artery stenosis
Event|Event|SIMPLE_SEGMENT|1531,1539|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|1531,1539|false|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1542,1549|false|false|false|C0028754|Obesity|OBESITY
Event|Event|SIMPLE_SEGMENT|1542,1549|false|false|false|||OBESITY
Finding|Finding|SIMPLE_SEGMENT|1542,1549|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|OBESITY
Event|Event|SIMPLE_SEGMENT|1552,1558|false|false|false|||MORBID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1561,1571|false|false|false|C0014852|Esophageal Diseases|ESOPHAGEAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1561,1578|false|false|false|C0017168|Gastroesophageal reflux disease|ESOPHAGEAL REFLUX
Finding|Finding|SIMPLE_SEGMENT|1561,1578|false|false|false|C0559234;C4317146|Acid reflux;Esophageal reflux observation|ESOPHAGEAL REFLUX
Event|Event|SIMPLE_SEGMENT|1572,1578|false|false|false|||REFLUX
Finding|Pathologic Function|SIMPLE_SEGMENT|1572,1578|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1581,1595|false|false|false|C0020676|Hypothyroidism|HYPOTHYROIDISM
Event|Event|SIMPLE_SEGMENT|1581,1595|false|false|false|||HYPOTHYROIDISM
Event|Event|SIMPLE_SEGMENT|1597,1603|false|false|false|||UNSPEC
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1606,1613|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|SIMPLE_SEGMENT|1606,1613|false|false|false|||ANXIETY
Finding|Sign or Symptom|SIMPLE_SEGMENT|1606,1613|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1606,1620|false|false|false|C0700613|Anxiety state|ANXIETY STATES
Event|Event|SIMPLE_SEGMENT|1614,1620|false|false|false|||STATES
Event|Event|SIMPLE_SEGMENT|1622,1628|false|false|false|||UNSPEC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1631,1641|false|false|false|C0011603|Dermatitis|DERMATITIS
Event|Event|SIMPLE_SEGMENT|1631,1641|false|false|false|||DERMATITIS
Event|Event|SIMPLE_SEGMENT|1644,1654|false|false|false|||ECZEMATOUS
Finding|Sign or Symptom|SIMPLE_SEGMENT|1657,1665|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1668,1675|false|false|false|C0009368|Colon structure (body structure)|COLONIC
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1668,1683|false|false|false|C4551463|Colon adenoma|COLONIC ADENOMA
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1676,1683|false|false|false|C0001430|Adenoma|ADENOMA
Event|Event|SIMPLE_SEGMENT|1676,1683|false|false|false|||ADENOMA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1686,1690|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|DISC
Anatomy|Cell Component|SIMPLE_SEGMENT|1686,1690|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|DISC
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1686,1690|false|false|false|C0993608|Disk Drug Form|DISC
Finding|Finding|SIMPLE_SEGMENT|1686,1690|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|DISC
Finding|Intellectual Product|SIMPLE_SEGMENT|1686,1690|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|DISC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1686,1698|false|false|false|C0012619|disc disorder|DISC DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1691,1698|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|1691,1698|false|false|false|||DISEASE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1701,1707|false|false|false|C0024090|Lumbar Region|LUMBAR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1710,1717|false|false|false|C0205065|Ovarian|Ovarian
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1718,1727|false|false|false|C1318143|Retention - dental|Retention
Finding|Cell Function|SIMPLE_SEGMENT|1718,1727|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|Retention
Finding|Functional Concept|SIMPLE_SEGMENT|1718,1727|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|Retention
Finding|Mental Process|SIMPLE_SEGMENT|1718,1727|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|Retention
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1718,1732|false|false|false|C0035281|Retention cyst|Retention Cyst
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1728,1732|false|false|false|C0010709|Cyst|Cyst
Event|Event|SIMPLE_SEGMENT|1728,1732|false|false|false|||Cyst
Finding|Body Substance|SIMPLE_SEGMENT|1728,1732|false|false|false|C1546594;C1550626|SpecimenType - Cyst|Cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|1728,1732|false|false|false|C1546594;C1550626|SpecimenType - Cyst|Cyst
Finding|Functional Concept|SIMPLE_SEGMENT|1742,1748|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1742,1756|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1749,1756|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1749,1756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1749,1756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1749,1756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1762,1768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1762,1768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1762,1768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1762,1768|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1762,1776|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1769,1776|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1769,1776|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1769,1776|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1769,1776|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Activity|SIMPLE_SEGMENT|1782,1794|false|false|false|C1880177|Contribution|contributory
Event|Event|SIMPLE_SEGMENT|1798,1806|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1798,1806|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1798,1806|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1798,1806|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1798,1811|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1798,1811|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1807,1811|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1807,1811|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1807,1811|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1813,1821|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1813,1821|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1813,1821|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1813,1821|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1813,1826|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1813,1826|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1822,1826|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1822,1826|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1822,1826|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1830,1839|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1830,1839|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|1846,1850|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1846,1850|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1846,1850|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|SIMPLE_SEGMENT|1899,1906|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1899,1906|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1899,1906|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1918,1923|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|1918,1923|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1934,1937|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1934,1937|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1934,1937|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1934,1937|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1934,1937|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1934,1937|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1934,1937|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|1939,1950|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1939,1950|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|SIMPLE_SEGMENT|1952,1963|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1967,1972|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|1982,1988|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|1982,1988|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|SIMPLE_SEGMENT|1990,1994|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|2004,2013|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2004,2013|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2036,2041|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2036,2041|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2044,2048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2044,2048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2044,2048|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2051,2057|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|2051,2057|false|false|false|C0332254|Supple|supple
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2062,2073|true|false|false|C0018021|Goiter|thyromegaly
Event|Event|SIMPLE_SEGMENT|2062,2073|false|false|false|||thyromegaly
Event|Event|SIMPLE_SEGMENT|2078,2081|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2078,2081|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2086,2093|false|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|SIMPLE_SEGMENT|2086,2100|true|false|false|C0007280|Carotid bruit|carotid bruits
Event|Event|SIMPLE_SEGMENT|2094,2100|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|2094,2100|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2103,2108|false|false|false|C0024109|Lung|LUNGS
Finding|Pathologic Function|SIMPLE_SEGMENT|2116,2123|false|false|false|C5441917|Distant Metastasis|distant
Finding|Body Substance|SIMPLE_SEGMENT|2124,2130|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2124,2137|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|2131,2137|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2131,2137|false|false|false|C0037709||sounds
Finding|Gene or Genome|SIMPLE_SEGMENT|2149,2152|false|false|false|C1417055|MBNL1 gene|exp
Event|Event|SIMPLE_SEGMENT|2153,2160|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2153,2160|false|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|2166,2174|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2166,2174|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2176,2180|false|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2176,2180|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|SIMPLE_SEGMENT|2181,2190|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|2181,2190|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2195,2211|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|2195,2215|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2205,2211|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2205,2211|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|2212,2215|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2212,2215|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2212,2215|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2218,2223|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2218,2223|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|SIMPLE_SEGMENT|2218,2223|false|false|false|||HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|2218,2223|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|SIMPLE_SEGMENT|2226,2229|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2234,2237|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|2234,2237|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2250,2257|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2250,2257|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2250,2257|false|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2260,2264|false|false|false|||NABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2266,2271|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2266,2271|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2273,2277|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2273,2277|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2288,2294|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|2298,2301|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2298,2301|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2307,2314|false|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|2315,2323|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2315,2323|false|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2326,2337|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|2340,2343|false|false|false|||WWP
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2358,2375|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|SIMPLE_SEGMENT|2369,2375|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2369,2375|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2369,2375|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2369,2375|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|2386,2389|false|false|false|||DPs
Finding|Gene or Genome|SIMPLE_SEGMENT|2386,2389|false|false|false|C1843919|PDSS1 gene|DPs
Anatomy|Body System|SIMPLE_SEGMENT|2394,2398|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|2394,2398|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|2404,2410|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2404,2410|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|2414,2421|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|2414,2421|true|false|false|C0221198|Lesion|lesions
Event|Event|SIMPLE_SEGMENT|2432,2437|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|2432,2437|false|false|false|C0234422|Awake (finding)|awake
Event|Event|SIMPLE_SEGMENT|2448,2456|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2448,2456|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2448,2456|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2448,2456|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2448,2461|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2448,2461|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2457,2461|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2457,2461|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2457,2461|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2465,2474|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|2465,2474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2465,2474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2465,2474|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2465,2474|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|SIMPLE_SEGMENT|2533,2540|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2533,2540|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2533,2540|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2552,2557|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2552,2557|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2568,2571|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2568,2571|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2568,2571|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2568,2571|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2568,2571|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2568,2571|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2568,2571|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|2573,2584|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|2573,2584|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|SIMPLE_SEGMENT|2586,2597|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2601,2606|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2616,2622|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|2616,2622|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|SIMPLE_SEGMENT|2624,2628|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|2638,2647|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2638,2647|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2670,2675|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2670,2675|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2678,2682|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2678,2682|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2678,2682|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2685,2691|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|2685,2691|false|false|false|C0332254|Supple|supple
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2696,2707|true|false|false|C0018021|Goiter|thyromegaly
Event|Event|SIMPLE_SEGMENT|2696,2707|false|false|false|||thyromegaly
Event|Event|SIMPLE_SEGMENT|2712,2715|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2712,2715|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2720,2727|false|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|SIMPLE_SEGMENT|2720,2734|true|false|false|C0007280|Carotid bruit|carotid bruits
Event|Event|SIMPLE_SEGMENT|2728,2734|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|2728,2734|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2737,2742|false|false|false|C0024109|Lung|LUNGS
Finding|Pathologic Function|SIMPLE_SEGMENT|2750,2757|false|false|false|C5441917|Distant Metastasis|distant
Finding|Body Substance|SIMPLE_SEGMENT|2758,2764|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2758,2771|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|2765,2771|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2765,2771|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|2791,2798|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2791,2798|false|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|2804,2812|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2804,2812|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2814,2818|true|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2814,2818|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|SIMPLE_SEGMENT|2819,2828|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|2819,2828|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2833,2849|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|2833,2853|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2843,2849|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2843,2849|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|2850,2853|false|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2850,2853|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2850,2853|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2856,2861|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2856,2861|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|SIMPLE_SEGMENT|2856,2861|false|false|false|||HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|2856,2861|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|SIMPLE_SEGMENT|2864,2867|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2872,2875|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|2872,2875|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2888,2895|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2888,2895|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2888,2895|false|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2898,2902|false|false|false|||NABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2904,2909|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2904,2909|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2911,2915|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2911,2915|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2926,2932|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|2936,2939|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2936,2939|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2945,2952|false|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|2953,2961|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2953,2961|false|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2964,2975|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|2978,2981|false|false|false|||WWP
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2996,3013|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|SIMPLE_SEGMENT|3007,3013|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3007,3013|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3007,3013|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3007,3013|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|3024,3027|false|false|false|||DPs
Finding|Gene or Genome|SIMPLE_SEGMENT|3024,3027|false|false|false|C1843919|PDSS1 gene|DPs
Anatomy|Body System|SIMPLE_SEGMENT|3032,3036|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3032,3036|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|3042,3048|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3042,3048|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|3052,3059|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|3052,3059|true|false|false|C0221198|Lesion|lesions
Event|Event|SIMPLE_SEGMENT|3070,3075|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|3070,3075|false|false|false|C0234422|Awake (finding)|awake
Event|Event|SIMPLE_SEGMENT|3107,3111|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3107,3111|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|3115,3124|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3115,3124|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Anatomy|Cell|SIMPLE_SEGMENT|3141,3144|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3149,3152|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3149,3152|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3149,3152|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3159,3162|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3159,3162|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|3159,3162|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|3159,3162|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3159,3162|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3169,3172|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3169,3172|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|3179,3182|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3179,3182|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3179,3182|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3179,3182|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3179,3182|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3187,3190|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3187,3190|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3187,3190|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3187,3190|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3187,3190|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3187,3190|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3196,3200|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3196,3200|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Finding|Body Substance|SIMPLE_SEGMENT|3241,3247|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|3254,3259|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3254,3259|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|3254,3259|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3264,3267|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|3264,3267|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|3264,3267|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3325,3331|false|false|false|C0023764|lipase|LIPASE
Drug|Enzyme|SIMPLE_SEGMENT|3325,3331|false|false|false|C0023764|lipase|LIPASE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3325,3331|false|false|false|C0023764|lipase|LIPASE
Event|Event|SIMPLE_SEGMENT|3325,3331|false|false|false|||LIPASE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3325,3331|false|false|false|C0373670|Lipase measurement|LIPASE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3349,3352|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3349,3352|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3349,3352|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3349,3352|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3349,3352|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3349,3352|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3349,3352|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3349,3352|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3353,3357|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|3353,3357|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|3353,3357|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|3353,3357|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3353,3357|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3363,3366|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3363,3366|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3363,3366|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3363,3366|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3363,3366|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3363,3366|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3363,3366|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3367,3371|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|3367,3371|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|3367,3371|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|3367,3371|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3367,3371|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3377,3380|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|3377,3380|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|3377,3380|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|3377,3380|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|3377,3380|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3377,3385|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|3377,3385|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3377,3385|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|3381,3385|false|false|false|||PHOS
Event|Event|SIMPLE_SEGMENT|3389,3392|false|false|false|||TOT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3417,3424|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|3417,3424|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3417,3424|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|3417,3424|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3417,3424|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3417,3424|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3430,3434|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|3430,3434|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3430,3434|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|3430,3434|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3430,3434|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3450,3456|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3450,3456|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3450,3456|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|3450,3456|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|3450,3456|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3450,3456|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3462,3471|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3462,3471|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|3462,3471|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3462,3471|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3462,3471|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|3462,3471|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|3462,3471|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3462,3471|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3476,3484|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|3476,3484|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|3476,3484|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3476,3484|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3494,3497|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3494,3497|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|SIMPLE_SEGMENT|3494,3497|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|3494,3497|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3501,3506|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3501,3510|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3501,3510|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3501,3510|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3507,3510|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3507,3510|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|3507,3510|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|3507,3510|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Organic Chemical|SIMPLE_SEGMENT|3528,3535|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3528,3535|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Event|Event|SIMPLE_SEGMENT|3528,3535|false|false|false|||LACTATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3528,3535|false|false|false|C0202115|Lactic acid measurement|LACTATE
Finding|Body Substance|SIMPLE_SEGMENT|3552,3557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3552,3557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3552,3557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|3552,3564|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3559,3564|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3559,3564|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Finding|Idea or Concept|SIMPLE_SEGMENT|3579,3584|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|3604,3609|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3604,3609|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3604,3609|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3604,3616|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3611,3616|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3611,3616|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3611,3616|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|3617,3620|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3617,3620|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3621,3628|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3621,3628|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3621,3628|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|SIMPLE_SEGMENT|3629,3632|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3633,3640|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3633,3640|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|SIMPLE_SEGMENT|3633,3640|false|false|false|||PROTEIN
Finding|Conceptual Entity|SIMPLE_SEGMENT|3633,3640|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3633,3640|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|SIMPLE_SEGMENT|3641,3644|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3641,3644|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3646,3653|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|3646,3653|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3646,3653|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|3646,3653|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3646,3653|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3646,3653|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|SIMPLE_SEGMENT|3654,3657|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3654,3657|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|3658,3664|false|false|false|C0022634|Ketones|KETONE
Event|Event|SIMPLE_SEGMENT|3665,3668|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3665,3668|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3669,3678|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|SIMPLE_SEGMENT|3669,3678|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3669,3678|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3669,3678|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|SIMPLE_SEGMENT|3679,3682|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3679,3682|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3693,3696|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3693,3696|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3705,3709|false|false|false|||LEUK
Event|Event|SIMPLE_SEGMENT|3710,3712|false|false|false|||TR
Finding|Body Substance|SIMPLE_SEGMENT|3725,3730|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3725,3730|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3725,3730|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3725,3735|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|SIMPLE_SEGMENT|3732,3735|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3732,3735|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3732,3735|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|3739,3742|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|3742,3743|false|false|false|||-
Event|Event|SIMPLE_SEGMENT|3745,3753|false|false|false|||BACTERIA
Finding|Functional Concept|SIMPLE_SEGMENT|3745,3753|false|false|false|C1510439|bacteria aspects|BACTERIA
Drug|Food|SIMPLE_SEGMENT|3759,3764|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|3759,3764|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3759,3764|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3759,3764|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|3759,3764|false|false|false|||YEAST
Event|Event|SIMPLE_SEGMENT|3765,3769|false|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3771,3774|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3771,3774|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3771,3774|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|SIMPLE_SEGMENT|3771,3774|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|SIMPLE_SEGMENT|3771,3774|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3771,3774|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|SIMPLE_SEGMENT|3771,3774|false|false|false|||EPI
Finding|Gene or Genome|SIMPLE_SEGMENT|3771,3774|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|SIMPLE_SEGMENT|3771,3774|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3771,3774|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|SIMPLE_SEGMENT|3789,3794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3789,3794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3789,3794|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|3789,3802|false|false|false|C0455910|Mucus in urine (finding)|URINE  MUCOUS
Finding|Body Substance|SIMPLE_SEGMENT|3796,3802|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|MUCOUS
Event|Event|SIMPLE_SEGMENT|3803,3807|false|false|false|||RARE
Finding|Gene or Genome|SIMPLE_SEGMENT|3803,3807|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Event|Event|SIMPLE_SEGMENT|3809,3816|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|3809,3816|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3809,3816|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|SIMPLE_SEGMENT|3819,3822|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3819,3822|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|3828,3838|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|3828,3838|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|3828,3838|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|3841,3845|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Event|Event|SIMPLE_SEGMENT|3856,3866|false|false|false|||prominence
Event|Event|SIMPLE_SEGMENT|3868,3877|false|false|false|||suspected
Event|Activity|SIMPLE_SEGMENT|3881,3890|false|false|false|C1882932|Representation (action)|represent
Event|Event|SIMPLE_SEGMENT|3881,3890|false|false|false|||represent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3909,3918|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3909,3918|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3909,3918|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3909,3926|false|false|false|C1508661|Pulmonary vessels|pulmonary vessels
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3919,3926|false|false|false|C0005847|Blood Vessel|vessels
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3944,3953|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|3944,3953|false|false|false|||pneumonia
Finding|Functional Concept|SIMPLE_SEGMENT|3965,3969|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|3978,3991|false|false|false|||opacification
Event|Event|SIMPLE_SEGMENT|3992,3996|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|4026,4034|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|SIMPLE_SEGMENT|4026,4034|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4042,4047|false|false|false|C1446899|minor (disease)|minor
Event|Event|SIMPLE_SEGMENT|4042,4047|false|false|false|||minor
Finding|Gene or Genome|SIMPLE_SEGMENT|4042,4047|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Event|Event|SIMPLE_SEGMENT|4048,4059|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4048,4059|false|false|false|C0004144|Atelectasis|atelectasis
Event|Event|SIMPLE_SEGMENT|4063,4071|false|false|false|||scarring
Finding|Pathologic Function|SIMPLE_SEGMENT|4063,4071|false|false|false|C0008767;C2004491|Cicatrix;Cicatrization|scarring
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4078,4082|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Drug|Enzyme|SIMPLE_SEGMENT|4078,4082|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Event|Event|SIMPLE_SEGMENT|4081,4082|false|false|false|||A
Finding|Intellectual Product|SIMPLE_SEGMENT|4098,4103|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Functional Concept|SIMPLE_SEGMENT|4104,4119|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Event|Event|SIMPLE_SEGMENT|4120,4129|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|4120,4129|true|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|4120,4129|true|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4120,4129|true|false|false|C0919386|Pathology procedure|pathology
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4140,4154|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|SIMPLE_SEGMENT|4140,4154|false|false|false|||diverticulosis
Event|Event|SIMPLE_SEGMENT|4160,4168|false|false|false|||sequelae
Finding|Pathologic Function|SIMPLE_SEGMENT|4160,4168|false|false|false|C0243088;C0543419|Sequela of disorder;sequelae aspects|sequelae
Event|Event|SIMPLE_SEGMENT|4178,4190|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|4178,4190|false|false|false|C0021368|Inflammation|inflammation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4207,4221|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|4207,4221|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|4240,4244|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|4255,4260|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4255,4274|false|false|false|C0929209|Right major fissure|right major fissure
Finding|Classification|SIMPLE_SEGMENT|4261,4266|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|major
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4261,4274|false|false|false|C0929208|Major fissure|major fissure
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4267,4274|false|false|false|C0332469|Fissure|fissure
Event|Event|SIMPLE_SEGMENT|4279,4284|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|4279,4284|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4286,4291|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4286,4291|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4286,4296|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4292,4296|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4292,4296|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|4316,4326|false|false|false|||guidelines
Finding|Intellectual Product|SIMPLE_SEGMENT|4316,4326|false|false|false|C0162791;C0220845;C0282423|Guideline (Publication Type);Guidelines;guiding characteristics|guidelines
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4335,4342|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|SIMPLE_SEGMENT|4335,4342|false|false|false|||absence
Finding|Functional Concept|SIMPLE_SEGMENT|4335,4342|false|false|false|C0332197|Absent|absence
Finding|Idea or Concept|SIMPLE_SEGMENT|4347,4351|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4347,4359|false|false|false|C1830376||risk factors
Finding|Finding|SIMPLE_SEGMENT|4347,4359|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|SIMPLE_SEGMENT|4347,4359|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|SIMPLE_SEGMENT|4352,4359|false|false|false|||factors
Event|Event|SIMPLE_SEGMENT|4372,4380|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|4372,4380|true|false|true|C1522577|follow-up|followup
Event|Event|SIMPLE_SEGMENT|4384,4390|false|false|false|||needed
Finding|Body Substance|SIMPLE_SEGMENT|4396,4403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4396,4403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4396,4403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|4396,4407|false|false|false|C0332310|Has patient|patient has
Finding|Idea or Concept|SIMPLE_SEGMENT|4409,4413|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4409,4421|false|false|false|C1830376||risk factors
Finding|Finding|SIMPLE_SEGMENT|4409,4421|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|SIMPLE_SEGMENT|4409,4421|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|SIMPLE_SEGMENT|4414,4421|false|false|false|||factors
Event|Event|SIMPLE_SEGMENT|4430,4437|false|false|false|||smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|4430,4437|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|4430,4437|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Event|Event|SIMPLE_SEGMENT|4439,4447|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|4439,4447|false|false|false|C1522577|follow-up|followup
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4448,4453|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|4448,4453|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4448,4456|false|false|false|C0202823|Chest CT|chest CT
Event|Event|SIMPLE_SEGMENT|4454,4456|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|4474,4485|false|false|false|||recommended
Finding|Intellectual Product|SIMPLE_SEGMENT|4489,4497|false|false|false|C1301746;C1547673;C1563337|ActClass - document;Document type;Documents|document
Event|Event|SIMPLE_SEGMENT|4498,4507|false|false|false|||stability
Event|Event|SIMPLE_SEGMENT|4511,4514|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4511,4514|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|SIMPLE_SEGMENT|4530,4533|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|4530,4533|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4534,4538|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4534,4538|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4534,4538|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4534,4538|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4534,4546|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|SIMPLE_SEGMENT|4539,4546|false|false|false|||volumes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4555,4565|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|4555,4565|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|4555,4565|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Event|SIMPLE_SEGMENT|4586,4594|false|false|false|||crowding
Finding|Finding|SIMPLE_SEGMENT|4586,4594|false|false|false|C0010383;C0040433|Crowding;Tooth Crowding|crowding
Finding|Social Behavior|SIMPLE_SEGMENT|4586,4594|false|false|false|C0010383;C0040433|Crowding;Tooth Crowding|crowding
Finding|Finding|SIMPLE_SEGMENT|4620,4626|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4620,4626|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Intellectual Product|SIMPLE_SEGMENT|4627,4631|false|true|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4632,4640|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|SIMPLE_SEGMENT|4642,4652|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|4642,4652|false|false|false|C0700148|Congestion|congestion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4657,4662|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4657,4662|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4657,4662|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4674,4687|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4674,4687|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|4691,4695|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|4719,4730|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4719,4730|false|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4737,4742|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4737,4742|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|4737,4742|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4737,4742|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|4750,4756|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4771,4777|false|false|false|C0003483|Aorta|aortic
Event|Event|SIMPLE_SEGMENT|4778,4787|false|false|false|||totuosity
Event|Event|SIMPLE_SEGMENT|4794,4804|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4794,4804|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4794,4804|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4807,4811|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4812,4821|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4812,4821|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|4812,4821|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|4812,4827|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4822,4827|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4822,4827|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4822,4827|false|false|false|C0013604|Edema|edema
Finding|Body Substance|SIMPLE_SEGMENT|4832,4837|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|4832,4837|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|4832,4837|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|SIMPLE_SEGMENT|4849,4857|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|4849,4857|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|4849,4857|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4849,4857|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|4860,4864|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4860,4864|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|4868,4877|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4868,4877|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4868,4877|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4868,4877|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4868,4877|false|false|false|C0030685|Patient Discharge|Discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4893,4898|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4893,4898|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4893,4898|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4899,4902|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4909,4912|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4909,4912|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4909,4912|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4919,4922|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4919,4922|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4919,4922|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4919,4922|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4928,4931|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4928,4931|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4939,4942|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4939,4942|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4939,4942|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4939,4942|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4939,4942|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4946,4949|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4946,4949|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4946,4949|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4946,4949|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4946,4949|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4946,4949|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4955,4959|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4955,4959|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|4965,4968|false|false|false|||RDW
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4975,4978|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4995,5000|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4995,5000|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4995,5000|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5005,5008|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|5005,5008|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5005,5008|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5030,5035|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5030,5035|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5030,5035|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5030,5043|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5030,5043|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5030,5043|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5036,5043|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5036,5043|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5036,5043|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5036,5043|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5036,5043|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5036,5043|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5088,5092|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5088,5092|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5088,5092|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5117,5122|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5117,5122|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5117,5122|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5123,5126|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5123,5126|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5123,5126|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|5123,5126|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5123,5126|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5123,5126|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5123,5126|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5123,5126|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5131,5134|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5131,5134|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5131,5134|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5131,5134|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5131,5134|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|5131,5134|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5131,5134|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5139,5146|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5139,5146|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5174,5179|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5174,5179|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5174,5179|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5174,5187|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5180,5187|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5180,5187|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5180,5187|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5180,5187|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5180,5187|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5180,5187|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5180,5187|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5180,5187|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Body Substance|SIMPLE_SEGMENT|5221,5226|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5221,5226|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5221,5226|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5221,5232|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5227,5232|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5227,5232|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Finding|Idea or Concept|SIMPLE_SEGMENT|5247,5252|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|5272,5277|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5272,5277|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5272,5277|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5272,5283|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5278,5283|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|5278,5283|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|SIMPLE_SEGMENT|5284,5287|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5284,5287|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5288,5295|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5288,5295|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5288,5295|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|SIMPLE_SEGMENT|5296,5299|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5296,5299|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5300,5307|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5300,5307|false|false|false|C0033684|Proteins|Protein
Event|Event|SIMPLE_SEGMENT|5300,5307|false|false|false|||Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|5300,5307|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5300,5307|false|false|false|C0202202|Protein measurement|Protein
Event|Event|SIMPLE_SEGMENT|5308,5311|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5308,5311|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5313,5320|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5313,5320|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5313,5320|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5313,5320|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5313,5320|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5313,5320|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|5321,5324|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5321,5324|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|5325,5331|false|false|false|C0022634|Ketones|Ketone
Event|Event|SIMPLE_SEGMENT|5332,5335|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5332,5335|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5344,5347|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5356,5359|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|5388,5393|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5388,5393|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5388,5393|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5388,5397|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|SIMPLE_SEGMENT|5394,5397|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5394,5397|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5394,5397|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|5401,5404|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|SIMPLE_SEGMENT|5420,5425|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|5420,5425|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5420,5425|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5420,5425|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|SIMPLE_SEGMENT|5420,5425|false|false|false|||Yeast
Event|Event|SIMPLE_SEGMENT|5426,5430|false|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5432,5435|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5432,5435|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5432,5435|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|5432,5435|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|5432,5435|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5432,5435|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|SIMPLE_SEGMENT|5432,5435|false|false|false|||Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|5432,5435|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|5432,5435|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5432,5435|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5445,5453|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|5445,5453|false|false|false|||diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5455,5469|false|false|false|C0028756|Morbid obesity|morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5462,5469|false|false|false|C0028754|Obesity|obesity
Event|Event|SIMPLE_SEGMENT|5462,5469|false|false|false|||obesity
Finding|Finding|SIMPLE_SEGMENT|5462,5469|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5479,5482|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|5479,5482|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|5487,5495|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|5512,5518|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|5512,5518|false|false|false|C0015967|Fever|fevers
Drug|Organic Chemical|SIMPLE_SEGMENT|5523,5528|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5523,5528|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|5523,5528|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5523,5528|false|false|false|C0010200|Coughing|cough
Finding|Finding|SIMPLE_SEGMENT|5523,5539|false|false|false|C0239134|Productive Cough|cough productive
Event|Event|SIMPLE_SEGMENT|5529,5539|false|false|false|||productive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5543,5547|false|false|false|C1321554|Bacterial shell rot|rust
Event|Event|SIMPLE_SEGMENT|5543,5547|false|false|false|||rust
Event|Event|SIMPLE_SEGMENT|5556,5562|false|false|false|||sputum
Finding|Body Substance|SIMPLE_SEGMENT|5556,5562|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|5556,5562|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|5580,5583|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|5580,5583|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|5593,5599|false|false|false|||Fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|5593,5599|false|false|false|C0015967|Fever|Fevers
Finding|Finding|SIMPLE_SEGMENT|5601,5607|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5601,5607|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5608,5617|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|5608,5617|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|5608,5617|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5621,5630|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|5621,5630|false|false|false|||pneumonia
Finding|Finding|SIMPLE_SEGMENT|5636,5644|false|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|5647,5652|false|false|false|||viral
Finding|Functional Concept|SIMPLE_SEGMENT|5647,5652|false|false|false|C0521026|Viral|viral
Event|Event|SIMPLE_SEGMENT|5654,5661|false|false|false|||illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|5654,5661|false|false|false|C0221423|Illness (finding)|illness
Finding|Idea or Concept|SIMPLE_SEGMENT|5663,5674|false|false|false|C0750501|most likely|Most likely
Finding|Finding|SIMPLE_SEGMENT|5668,5674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5668,5674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5679,5696|true|true|false|C2350512|Bacterial Processes|bacterial process
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5689,5696|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5689,5696|false|true|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|5689,5696|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|5689,5696|false|true|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5689,5696|false|true|false|C1522240|Process|process
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5704,5716|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|5704,5716|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|5704,5716|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|5724,5727|false|false|false|||PMN
Finding|Cell Function|SIMPLE_SEGMENT|5724,5727|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Finding|Intellectual Product|SIMPLE_SEGMENT|5724,5727|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Event|Event|SIMPLE_SEGMENT|5728,5740|false|false|false|||predominance
Finding|Body Substance|SIMPLE_SEGMENT|5742,5747|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|5742,5747|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|5742,5747|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|SIMPLE_SEGMENT|5748,5758|false|false|false|||legionella
Finding|Finding|SIMPLE_SEGMENT|5759,5762|false|false|false|C5848551|Neg - answer|neg
Event|Event|SIMPLE_SEGMENT|5764,5767|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5764,5767|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|5807,5811|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|5815,5821|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|5815,5821|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|5815,5821|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Intellectual Product|SIMPLE_SEGMENT|5826,5833|false|false|false|C0282416|Overall Publication Type|overall
Event|Event|SIMPLE_SEGMENT|5834,5847|false|false|false|||constellation
Event|Event|SIMPLE_SEGMENT|5852,5860|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|5852,5860|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|5852,5860|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|5886,5892|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|5886,5892|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|5886,5892|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|5886,5892|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Finding|SIMPLE_SEGMENT|5897,5900|false|false|false|C5848551|Neg - answer|neg
Event|Event|SIMPLE_SEGMENT|5901,5903|false|false|false|||CT
Finding|Body Substance|SIMPLE_SEGMENT|5909,5916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5909,5916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5909,5916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5921,5928|false|false|false|||treated
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5947,5950|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5947,5950|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|5947,5950|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|5947,5950|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5947,5950|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|SIMPLE_SEGMENT|5956,5960|false|false|false|||sats
Event|Event|SIMPLE_SEGMENT|5961,5967|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|5961,5967|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5972,5980|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5977,5980|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5977,5980|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|5977,5980|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|5977,5980|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|5977,5980|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|5977,5980|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|5977,5980|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Idea or Concept|SIMPLE_SEGMENT|5992,5995|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5992,5995|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|6010,6019|false|false|false|||de-satted
Event|Event|SIMPLE_SEGMENT|6025,6029|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|6025,6029|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|6025,6029|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6031,6036|false|false|false|C0024109|Lung|lungs
Finding|Finding|SIMPLE_SEGMENT|6043,6051|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|6043,6051|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|SIMPLE_SEGMENT|6052,6060|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|6052,6060|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|6083,6093|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6083,6093|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|6083,6093|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|6111,6117|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|6118,6121|false|false|false|||cxr
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6118,6121|false|false|false|C0039985|Plain chest X-ray|cxr
Procedure|Health Care Activity|SIMPLE_SEGMENT|6127,6131|false|false|false|C1315068|Pulmonary ventilator management|pulm
Finding|Pathologic Function|SIMPLE_SEGMENT|6127,6137|false|false|false|C0034063|Pulmonary Edema|pulm edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6132,6137|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6132,6137|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6132,6137|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|6138,6144|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6138,6144|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Substance|SIMPLE_SEGMENT|6152,6160|false|true|false|C1289919|Intravenous fluid|IV fluid
Drug|Substance|SIMPLE_SEGMENT|6155,6160|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6155,6160|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6155,6160|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|6161,6166|false|false|false|||bolus
Finding|Body Substance|SIMPLE_SEGMENT|6161,6166|false|true|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|SIMPLE_SEGMENT|6161,6166|false|true|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6161,6166|false|true|false|C1511237|bolus infusion|bolus
Finding|Idea or Concept|SIMPLE_SEGMENT|6168,6171|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6168,6171|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|6193,6198|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6193,6198|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|6204,6208|false|false|false|||POx1
Event|Event|SIMPLE_SEGMENT|6214,6217|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|6214,6217|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6214,6217|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6226,6230|false|false|false|C0312448|short-acting thyroid stimulator|sats
Drug|Hormone|SIMPLE_SEGMENT|6226,6230|false|false|false|C0312448|short-acting thyroid stimulator|sats
Event|Event|SIMPLE_SEGMENT|6226,6230|false|false|false|||sats
Event|Event|SIMPLE_SEGMENT|6274,6284|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6274,6284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|6274,6284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|SIMPLE_SEGMENT|6308,6311|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|6308,6311|false|false|false|C0013404|Dyspnea|SOB
Finding|Finding|SIMPLE_SEGMENT|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6328,6336|false|true|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|6328,6336|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6328,6336|false|true|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|6348,6355|false|false|false|||habitus
Event|Event|SIMPLE_SEGMENT|6359,6366|false|false|false|||Treated
Drug|Organic Chemical|SIMPLE_SEGMENT|6372,6381|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6372,6381|false|false|false|C0001927|albuterol|albuterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6382,6386|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|6382,6386|false|false|false|||nebs
Drug|Antibiotic|SIMPLE_SEGMENT|6391,6403|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|6391,6403|false|false|false|C0282386|levofloxacin|Levofloxacin
Event|Event|SIMPLE_SEGMENT|6404,6409|false|false|false|||750mg
Drug|Organic Chemical|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6435,6443|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|6435,6443|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|6435,6443|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6435,6443|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6446,6449|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6446,6449|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|6450,6456|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|6460,6472|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|6460,6472|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|6460,6472|false|false|false|||levofloxacin
Event|Event|SIMPLE_SEGMENT|6513,6522|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6513,6522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6513,6522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6513,6522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6513,6522|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|6524,6532|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|6524,6532|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|6524,6532|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Body Substance|SIMPLE_SEGMENT|6565,6570|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|6565,6570|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|6565,6570|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|6571,6576|false|false|false|||lytes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6577,6580|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6577,6580|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6577,6580|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Event|Event|SIMPLE_SEGMENT|6577,6580|false|false|false|||osm
Finding|Gene or Genome|SIMPLE_SEGMENT|6577,6580|false|false|false|C1335093;C1427709|CCM2 gene;OSM gene|osm
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6585,6590|false|false|false|C5575602|Cell Culture Serum|serum
Event|Event|SIMPLE_SEGMENT|6585,6590|false|false|false|||serum
Finding|Body Substance|SIMPLE_SEGMENT|6585,6590|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|6585,6590|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6591,6594|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6591,6594|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6591,6594|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Event|Event|SIMPLE_SEGMENT|6591,6594|false|false|false|||osm
Finding|Gene or Genome|SIMPLE_SEGMENT|6591,6594|false|false|false|C1335093;C1427709|CCM2 gene;OSM gene|osm
Finding|Idea or Concept|SIMPLE_SEGMENT|6596,6607|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|6601,6607|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6601,6607|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6609,6614|false|false|false|C0021141|Inappropriate ADH Syndrome|SIADH
Event|Event|SIMPLE_SEGMENT|6609,6614|false|false|false|||SIADH
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6615,6624|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|6615,6624|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6615,6624|false|false|false|C1522484|metastatic qualifier|secondary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6628,6637|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6628,6637|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6628,6637|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6628,6645|false|false|false|C0748169|PULMONARY PROCESS|pulmonary process
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6638,6645|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6638,6645|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|6638,6645|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|6638,6645|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6638,6645|false|false|false|C1522240|Process|process
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6651,6659|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|6651,6659|false|false|false|||Diabetes
Event|Event|SIMPLE_SEGMENT|6661,6667|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6661,6667|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|SIMPLE_SEGMENT|6670,6679|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6680,6684|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6680,6684|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6680,6684|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6685,6691|false|false|false|C0876064|Lantus|Lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6685,6691|false|false|false|C0876064|Lantus|Lantus
Event|Event|SIMPLE_SEGMENT|6685,6691|false|false|false|||Lantus
Event|Event|SIMPLE_SEGMENT|6705,6708|false|false|false|||ISS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6712,6716|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6712,6716|false|false|false|C0675390|ARID1A protein, human|Held
Finding|Gene or Genome|SIMPLE_SEGMENT|6712,6716|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|SIMPLE_SEGMENT|6712,6716|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Drug|Organic Chemical|SIMPLE_SEGMENT|6717,6726|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6717,6726|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|6717,6726|false|false|false|||metformin
Event|Event|SIMPLE_SEGMENT|6738,6741|false|false|false|||Was
Finding|Finding|SIMPLE_SEGMENT|6745,6753|false|false|false|C0241863|Diabetic|diabetic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6745,6758|false|false|false|C0011878|Diabetic Diet|diabetic diet
Drug|Food|SIMPLE_SEGMENT|6754,6758|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|6754,6758|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|6754,6758|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|6754,6758|false|false|false|C0012159|Diet therapy|diet
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6768,6771|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6768,6771|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6773,6782|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6783,6787|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6783,6787|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6783,6787|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6788,6798|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6788,6798|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|6788,6798|false|false|false|||lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|6800,6810|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6800,6810|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|6800,6810|false|false|false|||metoprolol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6813,6817|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6813,6817|false|false|false|C0675390|ARID1A protein, human|Held
Finding|Gene or Genome|SIMPLE_SEGMENT|6813,6817|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|SIMPLE_SEGMENT|6813,6817|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Drug|Organic Chemical|SIMPLE_SEGMENT|6818,6823|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6818,6823|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|6818,6823|false|false|false|||lasix
Finding|Mental Process|SIMPLE_SEGMENT|6838,6845|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6849,6860|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6849,6860|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|SIMPLE_SEGMENT|6849,6860|false|false|false|||dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6849,6860|false|false|false|C4284399|Dehydration procedure|dehydration
Event|Event|SIMPLE_SEGMENT|6873,6883|false|false|false|||Re-started
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6901,6904|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6901,6904|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6901,6904|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6901,6904|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6901,6904|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6901,6904|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6901,6904|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6901,6904|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6917,6920|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|6917,6920|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6917,6920|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|6917,6920|false|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|6917,6920|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6917,6920|false|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|6921,6926|false|false|false|||shows
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6932,6935|false|false|false|C0036916|Sexually Transmitted Diseases|STD
Drug|Organic Chemical|SIMPLE_SEGMENT|6932,6935|false|false|false|C0592138|STD brand of sodium tetradecyl sulfate|STD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6932,6935|false|false|false|C0592138|STD brand of sodium tetradecyl sulfate|STD
Event|Event|SIMPLE_SEGMENT|6932,6935|false|false|false|||STD
Finding|Gene or Genome|SIMPLE_SEGMENT|6932,6935|false|false|false|C1420519;C1421567;C1705831|SULT2A1 gene;ZAP70 gene;ZAP70 wt Allele|STD
Event|Event|SIMPLE_SEGMENT|6959,6968|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6969,6973|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6969,6973|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6969,6973|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6974,6977|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Enzyme|SIMPLE_SEGMENT|6974,6977|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Organic Chemical|SIMPLE_SEGMENT|6974,6977|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6974,6977|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Event|Event|SIMPLE_SEGMENT|6974,6977|false|false|false|||asa
Finding|Gene or Genome|SIMPLE_SEGMENT|6974,6977|false|false|false|C1412553|ARSA gene|asa
Drug|Organic Chemical|SIMPLE_SEGMENT|6979,6989|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6979,6989|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|6979,6989|false|false|false|||metoprolol
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6991,6996|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6991,6996|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6991,6996|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|6997,7009|false|false|false|C0452415|Diet, Healthy|healthy diet
Drug|Food|SIMPLE_SEGMENT|7005,7009|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|7005,7009|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|7005,7009|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|7005,7009|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|7022,7028|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|7022,7028|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|SIMPLE_SEGMENT|7031,7040|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7041,7045|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7041,7045|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7041,7045|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7046,7057|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7046,7057|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|SIMPLE_SEGMENT|7046,7057|false|false|false|||simvastatin
Event|Event|SIMPLE_SEGMENT|7058,7065|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|7058,7065|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|7066,7069|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|SIMPLE_SEGMENT|7066,7069|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|SIMPLE_SEGMENT|7066,7069|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7070,7073|false|false|false|C2606415|ZDHHC2 protein, human|rec
Drug|Enzyme|SIMPLE_SEGMENT|7070,7073|false|false|false|C2606415|ZDHHC2 protein, human|rec
Event|Event|SIMPLE_SEGMENT|7070,7073|false|false|false|||rec
Finding|Gene or Genome|SIMPLE_SEGMENT|7070,7073|false|false|false|C1422148;C1424025|MCM8 gene;RBPJP4 gene|rec
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7095,7102|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|SIMPLE_SEGMENT|7095,7102|false|false|false|||Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|7095,7102|false|false|false|C0860603|Anxiety symptoms|Anxiety
Event|Event|SIMPLE_SEGMENT|7104,7110|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|7104,7110|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|SIMPLE_SEGMENT|7113,7122|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7123,7127|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7128,7137|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7128,7137|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|SIMPLE_SEGMENT|7128,7137|false|false|false|||lorazepam
Drug|Organic Chemical|SIMPLE_SEGMENT|7139,7151|false|false|false|C1099456|escitalopram|escitalopram
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7139,7151|false|false|false|C1099456|escitalopram|escitalopram
Event|Event|SIMPLE_SEGMENT|7139,7151|false|false|false|||escitalopram
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7161,7167|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|7161,7167|false|false|false|||Anemia
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7169,7172|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7169,7172|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7180,7188|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|7180,7188|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7180,7188|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7202,7206|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|7202,7206|false|false|false|||GERD
Event|Event|SIMPLE_SEGMENT|7208,7214|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|7208,7214|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Drug|Organic Chemical|SIMPLE_SEGMENT|7229,7239|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7229,7239|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|SIMPLE_SEGMENT|7229,7239|false|false|false|||omeprazole
Finding|Idea or Concept|SIMPLE_SEGMENT|7244,7248|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7244,7248|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7244,7248|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7249,7261|false|false|false|C0937846|esomeprazole|esomeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7249,7261|false|false|false|C0937846|esomeprazole|esomeprazole
Event|Event|SIMPLE_SEGMENT|7249,7261|false|false|false|||esomeprazole
Finding|Functional Concept|SIMPLE_SEGMENT|7266,7276|false|false|false|C0444507|Incidental|incidental
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7277,7289|false|false|false|C0444708|Radiographic|radiographic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7290,7298|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|7290,7298|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|7290,7298|false|false|false|C2607943|findings aspects|findings
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7299,7308|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7299,7308|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7299,7308|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|7299,7315|false|false|false|C0034079||pulmonary nodule
Event|Event|SIMPLE_SEGMENT|7309,7315|false|false|false|||nodule
Event|Event|SIMPLE_SEGMENT|7322,7329|false|false|false|||require
Event|Event|SIMPLE_SEGMENT|7331,7337|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|7348,7359|false|false|false|||TRANSITIONS
Event|Activity|SIMPLE_SEGMENT|7363,7367|false|false|false|C1947933|care activity|CARE
Event|Event|SIMPLE_SEGMENT|7363,7367|false|false|false|||CARE
Finding|Finding|SIMPLE_SEGMENT|7363,7367|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|7363,7367|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Drug|Organic Chemical|SIMPLE_SEGMENT|7376,7384|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7376,7384|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7376,7384|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7376,7384|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7376,7384|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7376,7384|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7385,7388|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7385,7388|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|7385,7390|false|false|false|C3842674|Day 5|day 5
Event|Event|SIMPLE_SEGMENT|7389,7390|false|false|false|||5
Drug|Antibiotic|SIMPLE_SEGMENT|7394,7406|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|7394,7406|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|7407,7413|false|false|false|||course
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7433,7437|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|7438,7445|false|false|false|||checked
Event|Event|SIMPLE_SEGMENT|7468,7473|false|false|false|||faxed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7477,7480|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7477,7480|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7477,7480|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7477,7480|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|7477,7480|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7477,7480|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|7477,7480|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7477,7480|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|7477,7480|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|7477,7480|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|7477,7480|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|7497,7498|false|false|false|||f
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7506,7509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7506,7509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7506,7509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7506,7509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|7506,7509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7506,7509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|7506,7509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7506,7509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|7506,7509|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|7506,7509|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|7506,7509|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|SIMPLE_SEGMENT|7510,7514|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|SIMPLE_SEGMENT|7515,7519|false|false|false|||week
Finding|Intellectual Product|SIMPLE_SEGMENT|7515,7519|false|false|false|C1561540|Transaction counts and value totals - week|week
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7526,7530|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7526,7530|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7526,7530|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|7526,7530|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|7526,7537|false|false|false|C0034079||lung nodule
Event|Event|SIMPLE_SEGMENT|7531,7537|false|false|false|||nodule
Event|Event|SIMPLE_SEGMENT|7538,7542|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|7546,7549|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7546,7549|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|7558,7566|false|false|false|||followed
Event|Event|SIMPLE_SEGMENT|7578,7582|false|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|7578,7582|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|7578,7582|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Finding|Finding|SIMPLE_SEGMENT|7584,7593|false|false|false|C0750484|Confirmation|Confirmed
Event|Activity|SIMPLE_SEGMENT|7603,7610|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|7603,7610|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|7603,7610|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|7603,7610|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|7603,7610|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7603,7610|false|false|false|C0392367|Physical contact|CONTACT
Procedure|Health Care Activity|SIMPLE_SEGMENT|7640,7649|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7651,7658|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7651,7658|false|false|false|C0528249|Humalog|Humalog
Drug|Organic Chemical|SIMPLE_SEGMENT|7665,7670|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7665,7670|false|false|false|C0699992|Lasix|Lasix
Drug|Organic Chemical|SIMPLE_SEGMENT|7684,7695|false|false|false|C0012125|dicyclomine|Dicyclomine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7684,7695|false|false|false|C0012125|dicyclomine|Dicyclomine
Finding|Gene or Genome|SIMPLE_SEGMENT|7707,7710|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7713,7726|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7713,7726|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7713,7726|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7713,7726|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7741,7753|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7741,7753|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Organic Chemical|SIMPLE_SEGMENT|7767,7777|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7767,7777|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|7767,7787|false|false|false|C0724633|metoprolol succinate|Metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7767,7787|false|false|false|C0724633|metoprolol succinate|Metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|7778,7787|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7801,7807|false|false|false|C0876064|Lantus|Lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7801,7807|false|false|false|C0876064|Lantus|Lantus
Event|Event|SIMPLE_SEGMENT|7801,7807|false|false|false|||Lantus
Event|Event|SIMPLE_SEGMENT|7817,7820|false|false|false|||QHS
Drug|Organic Chemical|SIMPLE_SEGMENT|7823,7830|false|false|false|C0483514|Vicodin|Vicodin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7823,7830|false|false|false|C0483514|Vicodin|Vicodin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7833,7836|false|false|false|C0039225|Tablet Dosage Form|tab
Finding|Gene or Genome|SIMPLE_SEGMENT|7843,7846|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|7849,7858|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7849,7858|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|SIMPLE_SEGMENT|7863,7866|false|false|false|||QHS
Finding|Gene or Genome|SIMPLE_SEGMENT|7867,7870|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|7873,7885|false|false|false|C0937846|esomeprazole|Esomeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7873,7885|false|false|false|C0937846|esomeprazole|Esomeprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7891,7894|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7891,7894|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7891,7894|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7891,7894|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7891,7894|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7897,7907|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7897,7907|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|7921,7932|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7921,7932|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|7944,7953|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7944,7953|false|false|false|C0025598|metformin|Metformin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7961,7964|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7961,7964|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7961,7964|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7961,7964|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7961,7964|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7967,7974|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7967,7982|false|false|false|C0060282|ferrous sulfate|Ferrous sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7967,7982|false|false|false|C0060282|ferrous sulfate|Ferrous sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7975,7982|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7975,7982|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7975,7982|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|7989,7992|false|false|false|||TID
Event|Event|SIMPLE_SEGMENT|7998,8007|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7998,8007|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7998,8019|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8008,8019|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8008,8019|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8008,8019|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8008,8019|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8024,8036|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8024,8036|false|false|false|C1099456|escitalopram|Escitalopram
Event|Event|SIMPLE_SEGMENT|8024,8036|false|false|false|||Escitalopram
Drug|Organic Chemical|SIMPLE_SEGMENT|8024,8044|false|false|false|C1170746|escitalopram oxalate|Escitalopram Oxalate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8024,8044|false|false|false|C1170746|escitalopram oxalate|Escitalopram Oxalate
Drug|Organic Chemical|SIMPLE_SEGMENT|8037,8044|false|false|false|C0029988;C3669135|Oxalates;oxalate|Oxalate
Event|Event|SIMPLE_SEGMENT|8037,8044|false|false|false|||Oxalate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8037,8044|false|false|false|C0202153|Oxalate measurement|Oxalate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8064,8074|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8064,8074|false|false|false|C0065374|lisinopril|Lisinopril
Event|Activity|SIMPLE_SEGMENT|8091,8095|false|false|false|C1948035|Hold (action)|hold
Event|Event|SIMPLE_SEGMENT|8091,8095|false|false|false|||hold
Finding|Functional Concept|SIMPLE_SEGMENT|8091,8095|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|SIMPLE_SEGMENT|8091,8095|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8100,8103|false|false|false|C0871470|Systolic Pressure|sbp
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8100,8103|false|false|false|C0085805|Androgen Binding Protein|sbp
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8100,8103|false|false|false|C0085805|Androgen Binding Protein|sbp
Event|Event|SIMPLE_SEGMENT|8100,8103|false|false|false|||sbp
Finding|Gene or Genome|SIMPLE_SEGMENT|8100,8103|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|sbp
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8100,8103|false|false|false|C1306620|Systolic blood pressure measurement|sbp
Drug|Organic Chemical|SIMPLE_SEGMENT|8112,8124|false|false|false|C0937846|esomeprazole|esomeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8112,8124|false|false|false|C0937846|esomeprazole|esomeprazole
Event|Event|SIMPLE_SEGMENT|8112,8124|false|false|false|||esomeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|8112,8134|false|false|false|C0937622|esomeprazole magnesium|esomeprazole magnesium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8112,8134|false|false|false|C0937622|esomeprazole magnesium|esomeprazole magnesium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8125,8134|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8125,8134|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8125,8134|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8125,8134|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Event|Event|SIMPLE_SEGMENT|8125,8134|false|false|false|||magnesium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8125,8134|false|false|false|C0373675|Magnesium measurement|magnesium
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8146,8150|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8146,8150|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|8146,8150|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|8146,8150|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8151,8154|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8151,8154|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8151,8154|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8151,8154|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8151,8154|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8159,8166|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8159,8174|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8159,8174|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8167,8174|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8167,8174|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8167,8174|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|SIMPLE_SEGMENT|8167,8174|false|false|false|||Sulfate
Event|Event|SIMPLE_SEGMENT|8185,8188|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|8193,8204|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8193,8204|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Finding|Gene or Genome|SIMPLE_SEGMENT|8218,8221|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8222,8226|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8222,8226|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8222,8226|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8222,8226|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8231,8244|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|8231,8244|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|8231,8244|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8231,8244|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8231,8251|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|8231,8251|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8231,8251|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8245,8251|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8245,8251|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8245,8251|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|8245,8251|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8245,8251|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8245,8251|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|8272,8282|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8272,8282|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8272,8292|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8272,8292|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|8283,8292|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|8283,8292|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|8315,8324|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8315,8324|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|8336,8339|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8340,8348|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|SIMPLE_SEGMENT|8340,8348|false|false|false|||insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|8340,8348|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8353,8361|false|false|false|C0907402|insulin glargine|Glargine
Drug|Hormone|SIMPLE_SEGMENT|8353,8361|false|false|false|C0907402|insulin glargine|Glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8353,8361|false|false|false|C0907402|insulin glargine|Glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8380,8387|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|8380,8387|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8380,8387|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|8380,8387|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8380,8387|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8380,8387|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|8391,8398|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|8391,8398|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8391,8404|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8399,8404|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|8399,8404|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|8399,8404|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|8399,8404|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Event|Event|SIMPLE_SEGMENT|8431,8439|false|false|false|||Override
Finding|Functional Concept|SIMPLE_SEGMENT|8431,8439|false|false|false|C1547671|Override|Override
Event|Event|SIMPLE_SEGMENT|8441,8447|false|false|false|||Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|8441,8447|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|8449,8453|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8449,8453|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8449,8453|false|false|false|C1553498|home health encounter|home
Drug|Antibiotic|SIMPLE_SEGMENT|8466,8478|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|8466,8478|false|false|false|C0282386|levofloxacin|Levofloxacin
Event|Event|SIMPLE_SEGMENT|8495,8500|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|8514,8517|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8514,8517|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Antibiotic|SIMPLE_SEGMENT|8530,8542|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|8530,8542|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|8530,8542|false|false|false|||levofloxacin
Finding|Intellectual Product|SIMPLE_SEGMENT|8550,8554|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8550,8560|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|8557,8560|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8557,8560|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8570,8576|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8577,8584|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|8577,8584|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8592,8603|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8592,8603|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Organic Chemical|SIMPLE_SEGMENT|8604,8617|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8604,8617|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8604,8617|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8604,8617|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8631,8634|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8631,8634|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|8638,8641|false|false|false|||Q6H
Finding|Gene or Genome|SIMPLE_SEGMENT|8642,8645|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8646,8650|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8646,8650|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8646,8650|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8646,8650|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Activity|SIMPLE_SEGMENT|8652,8656|false|false|false|C1948035|Hold (action)|hold
Event|Event|SIMPLE_SEGMENT|8652,8656|false|false|false|||hold
Finding|Functional Concept|SIMPLE_SEGMENT|8652,8656|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|SIMPLE_SEGMENT|8652,8656|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Event|Event|SIMPLE_SEGMENT|8661,8669|false|false|false|||sedation
Finding|Finding|SIMPLE_SEGMENT|8661,8669|false|false|false|C0235195;C5400562|Sedated state;Sedation|sedation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8661,8669|false|false|false|C0344106|Sedation procedure|sedation
Drug|Organic Chemical|SIMPLE_SEGMENT|8682,8693|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8682,8693|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8714,8723|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8714,8723|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8725,8735|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8725,8735|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8748,8751|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8748,8751|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8748,8751|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8748,8751|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8748,8751|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8757,8767|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8757,8767|false|false|false|C0016860|furosemide|Furosemide
Finding|Classification|SIMPLE_SEGMENT|8788,8798|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8788,8798|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|SIMPLE_SEGMENT|8799,8802|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|SIMPLE_SEGMENT|8799,8802|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|SIMPLE_SEGMENT|8803,8807|false|false|false|||Work
Event|Occupational Activity|SIMPLE_SEGMENT|8803,8807|false|false|false|C0043227|Work|Work
Event|Event|SIMPLE_SEGMENT|8815,8820|false|false|false|||check
Anatomy|Cell Component|SIMPLE_SEGMENT|8831,8834|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8831,8834|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|8850,8857|false|false|false|||results
Event|Event|SIMPLE_SEGMENT|8862,8866|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|8862,8866|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Finding|Idea or Concept|SIMPLE_SEGMENT|8873,8876|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|Fax
Finding|Intellectual Product|SIMPLE_SEGMENT|8873,8876|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|Fax
Event|Event|SIMPLE_SEGMENT|8886,8895|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8886,8895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8886,8895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8886,8895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8886,8895|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8886,8907|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8886,8907|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8896,8907|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8896,8907|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8896,8907|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|8909,8913|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8909,8913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8909,8913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8909,8913|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|8916,8925|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8916,8925|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8916,8925|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8916,8925|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8916,8925|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8916,8935|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8926,8935|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8926,8935|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8926,8935|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8926,8935|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8926,8935|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8937,8965|false|false|false|C0694549|Community-Acquired Pneumonia|Community Acquired Pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8956,8965|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|SIMPLE_SEGMENT|8956,8965|false|false|false|||Pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8966,8974|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|8966,8974|false|false|false|||Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8966,8983|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8966,8990|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes Mellitus Type 2
Finding|Gene or Genome|SIMPLE_SEGMENT|8984,8988|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|8984,8988|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|8984,8990|false|false|false|C0441730|Type 2|Type 2
Event|Event|SIMPLE_SEGMENT|8994,9003|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8994,9003|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8994,9003|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8994,9003|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8994,9003|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9004,9013|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9004,9013|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9004,9013|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9004,9013|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9015,9021|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9015,9028|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9015,9028|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9022,9028|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9022,9028|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9030,9035|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9030,9035|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|9040,9048|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|9040,9048|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|9050,9055|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9050,9072|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9050,9072|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9059,9072|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9059,9072|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9059,9072|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9074,9079|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|9074,9079|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9074,9079|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|9074,9079|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|9074,9079|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|9074,9079|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|9074,9079|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|9084,9095|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|9084,9095|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|9097,9105|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9097,9105|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9097,9105|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9106,9112|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9106,9112|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9106,9112|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9114,9124|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|9114,9124|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9114,9124|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9114,9124|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9114,9124|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9127,9138|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|9127,9138|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|9127,9138|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|9143,9152|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9143,9152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9143,9152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9143,9152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9143,9152|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9143,9165|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9143,9165|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9143,9165|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9153,9165|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9153,9165|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9153,9165|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|9167,9171|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|9192,9200|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|9208,9216|false|false|false|C1547192|Organization unit type - Hospital|hospital
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9223,9232|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|9223,9232|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|9245,9252|false|false|false|||started
Drug|Antibiotic|SIMPLE_SEGMENT|9256,9267|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|9256,9267|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|9283,9287|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|9291,9299|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|9314,9317|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9314,9317|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|9352,9360|false|false|false|C2984078;C3889124|A little bit;Only a Little|a little
Finding|Finding|SIMPLE_SEGMENT|9352,9364|false|false|false|C2984078|A little bit|a little bit
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9354,9360|false|false|false|C0023882|Little's Disease|little
Event|Event|SIMPLE_SEGMENT|9354,9360|false|false|false|||little
Finding|Finding|SIMPLE_SEGMENT|9354,9360|false|false|false|C3889124|Only a Little|little
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9361,9364|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Organic Chemical|SIMPLE_SEGMENT|9361,9364|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9361,9364|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Event|Event|SIMPLE_SEGMENT|9361,9364|false|false|false|||bit
Finding|Gene or Genome|SIMPLE_SEGMENT|9361,9364|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Intellectual Product|SIMPLE_SEGMENT|9361,9364|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Receptor|SIMPLE_SEGMENT|9361,9364|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9366,9376|false|false|false|C0011175|Dehydration|dehydrated
Event|Event|SIMPLE_SEGMENT|9366,9376|false|false|false|||dehydrated
Event|Event|SIMPLE_SEGMENT|9386,9390|false|false|false|||came
Event|Event|SIMPLE_SEGMENT|9402,9410|false|false|false|||received
Drug|Substance|SIMPLE_SEGMENT|9419,9425|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|9419,9425|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|9419,9425|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9419,9425|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|9430,9434|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|9435,9442|false|false|false|||hydrate
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9454,9460|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9454,9460|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9454,9460|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|9454,9460|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9454,9460|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9454,9460|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|SIMPLE_SEGMENT|9461,9467|false|false|false|||levels
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9476,9481|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9476,9481|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9476,9481|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9489,9492|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Organic Chemical|SIMPLE_SEGMENT|9489,9492|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9489,9492|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Finding|Gene or Genome|SIMPLE_SEGMENT|9489,9492|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Intellectual Product|SIMPLE_SEGMENT|9489,9492|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Receptor|SIMPLE_SEGMENT|9489,9492|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Event|Event|SIMPLE_SEGMENT|9493,9496|false|false|false|||low
Finding|Finding|SIMPLE_SEGMENT|9493,9496|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|9493,9496|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|9514,9520|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9514,9520|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|9521,9524|false|false|false|||due
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9532,9541|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|9532,9541|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|9532,9541|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9550,9555|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|9564,9571|false|false|false|||treated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9578,9587|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|9578,9587|false|false|false|||pneumonia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9594,9600|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9594,9600|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9594,9600|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|9594,9600|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9594,9600|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9594,9600|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|SIMPLE_SEGMENT|9601,9607|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|9608,9616|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|9633,9640|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|9633,9640|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|9646,9650|false|false|false|||made
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9659,9670|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9659,9670|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9659,9670|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9659,9670|false|false|false|C4284232|Medications|medications
Drug|Food|SIMPLE_SEGMENT|9682,9687|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|9682,9687|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|9682,9687|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9682,9687|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Antibiotic|SIMPLE_SEGMENT|9688,9700|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|SIMPLE_SEGMENT|9688,9700|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|SIMPLE_SEGMENT|9701,9706|false|false|false|||750mg
Finding|Idea or Concept|SIMPLE_SEGMENT|9724,9727|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9724,9727|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Sign or Symptom|SIMPLE_SEGMENT|9755,9770|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|SIMPLE_SEGMENT|9764,9770|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|9779,9783|false|false|false|||sick
Finding|Sign or Symptom|SIMPLE_SEGMENT|9779,9783|false|false|false|C0221423|Illness (finding)|sick
Event|Event|SIMPLE_SEGMENT|9799,9807|false|false|false|||hesitate
Event|Event|SIMPLE_SEGMENT|9811,9815|false|false|false|||call
Finding|Intellectual Product|SIMPLE_SEGMENT|9821,9833|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|9821,9833|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|9829,9833|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|9829,9833|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|9829,9833|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9829,9833|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9834,9843|false|false|false|C0804815||physician
Event|Event|SIMPLE_SEGMENT|9853,9859|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|9873,9885|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|9873,9885|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|9881,9885|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|9881,9885|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|9881,9885|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9881,9885|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9886,9892|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|9896,9905|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9896,9905|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9896,9905|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9896,9905|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9896,9905|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|9910,9919|false|false|false|||scheduled
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9945,9949|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|9950,9957|false|false|false|||checked
Event|Activity|SIMPLE_SEGMENT|9970,9981|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|9970,9981|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|10022,10030|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|10022,10030|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|10022,10030|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|10038,10042|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10038,10042|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10038,10042|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10038,10042|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10038,10045|false|false|false|C1555558|care of - AddressPartType|care of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10071,10075|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|10071,10075|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|10071,10075|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|10079,10087|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10088,10100|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10088,10100|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10088,10100|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

