 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Codeine|179,186
<EOL>|186,187
<EOL>|188,189
Attending|189,198
:|198,199
_|200,201
_|201,202
_|202,203
.|203,204
<EOL>|204,205
<EOL>|206,207
Fever|224,229
<EOL>|229,230
<EOL>|231,232
Major|232,237
Surgical|238,246
or|247,249
Invasive|250,258
Procedure|259,268
:|268,269
<EOL>|269,270
None|270,274
<EOL>|274,275
<EOL>|276,277
_|305,306
_|306,307
_|307,308
woman|309,314
with|315,319
stage|320,325
IV|326,328
lung|329,333
adenocarcinoma|334,348
on|349,351
<EOL>|352,353
pemetrexed|353,363
,|363,364
CAD|365,368
,|368,369
CVA|370,373
presented|374,383
with|384,388
fever|389,394
from|395,399
home|400,404
.|404,405
Patient|406,413
was|414,417
<EOL>|418,419
found|419,424
to|425,427
have|428,432
temp|433,437
of|438,440
101.9|441,446
by|447,449
husband|450,457
on|458,460
_|461,462
_|462,463
_|463,464
,|464,465
down|466,470
to|471,473
100.4|474,479
<EOL>|480,481
with|481,485
cool|486,490
compresses|491,501
and|502,505
acetaminophen|506,519
.|519,520
Patient|521,528
reports|529,536
having|537,543
<EOL>|544,545
had|545,548
intermittent|549,561
nonproductive|562,575
coughs|576,582
,|582,583
mild|584,588
sore|589,593
throat|594,600
,|600,601
and|602,605
<EOL>|606,607
nasal|607,612
congestion|613,623
for|624,627
the|628,631
past|632,636
3|637,638
weeks|639,644
.|644,645
She|646,649
states|650,656
that|657,661
she|662,665
might|666,671
<EOL>|672,673
be|673,675
now|676,679
more|680,684
tired|685,690
than|691,695
usual|696,701
.|701,702
Patient|703,710
was|711,714
referred|715,723
to|724,726
the|727,730
ED|731,733
.|733,734
<EOL>|734,735
<EOL>|735,736
In|736,738
ED|739,741
,|741,742
T|743,744
99.2|745,749
,|749,750
HR|751,753
96|754,756
,|756,757
BP|758,760
132|761,764
/|764,765
64|765,767
,|767,768
RR|769,771
16|772,774
,|774,775
95|776,778
%|778,779
RA|779,781
.|781,782
Exam|783,787
<EOL>|788,789
unremarkable|789,801
.|801,802
Labs|803,807
notable|808,815
for|816,819
ANC|820,823
1200|824,828
,|828,829
Na|830,832
129|833,836
,|836,837
Cr|838,840
2.5|841,844
(|845,846
recent|846,852
<EOL>|853,854
baseline|854,862
1.5|863,866
-|866,867
2.0|867,870
)|870,871
.|871,872
CXR|873,876
showed|877,883
old|884,887
LLL|888,891
consolidation|892,905
and|906,909
no|910,912
new|913,916
<EOL>|917,918
process|918,925
.|925,926
Admitted|927,935
to|936,938
OMED|939,943
for|944,947
further|948,955
management|956,966
.|966,967
<EOL>|968,969
<EOL>|970,971
ONCOLOGIC|993,1002
Stage|1013,1018
IV|1019,1021
lung|1022,1026
adenocarcinoma|1027,1041
:|1041,1042
<EOL>|1042,1043
-|1043,1044
In|1045,1047
_|1048,1049
_|1049,1050
_|1050,1051
:|1051,1052
diagnosed|1053,1062
with|1063,1067
stage|1068,1073
IV|1074,1076
lung|1077,1081
adenoca|1082,1089
after|1090,1095
<EOL>|1096,1097
admission|1097,1106
for|1107,1110
STEMI|1111,1116
.|1116,1117
Received|1118,1126
the|1127,1130
first|1131,1136
cycle|1137,1142
of|1143,1145
pemetrexed|1146,1156
on|1157,1159
<EOL>|1160,1161
_|1161,1162
_|1162,1163
_|1163,1164
.|1164,1165
Most|1166,1170
recent|1171,1177
chemo|1178,1183
was|1184,1187
C6|1188,1190
of|1191,1193
pemetrexed|1194,1204
on|1205,1207
_|1208,1209
_|1209,1210
_|1210,1211
<EOL>|1211,1212
-|1212,1213
She|1214,1217
had|1218,1221
been|1222,1226
treated|1227,1234
over|1235,1239
the|1240,1243
course|1244,1250
of|1251,1253
the|1254,1257
last|1258,1262
year|1263,1267
with|1268,1272
<EOL>|1273,1274
multiple|1274,1282
courses|1283,1290
of|1291,1293
antibiotics|1294,1305
for|1306,1309
RLL|1310,1313
pneumonia|1314,1323
,|1323,1324
which|1325,1330
failed|1331,1337
<EOL>|1338,1339
to|1339,1341
resolve|1342,1349
on|1350,1352
serial|1353,1359
chest|1360,1365
imaging|1366,1373
.|1373,1374
<EOL>|1375,1376
<EOL>|1376,1377
NON-ONCOLOGIC|1377,1390
#|1400,1401
Dyslipidemia|1402,1414
<EOL>|1414,1415
#|1415,1416
Hypertension|1417,1429
<EOL>|1431,1432
#|1432,1433
CAD|1434,1437
:|1437,1438
MI|1439,1441
in|1442,1444
_|1445,1446
_|1446,1447
_|1447,1448
and|1449,1452
subsequent|1453,1463
1|1464,1465
vessel|1466,1472
CABG|1473,1477
SVG|1478,1481
-|1482,1483
>|1483,1484
LAD|1484,1487
,|1487,1488
s|1489,1490
/|1490,1491
p|1491,1492
<EOL>|1493,1494
BMS|1494,1497
in|1498,1500
LAD|1501,1504
in|1505,1507
_|1508,1509
_|1509,1510
_|1510,1511
after|1512,1517
anterior|1518,1526
STEMI|1527,1532
<EOL>|1532,1533
#|1533,1534
CVA|1535,1538
-|1539,1540
small|1541,1546
left|1547,1551
posterior|1552,1561
frontal|1562,1569
infarct|1570,1577
in|1578,1580
_|1581,1582
_|1582,1583
_|1583,1584
<EOL>|1584,1585
small|1585,1590
PFO|1591,1594
<EOL>|1594,1595
#|1595,1596
Macular|1597,1604
Degereration|1605,1617
<EOL>|1617,1618
<EOL>|1619,1620
:|1634,1635
<EOL>|1635,1636
_|1636,1637
_|1637,1638
_|1638,1639
<EOL>|1639,1640
:|1654,1655
<EOL>|1655,1656
Her|1656,1659
father|1660,1666
died|1667,1671
due|1672,1675
to|1676,1678
CAD|1679,1682
at|1683,1685
age|1686,1689
_|1690,1691
_|1691,1692
_|1692,1693
.|1693,1694
Her|1695,1698
mother|1699,1705
had|1706,1709
stomach|1710,1717
<EOL>|1718,1719
cancer|1719,1725
and|1726,1729
osteosarcoma|1730,1742
.|1742,1743
No|1744,1746
history|1747,1754
of|1755,1757
lung|1758,1762
cancer|1763,1769
,|1769,1770
colon|1771,1776
cancer|1777,1783
<EOL>|1784,1785
or|1785,1787
breast|1788,1794
cancer|1795,1801
.|1801,1802
<EOL>|1802,1803
<EOL>|1804,1805
Gen|1820,1823
:|1823,1824
elderly|1825,1832
woman|1833,1838
in|1839,1841
NAD|1842,1845
<EOL>|1845,1846
HEENT|1846,1851
:|1851,1852
EOMI|1853,1857
,|1857,1858
OP|1859,1861
moist|1862,1867
without|1868,1875
lesion|1876,1882
<EOL>|1882,1883
Neck|1883,1887
:|1887,1888
supple|1889,1895
,|1895,1896
no|1897,1899
LAD|1900,1903
<EOL>|1903,1904
CV|1904,1906
:|1906,1907
RRR|1908,1911
,|1911,1912
normal|1913,1919
S1|1920,1922
/|1922,1923
S2|1923,1925
,|1925,1926
no|1927,1929
m|1930,1931
/|1931,1932
r|1932,1933
/|1933,1934
g|1934,1935
<EOL>|1935,1936
Lungs|1936,1941
:|1941,1942
Poor|1943,1947
aeration|1948,1956
at|1957,1959
L|1960,1961
base|1962,1966
<EOL>|1966,1967
Abd|1967,1970
:|1970,1971
soft|1972,1976
,|1976,1977
NT|1978,1980
,|1980,1981
ND|1982,1984
,|1984,1985
BS|1986,1988
present|1989,1996
<EOL>|1996,1997
Ext|1997,2000
:|2000,2001
no|2002,2004
c|2005,2006
/|2006,2007
c|2007,2008
/|2008,2009
e|2009,2010
<EOL>|2010,2011
<EOL>|2012,2013
Pertinent|2013,2022
Results|2023,2030
:|2030,2031
<EOL>|2031,2032
WBC|2032,2035
-|2035,2036
2|2036,2037
.|2037,2038
0|2038,2039
*|2039,2040
#|2040,2041
RBC|2042,2045
-|2045,2046
2|2046,2047
.|2047,2048
39|2048,2050
*|2050,2051
HGB|2052,2055
-|2055,2056
7|2056,2057
.|2057,2058
4|2058,2059
*|2059,2060
HCT|2061,2064
-|2064,2065
22|2065,2067
.|2067,2068
7|2068,2069
*|2069,2070
MCV|2071,2074
-|2074,2075
95|2075,2077
<EOL>|2077,2078
NEUTS|2078,2083
-|2083,2084
62|2084,2086
BANDS|2087,2092
-|2092,2093
2|2093,2094
LYMPHS|2095,2101
-|2101,2102
14|2102,2104
*|2104,2105
MONOS|2106,2111
-|2111,2112
13|2112,2114
*|2114,2115
EOS|2116,2119
-|2119,2120
4|2120,2121
BASOS|2122,2127
-|2127,2128
1|2128,2129
ATYPS|2130,2135
-|2135,2136
4|2136,2137
*|2137,2138
<EOL>|2139,2140
_|2140,2141
_|2141,2142
_|2142,2143
MYELOS|2144,2150
-|2150,2151
0|2151,2152
<EOL>|2152,2153
PLT|2153,2156
COUNT|2157,2162
-|2162,2163
111|2163,2166
*|2166,2167
#|2167,2168
<EOL>|2168,2169
GLUCOSE|2169,2176
-|2176,2177
124|2177,2180
*|2180,2181
UREA|2182,2186
N|2187,2188
-|2188,2189
57|2189,2191
*|2191,2192
CREAT|2193,2198
-|2198,2199
2|2199,2200
.|2200,2201
5|2201,2202
*|2202,2203
SODIUM|2204,2210
-|2210,2211
129|2211,2214
*|2214,2215
POTASSIUM|2216,2225
-|2225,2226
4.9|2226,2229
<EOL>|2230,2231
CHLORIDE|2231,2239
-|2239,2240
96|2240,2242
TOTAL|2243,2248
CO2|2249,2252
-|2252,2253
25|2253,2255
<EOL>|2255,2256
LACTATE|2256,2263
-|2263,2264
0.6|2264,2267
<EOL>|2267,2268
<EOL>|2268,2269
URINE|2269,2274
COLOR|2276,2281
-|2281,2282
Yellow|2282,2288
APPEAR|2289,2295
-|2295,2296
Clear|2296,2301
SP|2302,2304
_|2305,2306
_|2306,2307
_|2307,2308
<EOL>|2308,2309
URINE|2309,2314
BLOOD|2316,2321
-|2321,2322
TR|2322,2324
NITRITE|2325,2332
-|2332,2333
NEG|2333,2336
PROTEIN|2337,2344
-|2344,2345
25|2345,2347
GLUCOSE|2348,2355
-|2355,2356
NEG|2356,2359
KETONE|2360,2366
-|2366,2367
NEG|2367,2370
<EOL>|2371,2372
BILIRUBIN|2372,2381
-|2381,2382
NEG|2382,2385
UROBILNGN|2386,2395
-|2395,2396
NEG|2396,2399
PH|2400,2402
-|2402,2403
5.0|2403,2406
LEUK|2407,2411
-|2411,2412
NEG|2412,2415
<EOL>|2415,2416
URINE|2416,2421
_|2423,2424
_|2424,2425
_|2425,2426
BACTERIA|2427,2435
-|2435,2436
FEW|2436,2439
YEAST|2440,2445
-|2445,2446
NONE|2446,2450
_|2451,2452
_|2452,2453
_|2453,2454
TRANS|2455,2460
<EOL>|2461,2462
_|2462,2463
_|2463,2464
_|2464,2465
<EOL>|2465,2466
<EOL>|2466,2467
STUDIES|2467,2474
:|2474,2475
<EOL>|2475,2476
<EOL>|2476,2477
Chest|2477,2482
Xray|2483,2487
_|2488,2489
_|2489,2490
_|2490,2491
:|2491,2492
<EOL>|2493,2494
1|2494,2495
.|2495,2496
In|2497,2499
setting|2500,2507
of|2508,2510
extensive|2511,2520
bronchoalveolar|2521,2536
carcinoma|2537,2546
,|2546,2547
and|2548,2551
the|2552,2555
<EOL>|2556,2557
absence|2557,2564
of|2565,2567
<EOL>|2568,2569
recent|2569,2575
comparable|2576,2586
studies|2587,2594
,|2594,2595
new|2596,2599
pneumonia|2600,2609
would|2610,2615
be|2616,2618
difficult|2619,2628
to|2629,2631
<EOL>|2632,2633
recognize|2633,2642
in|2643,2645
the|2646,2649
right|2650,2655
lower|2656,2661
and|2662,2665
middle|2666,2672
lobes|2673,2678
.|2678,2679
<EOL>|2680,2681
<EOL>|2681,2682
CT|2682,2684
Chest|2685,2690
_|2691,2692
_|2692,2693
_|2693,2694
:|2694,2695
<EOL>|2696,2697
1.|2697,2699
Increased|2700,2709
bronchial|2710,2719
and|2720,2723
peribronchial|2724,2737
nodules|2738,2745
with|2746,2750
<EOL>|2751,2752
ground|2752,2758
-|2758,2759
glass|2759,2764
halos|2765,2770
<EOL>|2771,2772
since|2772,2777
_|2778,2779
_|2779,2780
_|2780,2781
,|2781,2782
predominating|2783,2796
upper|2797,2802
and|2803,2806
middle|2807,2813
lobes|2814,2819
,|2819,2820
most|2821,2825
<EOL>|2826,2827
consistent|2827,2837
with|2838,2842
infection|2843,2852
.|2852,2853
<EOL>|2854,2855
2.|2855,2857
Stable|2858,2864
right|2865,2870
lower|2871,2876
lobe|2877,2881
reticular|2882,2891
opacities|2892,2901
with|2902,2906
areas|2907,2912
of|2913,2915
<EOL>|2916,2917
consolidation|2917,2930
<EOL>|2931,2932
and|2932,2935
widespread|2936,2946
nodules|2947,2954
predominantly|2955,2968
involving|2969,2978
the|2979,2982
right|2983,2988
upper|2989,2994
<EOL>|2995,2996
and|2996,2999
middle|3000,3006
<EOL>|3007,3008
lobes|3008,3013
,|3013,3014
consistent|3015,3025
with|3026,3030
known|3031,3036
bronchioalveolar|3037,3053
cell|3054,3058
carcinoma|3059,3068
.|3068,3069
<EOL>|3070,3071
3.|3071,3073
Stable|3074,3080
large|3081,3086
left|3087,3091
thyroid|3092,3099
mass|3100,3104
.|3104,3105
<EOL>|3106,3107
4.|3107,3109
Stable|3110,3116
abdominal|3117,3126
aortic|3127,3133
intimal|3134,3141
calcification|3142,3155
displacement|3156,3168
.|3168,3169
<EOL>|3170,3171
5.|3171,3173
Stable|3174,3180
renal|3181,3186
cysts|3187,3192
.|3192,3193
Miniscule|3194,3203
nonobstructive|3204,3218
right|3219,3224
renal|3225,3230
<EOL>|3231,3232
calculus|3232,3240
.|3240,3241
<EOL>|3242,3243
6.|3243,3245
Moderate|3246,3254
emphysema|3255,3264
.|3264,3265
<EOL>|3265,3266
<EOL>|3267,3268
_|3291,3292
_|3292,3293
_|3293,3294
year|3295,3299
old|3300,3303
woman|3304,3309
with|3310,3314
stage|3315,3320
IV|3321,3323
lung|3324,3328
adenoca|3329,3336
,|3336,3337
CAD|3338,3341
who|3342,3345
presented|3346,3355
<EOL>|3356,3357
with|3357,3361
fever|3362,3367
at|3368,3370
home|3371,3375
.|3375,3376
<EOL>|3376,3377
<EOL>|3377,3378
#|3378,3379
.|3379,3380
Fever|3381,3386
:|3386,3387
She|3388,3391
presented|3392,3401
with|3402,3406
_|3407,3408
_|3408,3409
_|3409,3410
weeks|3411,3416
of|3417,3419
fatigue|3420,3427
,|3427,3428
nonproductive|3429,3442
<EOL>|3443,3444
cough|3444,3449
that|3450,3454
is|3455,3457
chronic|3458,3465
,|3465,3466
and|3467,3470
1|3471,3472
day|3473,3476
of|3477,3479
fevers|3480,3486
.|3486,3487
Chest|3489,3494
xray|3495,3499
was|3500,3503
<EOL>|3504,3505
unremarkable|3505,3517
but|3518,3521
could|3522,3527
not|3528,3531
rule|3532,3536
out|3537,3540
infection|3541,3550
given|3551,3556
the|3557,3560
location|3561,3569
<EOL>|3570,3571
of|3571,3573
her|3574,3577
lung|3578,3582
cancer|3583,3589
.|3589,3590
She|3592,3595
had|3596,3599
negative|3600,3608
blood|3609,3614
and|3615,3618
urine|3619,3624
cultures|3625,3633
.|3633,3634
<EOL>|3636,3637
She|3637,3640
underwent|3641,3650
CT|3651,3653
chest|3654,3659
on|3660,3662
admission|3663,3672
,|3672,3673
as|3674,3676
she|3677,3680
was|3681,3684
due|3685,3688
for|3689,3692
a|3693,3694
repeat|3695,3701
<EOL>|3702,3703
CT|3703,3705
scan|3706,3710
the|3711,3714
following|3715,3724
week|3725,3729
routinely|3730,3739
.|3739,3740
The|3742,3745
CT|3746,3748
chest|3749,3754
was|3755,3758
<EOL>|3759,3760
concerning|3760,3770
for|3771,3774
a|3775,3776
new|3777,3780
infectious|3781,3791
process|3792,3799
in|3800,3802
the|3803,3806
right|3807,3812
upper|3813,3818
and|3819,3822
<EOL>|3823,3824
middle|3824,3830
lobes|3831,3836
,|3836,3837
as|3838,3840
well|3841,3845
as|3846,3848
stable|3849,3855
areas|3856,3861
of|3862,3864
consolidation|3865,3878
and|3879,3882
<EOL>|3883,3884
nodules|3884,3891
consistent|3892,3902
with|3903,3907
bronchioalveolar|3908,3924
carcinoma|3925,3934
.|3934,3935
She|3937,3940
was|3941,3944
<EOL>|3945,3946
started|3946,3953
on|3954,3956
ceftriaxone|3957,3968
and|3969,3972
azithromycin|3973,3985
and|3986,3989
was|3990,3993
discharged|3994,4004
on|4005,4007
<EOL>|4008,4009
cefuroxime|4009,4019
and|4020,4023
azithromycin|4024,4036
.|4036,4037
She|4039,4042
was|4043,4046
also|4047,4051
discharged|4052,4062
on|4063,4065
home|4066,4070
<EOL>|4071,4072
oxygen|4072,4078
(|4079,4080
she|4080,4083
already|4084,4091
used|4092,4096
oxygen|4097,4103
sometimes|4104,4113
at|4114,4116
home|4117,4121
and|4122,4125
was|4126,4129
<EOL>|4130,4131
instructed|4131,4141
to|4142,4144
use|4145,4148
it|4149,4151
full|4152,4156
-|4156,4157
time|4157,4161
after|4162,4167
discharge|4168,4177
)|4177,4178
.|4178,4179
<EOL>|4179,4180
<EOL>|4180,4181
#|4181,4182
.|4182,4183
Acute|4184,4189
renal|4190,4195
failure|4196,4203
:|4203,4204
She|4205,4208
had|4209,4212
an|4213,4215
elevated|4216,4224
creatinine|4225,4235
on|4236,4238
<EOL>|4239,4240
admission|4240,4249
to|4250,4252
2.5|4253,4256
from|4257,4261
a|4262,4263
recent|4264,4270
baseline|4271,4279
of|4280,4282
1.3|4283,4286
-|4286,4287
1.8|4287,4290
.|4290,4291
This|4293,4297
was|4298,4301
<EOL>|4302,4303
felt|4303,4307
to|4308,4310
be|4311,4313
prerenal|4314,4322
azotemia|4323,4331
and|4332,4335
it|4336,4338
improved|4339,4347
with|4348,4352
IV|4353,4355
hydration|4356,4365
.|4365,4366
<EOL>|4368,4369
However|4369,4376
,|4376,4377
she|4378,4381
still|4382,4387
has|4388,4391
new|4392,4395
renal|4396,4401
insufficiency|4402,4415
and|4416,4419
would|4420,4425
likely|4426,4432
<EOL>|4433,4434
benefit|4434,4441
from|4442,4446
follow|4447,4453
-|4453,4454
up|4454,4456
with|4457,4461
nephrology|4462,4472
after|4473,4478
discharge|4479,4488
.|4488,4489
She|4491,4494
was|4495,4498
<EOL>|4499,4500
also|4500,4504
instructed|4505,4515
to|4516,4518
follow|4519,4525
a|4526,4527
low|4528,4531
potassium|4532,4541
diet|4542,4546
.|4546,4547
<EOL>|4547,4548
<EOL>|4548,4549
#|4549,4550
.|4550,4551
Hyponatremia|4552,4564
:|4564,4565
She|4566,4569
had|4570,4573
low|4574,4577
serum|4578,4583
sodium|4584,4590
on|4591,4593
admission|4594,4603
,|4603,4604
felt|4605,4609
to|4610,4612
<EOL>|4613,4614
be|4614,4616
related|4617,4624
to|4625,4627
hypovolemia|4628,4639
in|4640,4642
the|4643,4646
setting|4647,4654
of|4655,4657
her|4658,4661
illness|4662,4669
.|4669,4670
Her|4672,4675
<EOL>|4676,4677
sodium|4677,4683
improved|4684,4692
to|4693,4695
normal|4696,4702
levels|4703,4709
with|4710,4714
IV|4715,4717
fluids|4718,4724
.|4724,4725
<EOL>|4725,4726
<EOL>|4726,4727
#|4727,4728
.|4728,4729
Stage|4730,4735
IV|4736,4738
Lung|4739,4743
Adenocarcinoma|4744,4758
:|4758,4759
She|4760,4763
is|4764,4766
s|4767,4768
/|4768,4769
p|4769,4770
6|4771,4772
cycles|4773,4779
of|4780,4782
<EOL>|4783,4784
pemetrexed|4784,4794
.|4794,4795
She|4797,4800
should|4801,4807
follow|4808,4814
-|4814,4815
up|4815,4817
with|4818,4822
her|4823,4826
primary|4827,4834
oncologist|4835,4845
<EOL>|4846,4847
for|4847,4850
further|4851,4858
treatment|4859,4868
.|4868,4869
<EOL>|4869,4870
<EOL>|4870,4871
#|4871,4872
.|4872,4873
Anemia|4874,4880
:|4880,4881
She|4882,4885
was|4886,4889
given|4890,4895
1|4896,4897
unit|4898,4902
of|4903,4905
PRBCs|4906,4911
for|4912,4915
anemia|4916,4922
on|4923,4925
<EOL>|4926,4927
admission|4927,4936
.|4936,4937
Her|4939,4942
anemia|4943,4949
was|4950,4953
felt|4954,4958
to|4959,4961
be|4962,4964
related|4965,4972
to|4973,4975
her|4976,4979
recent|4980,4986
<EOL>|4987,4988
chemotherapy|4988,5000
.|5000,5001
<EOL>|5001,5002
<EOL>|5002,5003
#|5003,5004
.|5004,5005
CAD|5006,5009
:|5009,5010
She|5011,5014
was|5015,5018
continued|5019,5028
on|5029,5031
a|5032,5033
statin|5034,5040
,|5040,5041
aspirin|5042,5049
,|5049,5050
and|5051,5054
clopidogrel|5055,5066
.|5066,5067
<EOL>|5067,5068
<EOL>|5068,5069
#|5069,5070
.|5070,5071
HTN|5072,5075
:|5075,5076
She|5077,5080
was|5081,5084
continued|5085,5094
on|5095,5097
amlodipine|5098,5108
.|5108,5109
<EOL>|5109,5110
<EOL>|5111,5112
Medications|5112,5123
on|5124,5126
Admission|5127,5136
:|5136,5137
<EOL>|5137,5138
amlodipine|5138,5148
5|5149,5150
mg|5151,5153
daily|5154,5159
<EOL>|5159,5160
atorvastatin|5160,5172
80|5173,5175
mg|5176,5178
daily|5179,5184
<EOL>|5184,5185
clopidogrel|5185,5196
75|5197,5199
mg|5200,5202
daily|5203,5208
<EOL>|5208,5209
aspirin|5209,5216
81|5217,5219
mg|5220,5222
daily|5223,5228
<EOL>|5228,5229
ranitidine|5229,5239
150|5240,5243
mg|5244,5246
daily|5247,5252
<EOL>|5252,5253
folate|5253,5259
<EOL>|5259,5260
loperamide|5260,5270
prn|5271,5274
<EOL>|5274,5275
lorazepam|5275,5284
prn|5285,5288
<EOL>|5288,5289
metoclopramide|5289,5303
prn|5304,5307
<EOL>|5307,5308
ondansetron|5308,5319
prn|5320,5323
<EOL>|5323,5324
trazodone|5324,5333
50|5334,5336
mg|5337,5339
daily|5340,5345
prn|5346,5349
<EOL>|5349,5350
<EOL>|5350,5351
<EOL>|5352,5353
Discharge|5353,5362
Medications|5363,5374
:|5374,5375
<EOL>|5375,5376
1.|5376,5378
Amlodipine|5379,5389
5|5390,5391
mg|5392,5394
Tablet|5395,5401
Sig|5402,5405
:|5405,5406
One|5407,5410
(|5411,5412
1|5412,5413
)|5413,5414
Tablet|5415,5421
PO|5422,5424
DAILY|5425,5430
(|5431,5432
Daily|5432,5437
)|5437,5438
.|5438,5439
<EOL>|5441,5442
<EOL>|5442,5443
2.|5443,5445
Atorvastatin|5446,5458
80|5459,5461
mg|5462,5464
Tablet|5465,5471
Sig|5472,5475
:|5475,5476
One|5477,5480
(|5481,5482
1|5482,5483
)|5483,5484
Tablet|5485,5491
PO|5492,5494
once|5495,5499
a|5500,5501
day|5502,5505
.|5505,5506
<EOL>|5508,5509
<EOL>|5509,5510
3.|5510,5512
Clopidogrel|5513,5524
75|5525,5527
mg|5528,5530
Tablet|5531,5537
Sig|5538,5541
:|5541,5542
One|5543,5546
(|5547,5548
1|5548,5549
)|5549,5550
Tablet|5551,5557
PO|5558,5560
DAILY|5561,5566
<EOL>|5567,5568
(|5568,5569
Daily|5569,5574
)|5574,5575
.|5575,5576
<EOL>|5578,5579
4.|5579,5581
Aspirin|5582,5589
81|5590,5592
mg|5593,5595
Tablet|5596,5602
,|5602,5603
Chewable|5604,5612
Sig|5613,5616
:|5616,5617
One|5618,5621
(|5622,5623
1|5623,5624
)|5624,5625
Tablet|5626,5632
,|5632,5633
Chewable|5634,5642
<EOL>|5643,5644
PO|5644,5646
DAILY|5647,5652
(|5653,5654
Daily|5654,5659
)|5659,5660
.|5660,5661
<EOL>|5663,5664
5.|5664,5666
Ranitidine|5667,5677
HCl|5678,5681
150|5682,5685
mg|5686,5688
Tablet|5689,5695
Sig|5696,5699
:|5699,5700
One|5701,5704
(|5705,5706
1|5706,5707
)|5707,5708
Tablet|5709,5715
PO|5716,5718
DAILY|5719,5724
<EOL>|5725,5726
(|5726,5727
Daily|5727,5732
)|5732,5733
.|5733,5734
<EOL>|5736,5737
6.|5737,5739
Folic|5740,5745
Acid|5746,5750
1|5751,5752
mg|5753,5755
Tablet|5756,5762
Sig|5763,5766
:|5766,5767
One|5768,5771
(|5772,5773
1|5773,5774
)|5774,5775
Tablet|5776,5782
PO|5783,5785
DAILY|5786,5791
(|5792,5793
Daily|5793,5798
)|5798,5799
.|5799,5800
<EOL>|5802,5803
<EOL>|5803,5804
7.|5804,5806
Loperamide|5807,5817
2|5818,5819
mg|5820,5822
Tablet|5823,5829
Sig|5830,5833
:|5833,5834
One|5835,5838
(|5839,5840
1|5840,5841
)|5841,5842
Tablet|5843,5849
PO|5850,5852
four|5853,5857
times|5858,5863
a|5864,5865
<EOL>|5866,5867
day|5867,5870
as|5871,5873
needed|5874,5880
for|5881,5884
diarrhea|5885,5893
.|5893,5894
<EOL>|5896,5897
8.|5897,5899
Lorazepam|5900,5909
Oral|5911,5915
<EOL>|5915,5916
9.|5916,5918
Metoclopramide|5919,5933
Oral|5935,5939
<EOL>|5939,5940
10.|5940,5943
Zofran|5944,5950
Oral|5952,5956
<EOL>|5956,5957
11.|5957,5960
Trazodone|5961,5970
50|5971,5973
mg|5974,5976
Tablet|5977,5983
Sig|5984,5987
:|5987,5988
One|5989,5992
(|5993,5994
1|5994,5995
)|5995,5996
Tablet|5997,6003
PO|6004,6006
at|6007,6009
bedtime|6010,6017
as|6018,6020
<EOL>|6021,6022
needed|6022,6028
for|6029,6032
insomnia|6033,6041
.|6041,6042
<EOL>|6044,6045
12.|6045,6048
Azithromycin|6049,6061
250|6062,6065
mg|6066,6068
Tablet|6069,6075
Sig|6076,6079
:|6079,6080
One|6081,6084
(|6085,6086
1|6086,6087
)|6087,6088
Tablet|6089,6095
PO|6096,6098
Q24H|6099,6103
<EOL>|6104,6105
(|6105,6106
every|6106,6111
24|6112,6114
hours|6115,6120
)|6120,6121
for|6122,6125
3|6126,6127
days|6128,6132
:|6132,6133
First|6134,6139
dose|6140,6144
on|6145,6147
_|6148,6149
_|6149,6150
_|6150,6151
.|6151,6152
<EOL>|6152,6153
Disp|6153,6157
:|6157,6158
*|6158,6159
3|6159,6160
Tablet|6161,6167
(|6167,6168
s|6168,6169
)|6169,6170
*|6170,6171
Refills|6172,6179
:|6179,6180
*|6180,6181
0|6181,6182
*|6182,6183
<EOL>|6183,6184
13.|6184,6187
Cefuroxime|6188,6198
Axetil|6199,6205
500|6206,6209
mg|6210,6212
Tablet|6213,6219
Sig|6220,6223
:|6223,6224
One|6225,6228
(|6229,6230
1|6230,6231
)|6231,6232
Tablet|6233,6239
PO|6240,6242
twice|6243,6248
<EOL>|6249,6250
a|6250,6251
day|6252,6255
for|6256,6259
8|6260,6261
days|6262,6266
:|6266,6267
First|6268,6273
dose|6274,6278
on|6279,6281
night|6282,6287
of|6288,6290
_|6291,6292
_|6292,6293
_|6293,6294
.|6294,6295
Please|6296,6302
take|6303,6307
<EOL>|6308,6309
antibiotic|6309,6319
to|6320,6322
its|6323,6326
completion|6327,6337
.|6337,6338
<EOL>|6338,6339
Disp|6339,6343
:|6343,6344
*|6344,6345
17|6345,6347
Tablet|6348,6354
(|6354,6355
s|6355,6356
)|6356,6357
*|6357,6358
Refills|6359,6366
:|6366,6367
*|6367,6368
0|6368,6369
*|6369,6370
<EOL>|6370,6371
14.|6371,6374
Senna|6375,6380
8.6|6381,6384
mg|6385,6387
Tablet|6388,6394
Sig|6395,6398
:|6398,6399
One|6400,6403
(|6404,6405
1|6405,6406
)|6406,6407
Tablet|6408,6414
PO|6415,6417
twice|6418,6423
a|6424,6425
day|6426,6429
as|6430,6432
<EOL>|6433,6434
needed|6434,6440
for|6441,6444
constipation|6445,6457
.|6457,6458
<EOL>|6460,6461
15.|6461,6464
Metoprolol|6465,6475
Tartrate|6476,6484
50|6485,6487
mg|6488,6490
Tablet|6491,6497
Sig|6498,6501
:|6501,6502
One|6503,6506
(|6507,6508
1|6508,6509
)|6509,6510
Tablet|6511,6517
PO|6518,6520
BID|6521,6524
<EOL>|6525,6526
(|6526,6527
2|6527,6528
times|6529,6534
a|6535,6536
day|6537,6540
)|6540,6541
.|6541,6542
<EOL>|6544,6545
16|6545,6547
.|6547,6548
Polyethylene|6549,6561
Glycol|6562,6568
3350|6569,6573
17|6574,6576
gram|6577,6581
/|6581,6582
dose|6582,6586
Powder|6587,6593
Sig|6594,6597
:|6597,6598
One|6599,6602
(|6603,6604
1|6604,6605
)|6605,6606
<EOL>|6608,6609
PO|6609,6611
DAILY|6612,6617
(|6618,6619
Daily|6619,6624
)|6624,6625
as|6626,6628
needed|6629,6635
for|6636,6639
constipation|6640,6652
.|6652,6653
<EOL>|6655,6656
<EOL>|6657,6658
Discharge|6658,6667
Disposition|6668,6679
:|6679,6680
<EOL>|6680,6681
Home|6681,6685
With|6686,6690
Service|6691,6698
<EOL>|6698,6699
<EOL>|6700,6701
Facility|6701,6709
:|6709,6710
<EOL>|6710,6711
_|6711,6712
_|6712,6713
_|6713,6714
<EOL>|6715,6716
<EOL>|6717,6718
Discharge|6718,6727
Diagnosis|6728,6737
:|6737,6738
<EOL>|6738,6739
Community|6758,6767
-|6767,6768
Acquired|6768,6776
Pneumonia|6777,6786
<EOL>|6786,6787
<EOL>|6787,6788
Secondary|6788,6797
Diagnosis|6798,6807
:|6807,6808
<EOL>|6808,6809
Non-small|6809,6818
cell|6819,6823
lung|6824,6828
cancer|6829,6835
<EOL>|6835,6836
Coronary|6836,6844
Artery|6845,6851
Disease|6852,6859
<EOL>|6859,6860
<EOL>|6860,6861
<EOL>|6862,6863
Mental|6884,6890
Status|6891,6897
:|6897,6898
Clear|6899,6904
and|6905,6908
coherent|6909,6917
.|6917,6918
<EOL>|6918,6919
Level|6919,6924
of|6925,6927
Consciousness|6928,6941
:|6941,6942
Alert|6943,6948
and|6949,6952
interactive|6953,6964
.|6964,6965
<EOL>|6965,6966
Activity|6966,6974
Status|6975,6981
:|6981,6982
Ambulatory|6983,6993
-|6994,6995
Independent|6996,7007
.|7007,7008
<EOL>|7008,7009
<EOL>|7009,7010
<EOL>|7011,7012
You|7036,7039
were|7040,7044
admitted|7045,7053
to|7054,7056
the|7057,7060
hospital|7061,7069
after|7070,7075
a|7076,7077
fever|7078,7083
.|7083,7084
You|7086,7089
underwent|7090,7099
<EOL>|7100,7101
a|7101,7102
CT|7103,7105
scan|7106,7110
of|7111,7113
your|7114,7118
chest|7119,7124
that|7125,7129
showed|7130,7136
that|7137,7141
you|7142,7145
likely|7146,7152
have|7153,7157
<EOL>|7158,7159
pneumonia|7159,7168
in|7169,7171
your|7172,7176
right|7177,7182
lung|7183,7187
.|7187,7188
You|7190,7193
were|7194,7198
started|7199,7206
on|7207,7209
antibiotics|7210,7221
<EOL>|7222,7223
to|7223,7225
treat|7226,7231
this|7232,7236
pneumonia|7237,7246
.|7246,7247
<EOL>|7247,7248
<EOL>|7248,7249
You|7249,7252
now|7253,7256
have|7257,7261
an|7262,7264
increased|7265,7274
oxygen|7275,7281
requirement|7282,7293
and|7294,7297
should|7298,7304
ALWAYS|7305,7311
<EOL>|7312,7313
wear|7313,7317
supplemental|7318,7330
oxygen|7331,7337
at|7338,7340
rate|7341,7345
of|7346,7348
2|7349,7350
liters|7351,7357
per|7358,7361
minute|7362,7368
.|7368,7369
<EOL>|7369,7370
<EOL>|7370,7371
You|7371,7374
also|7375,7379
had|7380,7383
a|7384,7385
low|7386,7389
blood|7390,7395
count|7396,7401
and|7402,7405
were|7406,7410
given|7411,7416
a|7417,7418
blood|7419,7424
<EOL>|7425,7426
transfusion|7426,7437
.|7437,7438
It|7440,7442
was|7443,7446
felt|7447,7451
that|7452,7456
your|7457,7461
blood|7462,7467
count|7468,7473
was|7474,7477
low|7478,7481
due|7482,7485
to|7486,7488
<EOL>|7489,7490
chemotherapy|7490,7502
.|7502,7503
<EOL>|7503,7504
<EOL>|7504,7505
You|7505,7508
should|7509,7515
weigh|7516,7521
yourself|7522,7530
every|7531,7536
morning|7537,7544
and|7545,7548
call|7549,7553
your|7554,7558
doctor|7559,7565
if|7566,7568
<EOL>|7569,7570
you|7570,7573
gain|7574,7578
more|7579,7583
than|7584,7588
3|7589,7590
pounds|7591,7597
or|7598,7600
notice|7601,7607
increasing|7608,7618
shortness|7619,7628
of|7629,7631
<EOL>|7632,7633
breath|7633,7639
,|7639,7640
or|7641,7643
leg|7644,7647
swelling|7648,7656
.|7656,7657
<EOL>|7657,7658
<EOL>|7658,7659
Changes|7659,7666
to|7667,7669
your|7670,7674
medications|7675,7686
:|7686,7687
<EOL>|7687,7688
ADDED|7688,7693
continuous|7694,7704
supplemental|7705,7717
oxygen|7718,7724
at|7725,7727
2|7728,7729
liters|7730,7736
per|7737,7740
minute|7741,7747
<EOL>|7747,7748
ADDED|7748,7753
cefuroxime|7754,7764
500|7765,7768
mg|7769,7771
BID|7772,7775
for|7776,7779
8|7780,7781
more|7782,7786
days|7787,7791
<EOL>|7791,7792
ADDED|7792,7797
azithromycin|7798,7810
250mg|7811,7816
by|7817,7819
mouth|7820,7825
for|7826,7829
3|7830,7831
more|7832,7836
days|7837,7841
<EOL>|7841,7842
ADDED|7842,7847
Senna|7848,7853
1|7854,7855
tab|7856,7859
twice|7860,7865
daily|7866,7871
as|7872,7874
needed|7875,7881
for|7882,7885
constipation|7886,7898
<EOL>|7898,7899
ADDED|7899,7904
Polyethylene|7905,7917
Glycol|7918,7924
(|7925,7926
Miralax|7926,7933
)|7933,7934
1|7935,7936
packet|7937,7943
daily|7944,7949
as|7950,7952
needed|7953,7959
for|7960,7963
<EOL>|7964,7965
constipation|7965,7977
<EOL>|7977,7978
<EOL>|7979,7980
Followup|7980,7988
Instructions|7989,8001
:|8001,8002
<EOL>|8002,8003
_|8003,8004
_|8004,8005
_|8005,8006
<EOL>|8006,8007

