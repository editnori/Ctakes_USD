 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|210,225|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|216,225|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|216,225|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Functional Concept|SIMPLE_SEGMENT|227,231|false|true|false|C1552822|Table Cell Horizontal Align - left|Left
Finding|Finding|SIMPLE_SEGMENT|232,240|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|232,245|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|232,251|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|241,245|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|241,245|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|241,251|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|246,251|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|246,251|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|246,251|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Classification|SIMPLE_SEGMENT|254,259|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|272,290|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|281,290|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|281,290|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|281,290|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|281,290|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|292,296|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Finding|Idea or Concept|SIMPLE_SEGMENT|297,304|false|false|false|C1550516|Target Awareness - partial|partial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|305,311|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|312,322|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|312,322|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|312,322|false|false|false|C0002688|Amputation|amputation
Finding|Conceptual Entity|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|326,333|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|326,336|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|326,352|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|326,352|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|337,344|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|337,344|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|337,352|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|345,352|false|false|false|C0221423|Illness (finding)|Illness
Finding|Functional Concept|SIMPLE_SEGMENT|363,380|false|false|false|C3853134|Poorly controlled|poorly controlled
Finding|Finding|SIMPLE_SEGMENT|370,380|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Functional Concept|SIMPLE_SEGMENT|370,380|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Idea or Concept|SIMPLE_SEGMENT|370,380|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|381,389|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|406,417|false|false|false|C0035309|Retinal Diseases|retinopathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|419,429|false|false|false|C0442874|Neuropathy|neuropathy
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|431,434|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|431,434|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|431,434|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|431,434|false|false|false|C2347441|Pad Dosage Form|PAD
Finding|Gene or Genome|SIMPLE_SEGMENT|431,434|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|431,434|false|false|false|C3814046|PAD Regimen|PAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|436,440|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|436,440|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|436,446|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|441,446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|441,446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|441,446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|449,455|false|false|false|C0018534|Hallux structure|hallux
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|458,461|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|458,461|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|458,461|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|458,461|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|476,480|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|486,495|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|486,495|false|false|false|C0027415|Narcotics|narcotics
Attribute|Clinical Attribute|SIMPLE_SEGMENT|496,505|false|false|false|C4255433||agreement
Finding|Intellectual Product|SIMPLE_SEGMENT|496,505|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Social Behavior|SIMPLE_SEGMENT|496,505|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|530,540|false|false|false|C2979880||subjective
Finding|Finding|SIMPLE_SEGMENT|530,540|false|false|false|C2266644|subjective (symptom)|subjective
Finding|Finding|SIMPLE_SEGMENT|542,547|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|542,547|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|549,555|false|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|SIMPLE_SEGMENT|567,571|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|567,571|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|567,571|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|SIMPLE_SEGMENT|577,582|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|577,586|false|false|false|C0018534|Hallux structure|great toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|583,586|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Body Substance|SIMPLE_SEGMENT|604,609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|604,609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|604,609|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Body Substance|SIMPLE_SEGMENT|639,644|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|639,644|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|639,644|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|673,676|false|false|false|C0282612|Prostatic Intraepithelial Neoplasias|pin
Finding|Gene or Genome|SIMPLE_SEGMENT|673,676|false|false|false|C1825012|DYNLL1 gene|pin
Finding|Conceptual Entity|SIMPLE_SEGMENT|693,697|false|false|false|C1711300;C2243104|Span - parameter;span - body measurement finding|span
Finding|Finding|SIMPLE_SEGMENT|693,697|false|false|false|C1711300;C2243104|Span - parameter;span - body measurement finding|span
Finding|Intellectual Product|SIMPLE_SEGMENT|703,707|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|730,736|false|false|false|C0039515|Tennis (activity)|tennis
Finding|Idea or Concept|SIMPLE_SEGMENT|743,752|false|false|false|C0449450|Presentation|Presented
Finding|Intellectual Product|SIMPLE_SEGMENT|760,766|false|false|false|C1546403;C1546845;C1547230;C1561556|Admission Type - Urgent;Certification patient type - Urgent;Triage Code - Urgent;Visit Priority Code - Urgent|urgent
Event|Activity|SIMPLE_SEGMENT|767,771|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|767,771|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|767,771|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Sign or Symptom|SIMPLE_SEGMENT|792,799|false|false|false|C0015967|Fever|febrile
Drug|Organic Chemical|SIMPLE_SEGMENT|814,821|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|814,821|false|false|false|C0699142|Tylenol|Tylenol
Finding|Finding|SIMPLE_SEGMENT|842,850|false|false|false|C0277797|Apyrexial|afebrile
Event|Activity|SIMPLE_SEGMENT|873,880|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|873,880|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Functional Concept|SIMPLE_SEGMENT|889,898|false|false|false|C0443318|Sustained|sustained
Finding|Finding|SIMPLE_SEGMENT|899,910|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Finding|SIMPLE_SEGMENT|914,917|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|914,917|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|950,955|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|950,955|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|950,955|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|950,955|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|959,963|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|971,977|false|false|false|C0018534|Hallux structure|hallux
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|988,992|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|988,992|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|988,992|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Finding|SIMPLE_SEGMENT|996,1000|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|996,1000|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|996,1000|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1005,1018|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1020,1026|false|false|false|C0885876|X-rays, Homeopathic Preparations|X-rays
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1020,1026|false|false|false|C0043309|Roentgen Rays|X-rays
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1020,1026|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|X-rays
Finding|Functional Concept|SIMPLE_SEGMENT|1032,1036|false|false|false|C0443157|Bony|bony
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1037,1044|false|false|false|C0333307|Superficial ulcer|erosion
Finding|Pathologic Function|SIMPLE_SEGMENT|1037,1044|false|false|false|C1959609|Erosion lesion|erosion
Finding|Functional Concept|SIMPLE_SEGMENT|1052,1064|true|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1065,1068|true|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1065,1068|true|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|SIMPLE_SEGMENT|1065,1068|true|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Finding|Gene or Genome|SIMPLE_SEGMENT|1065,1068|true|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|SIMPLE_SEGMENT|1065,1068|true|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|SIMPLE_SEGMENT|1065,1068|true|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|SIMPLE_SEGMENT|1065,1068|true|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1070,1074|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Finding|Functional Concept|SIMPLE_SEGMENT|1070,1074|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|SIMPLE_SEGMENT|1070,1074|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|SIMPLE_SEGMENT|1070,1074|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Drug|Antibiotic|SIMPLE_SEGMENT|1082,1093|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Idea or Concept|SIMPLE_SEGMENT|1098,1105|false|false|false|C1550516|Target Awareness - partial|partial
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|1106,1116|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|1106,1116|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1106,1116|false|false|false|C0002688|Amputation|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1106,1134|false|false|false|C4316611|Amputation of left great toe|amputation of left great toe
Finding|Functional Concept|SIMPLE_SEGMENT|1120,1124|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Gene or Genome|SIMPLE_SEGMENT|1125,1130|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1125,1134|false|false|false|C0018534|Hallux structure|great toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1131,1134|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1160,1163|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1160,1163|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1164,1168|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1164,1168|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1164,1168|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1170,1178|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1170,1178|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1180,1199|false|false|false|C0848390|excessive urination|excessive urination
Finding|Organism Function|SIMPLE_SEGMENT|1190,1199|false|false|false|C0042034|Urination|urination
Finding|Finding|SIMPLE_SEGMENT|1201,1212|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Sign or Symptom|SIMPLE_SEGMENT|1201,1212|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Finding|SIMPLE_SEGMENT|1214,1221|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1214,1221|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1223,1228|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1223,1228|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1223,1233|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1223,1233|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1229,1233|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1229,1233|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1229,1233|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|1248,1255|false|false|false|C1555582|Initial (abbreviation)|Initial
Drug|Food|SIMPLE_SEGMENT|1256,1261|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1256,1267|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|1256,1267|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|1262,1267|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1262,1267|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|SIMPLE_SEGMENT|1286,1294|false|false|false|C0277797|Apyrexial|afebrile
Finding|Finding|SIMPLE_SEGMENT|1296,1307|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Finding|Functional Concept|SIMPLE_SEGMENT|1330,1334|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1330,1334|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|1352,1356|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1352,1356|false|false|false|C0687712|warming process|warm
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1395,1399|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1395,1399|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1401,1406|false|false|false|C0024109|Lung|lungs
Finding|Idea or Concept|SIMPLE_SEGMENT|1407,1412|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1417,1420|false|false|false|C0022681|Medullary sponge kidney|MSK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1417,1420|false|false|false|C0022681|Medullary sponge kidney|MSK
Finding|Gene or Genome|SIMPLE_SEGMENT|1417,1420|false|false|false|C1420279|SIK1 gene|MSK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1422,1430|false|false|false|C0041834|Erythema|erythema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1443,1450|false|false|false|C0018534|Hallux structure|big toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1447,1450|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Social Behavior|SIMPLE_SEGMENT|1467,1475|false|false|false|C0678975|inferiority|inferior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1476,1480|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1476,1480|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|1476,1480|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1476,1480|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|1476,1480|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|1476,1480|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Mental Process|SIMPLE_SEGMENT|1482,1492|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1482,1492|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Finding|Intellectual Product|SIMPLE_SEGMENT|1508,1512|false|false|false|C1705483|Pathname|path
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1508,1512|false|false|false|C0919386|Pathology procedure|path
Finding|Gene or Genome|SIMPLE_SEGMENT|1516,1521|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1535,1541|false|false|false|C0489800|Posterior part of left leg|L calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1537,1541|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1537,1541|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Functional Concept|SIMPLE_SEGMENT|1543,1550|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Intellectual Product|SIMPLE_SEGMENT|1543,1550|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1568,1575|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|plantar
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1568,1583|false|false|false|C0231784|Plantar flexion|plantar flexion
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1576,1583|false|false|false|C1525443|W flexion|flexion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1576,1583|false|false|false|C0231452||flexion
Finding|Functional Concept|SIMPLE_SEGMENT|1585,1592|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Intellectual Product|SIMPLE_SEGMENT|1585,1592|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Finding|SIMPLE_SEGMENT|1593,1596|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|SIMPLE_SEGMENT|1593,1596|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1593,1596|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1600,1605|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1600,1605|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1610,1613|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Mental Process|SIMPLE_SEGMENT|1615,1621|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1615,1628|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|1615,1628|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1622,1628|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|1622,1628|false|false|false|C1546481|What subject filter - Status|Status
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1636,1641|false|false|false|C1517938|Long Interspersed Elements|Lines
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1636,1641|false|false|false|C1517938|Long Interspersed Elements|Lines
Finding|Idea or Concept|SIMPLE_SEGMENT|1636,1641|false|false|false|C1548328|Lines Quantity Limit Request|Lines
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1656,1662|false|false|false|C0230371|Structure of left hand|L hand
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1658,1662|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|SIMPLE_SEGMENT|1658,1662|false|false|false|C0741992|Hand problem|hand
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1664,1668|false|false|false|C0587081|Laboratory test finding|Labs
Drug|Organic Chemical|SIMPLE_SEGMENT|1750,1757|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1750,1757|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1750,1757|false|false|false|C0202115|Lactic acid measurement|Lactate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1795,1799|false|false|false|C0722071|Neut brand of sodium bicarbonate|neut
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1795,1799|false|false|false|C0722071|Neut brand of sodium bicarbonate|neut
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1795,1799|false|false|false|C0027944|Neutralization Tests|neut
Procedure|Research Activity|SIMPLE_SEGMENT|1814,1821|false|false|false|C0947630|Scientific Study|Studies
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1842,1846|false|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1842,1846|false|false|false|C0043299|Diagnostic radiologic examination|Xray
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1847,1851|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|Foot
Finding|Finding|SIMPLE_SEGMENT|1847,1851|false|false|false|C0555980|Foot problem|Foot
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1855,1858|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|Lat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1855,1858|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|Lat
Drug|Immunologic Factor|SIMPLE_SEGMENT|1855,1858|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|Lat
Finding|Gene or Genome|SIMPLE_SEGMENT|1855,1858|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|Lat
Finding|Functional Concept|SIMPLE_SEGMENT|1865,1869|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Finding|Conceptual Entity|SIMPLE_SEGMENT|1878,1882|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1878,1882|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Intellectual Product|SIMPLE_SEGMENT|1878,1882|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1878,1882|false|false|false|C4723641|Nucleotide Sequence Read|read
Finding|Pathologic Function|SIMPLE_SEGMENT|1905,1915|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1933,1939|false|false|false|C4522154|Distal Resection Margin|distal
Finding|Gene or Genome|SIMPLE_SEGMENT|1954,1959|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1954,1963|false|false|false|C0018534|Hallux structure|great toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1960,1963|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1968,1975|false|false|false|C0333307|Superficial ulcer|erosion
Finding|Pathologic Function|SIMPLE_SEGMENT|1968,1975|false|false|false|C1959609|Erosion lesion|erosion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1993,1997|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1993,1997|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|1993,1997|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1993,1997|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|1993,1997|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|1993,1997|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2005,2011|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2005,2019|false|false|false|C0576464;C3669027|Bone structure of distal phalanx|distal phalanx
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2012,2019|false|false|false|C0222682;C0223792|Phalanx of hand;Phalanx structure|phalanx
Finding|Gene or Genome|SIMPLE_SEGMENT|2027,2032|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2033,2036|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Intellectual Product|SIMPLE_SEGMENT|2072,2080|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2082,2090|false|false|false|C2926606||Findings
Finding|Functional Concept|SIMPLE_SEGMENT|2082,2090|false|false|false|C2607943|findings aspects|Findings
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2120,2133|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Gene or Genome|SIMPLE_SEGMENT|2138,2141|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2138,2141|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|2138,2141|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2138,2155|false|false|false|C0202671|MRI with contrast|MRI with contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|2147,2155|false|false|false|C0009924|Contrast Media|contrast
Event|Activity|SIMPLE_SEGMENT|2187,2197|false|false|false|C1516048|Assessed|assessment
Finding|Intellectual Product|SIMPLE_SEGMENT|2187,2197|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2187,2197|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|SIMPLE_SEGMENT|2187,2197|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Finding|Body Substance|SIMPLE_SEGMENT|2201,2208|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2201,2208|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2201,2208|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Antibiotic|SIMPLE_SEGMENT|2220,2232|false|false|false|C0031955|piperacillin|Piperacillin
Drug|Organic Chemical|SIMPLE_SEGMENT|2220,2232|false|false|false|C0031955|piperacillin|Piperacillin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2220,2243|false|false|false|C0250480|piperacillin-tazobactam combination|Piperacillin-Tazobactam
Drug|Antibiotic|SIMPLE_SEGMENT|2233,2243|false|false|false|C0075870|tazobactam|Tazobactam
Drug|Organic Chemical|SIMPLE_SEGMENT|2233,2243|false|false|false|C0075870|tazobactam|Tazobactam
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2246,2256|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|2246,2256|false|false|false|C0042313|vancomycin|Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2246,2256|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Procedure|Health Care Activity|SIMPLE_SEGMENT|2258,2266|false|false|false|C0009818|Consultation|Consults
Finding|Functional Concept|SIMPLE_SEGMENT|2288,2296|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|2288,2296|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|2288,2296|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|SIMPLE_SEGMENT|2343,2350|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2343,2350|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2358,2363|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2396,2399|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2396,2399|false|false|false|C2346952|Bachelor of Education|bed
Finding|Sign or Symptom|SIMPLE_SEGMENT|2414,2420|false|false|false|C0085593|Chills|chills
Finding|Functional Concept|SIMPLE_SEGMENT|2451,2455|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2451,2460|false|false|false|C0230461|Structure of left foot|Left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2456,2460|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|2456,2460|false|false|false|C0555980|Foot problem|foot
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2478,2486|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|2478,2486|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|2478,2486|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|2478,2486|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2478,2486|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Idea or Concept|SIMPLE_SEGMENT|2516,2522|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|2516,2522|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|2516,2525|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2516,2533|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2516,2533|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|2526,2533|false|false|false|C0449913|System|SYSTEMS
Drug|Organic Chemical|SIMPLE_SEGMENT|2536,2544|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2536,2544|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Vitamin|SIMPLE_SEGMENT|2536,2544|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Finding|Functional Concept|SIMPLE_SEGMENT|2536,2544|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Finding|Idea or Concept|SIMPLE_SEGMENT|2536,2544|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2545,2548|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2545,2548|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2545,2548|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|SIMPLE_SEGMENT|2545,2548|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2545,2548|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Finding|Gene or Genome|SIMPLE_SEGMENT|2545,2548|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2545,2548|false|false|false|C0489633|Review of systems (procedure)|ROS
Finding|Classification|SIMPLE_SEGMENT|2575,2583|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2575,2583|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2575,2583|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|2586,2606|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|2591,2598|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2591,2598|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2591,2598|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2591,2598|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2591,2606|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2599,2606|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2599,2606|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2599,2606|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2609,2613|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2609,2613|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2609,2613|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2615,2618|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2615,2618|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2615,2618|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2615,2618|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2615,2618|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2615,2618|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2615,2618|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2623,2626|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2627,2635|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2636,2639|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2636,2639|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2636,2639|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2645,2648|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2645,2648|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2645,2648|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2645,2648|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2645,2648|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2645,2648|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2645,2648|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2656,2659|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2656,2659|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2656,2659|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2665,2668|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2665,2668|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2665,2668|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2665,2668|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2665,2668|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2665,2668|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2665,2668|false|false|false|C1413980|DES gene|DES
Finding|Conceptual Entity|SIMPLE_SEGMENT|2672,2676|false|false|false|C2697523|Graph Edge|edge
Finding|Cell Function|SIMPLE_SEGMENT|2678,2681|false|false|false|C5445058|integrated stress response signaling|ISR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2689,2692|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2689,2692|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2689,2692|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2693,2696|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2693,2696|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2693,2696|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2693,2696|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2693,2696|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2693,2696|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2693,2696|false|false|false|C1413980|DES gene|DES
Finding|Pathologic Function|SIMPLE_SEGMENT|2701,2709|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2710,2716|false|false|false|C4522154|Distal Resection Margin|distal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2731,2734|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2731,2734|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2731,2734|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2731,2734|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2731,2734|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2731,2734|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2731,2734|false|false|false|C1413980|DES gene|DES
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2756,2760|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2766,2769|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2766,2769|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2766,2769|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2794,2804|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2794,2804|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2794,2804|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2814,2818|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2822,2834|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2836,2845|false|false|false|C0149931|Migraine Disorders|Migraines
Finding|Intellectual Product|SIMPLE_SEGMENT|2847,2854|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|2847,2854|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2847,2868|false|false|false|C0748678|shoulder pain chronic|Chronic shoulder pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2855,2863|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2855,2863|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2855,2863|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Sign or Symptom|SIMPLE_SEGMENT|2855,2868|false|false|false|C0037011|Shoulder Pain|shoulder pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2864,2868|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2864,2868|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2864,2868|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2872,2881|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2872,2881|false|false|false|C0027415|Narcotics|narcotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2883,2886|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2883,2886|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2883,2886|false|false|false|C0764906|OSA protein, Drosophila|OSA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2888,2909|false|false|false|C0031117;C4721453|Peripheral Nervous System Diseases;Peripheral Neuropathy|Peripheral neuropathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2899,2909|false|false|false|C0442874|Neuropathy|neuropathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|2911,2919|false|false|false|C0085631;C3887611|Agitation;Restlessness|Restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2911,2923|false|false|false|C0035258|Restless Legs Syndrome|Restless leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2920,2923|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|SIMPLE_SEGMENT|2926,2932|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2926,2940|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2933,2940|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2933,2940|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2933,2940|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2946,2952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2946,2952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2946,2952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2946,2952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2946,2960|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2953,2960|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2953,2960|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2953,2960|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Body Substance|SIMPLE_SEGMENT|2962,2969|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2962,2969|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2962,2969|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Classification|SIMPLE_SEGMENT|3021,3027|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3021,3027|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3021,3027|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3021,3027|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|3021,3035|false|false|false|C0241889|Family Medical History|family history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3028,3035|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3028,3035|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3028,3035|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Idea or Concept|SIMPLE_SEGMENT|3037,3043|false|false|false|C1546508|Relationship - Mother|Mother
Finding|Finding|SIMPLE_SEGMENT|3049,3057|false|false|false|C0332149|Possible|possible
Drug|Organic Chemical|SIMPLE_SEGMENT|3058,3065|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3058,3065|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|3058,3065|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3058,3071|false|true|false|C0085762|Alcohol abuse|alcohol abuse
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3066,3071|false|false|false|C0013146|Drug abuse|abuse
Event|Event|SIMPLE_SEGMENT|3066,3071|false|false|false|C1546935|Abuse|abuse
Finding|Finding|SIMPLE_SEGMENT|3066,3071|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Conceptual Entity|SIMPLE_SEGMENT|3073,3079|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3073,3079|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Finding|SIMPLE_SEGMENT|3081,3089|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Finding|Organism Function|SIMPLE_SEGMENT|3081,3089|false|false|false|C0011065;C1549464;C1704456|Cessation of life;Deceased - ActIneligibilityReason;Deceased - Military Status|deceased
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3102,3109|false|false|false|C0019829|Hodgkin Disease|Hodgkin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3102,3119|false|false|false|C0019829|Hodgkin Disease|Hodgkin's Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3112,3119|false|false|false|C0012634|Disease|Disease
Finding|Idea or Concept|SIMPLE_SEGMENT|3128,3135|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|3128,3135|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Finding|SIMPLE_SEGMENT|3139,3147|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3139,3147|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3139,3147|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3139,3152|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3139,3152|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3148,3152|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3148,3152|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3154,3163|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|SIMPLE_SEGMENT|3164,3168|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3164,3168|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|SIMPLE_SEGMENT|3231,3238|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3231,3238|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3240,3245|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3240,3245|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3240,3245|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|3240,3245|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3240,3245|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3240,3245|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3250,3261|false|false|false|C1704675|Interaction|interactive
Finding|Finding|SIMPLE_SEGMENT|3263,3283|false|false|false|C2051415|patient appears in no acute distress (physical finding)|In no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|3269,3274|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|3275,3283|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3275,3283|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3285,3290|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3298,3301|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3298,3301|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3303,3310|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3303,3310|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Gene or Genome|SIMPLE_SEGMENT|3320,3323|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3324,3329|false|false|false|C0024109|Lung|LUNGS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3343,3346|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|3343,3346|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3343,3346|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3351,3358|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3351,3358|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3351,3358|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3360,3364|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3379,3383|false|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3379,3393|false|false|false|C0278328|Deep palpation|deep palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3384,3393|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3421,3426|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|3421,3433|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3427,3433|false|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3435,3446|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Functional Concept|SIMPLE_SEGMENT|3448,3452|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3448,3457|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3453,3457|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|3453,3457|false|false|false|C0555980|Foot problem|foot
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3475,3483|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3475,3483|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|3475,3483|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|3475,3483|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3475,3483|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Functional Concept|SIMPLE_SEGMENT|3492,3504|false|false|false|C0332476|erythematous|erythematous
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3527,3532|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3527,3532|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3533,3537|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3533,3537|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3546,3551|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3546,3551|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|3564,3570|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3564,3570|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3564,3570|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|SIMPLE_SEGMENT|3595,3600|false|false|false|C1513492|motor movement|motor
Finding|Finding|SIMPLE_SEGMENT|3595,3609|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3595,3609|false|false|false|C0234130|Motor function (observable entity)|motor function
Finding|Finding|SIMPLE_SEGMENT|3601,3609|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3601,3609|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3601,3609|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3601,3609|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|SIMPLE_SEGMENT|3618,3624|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Body Substance|SIMPLE_SEGMENT|3627,3636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3627,3636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3627,3636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3627,3636|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|SIMPLE_SEGMENT|3637,3641|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3637,3641|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|SIMPLE_SEGMENT|3691,3698|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3691,3698|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3691,3709|false|false|false|C1148118||General Appearance
Finding|Finding|SIMPLE_SEGMENT|3691,3709|false|false|false|C1148438|general appearance (physical finding)|General Appearance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3699,3709|false|false|false|C0550215||Appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|3699,3709|false|false|false|C2051406|patient appearance regarding mental status exam|Appearance
Finding|Finding|SIMPLE_SEGMENT|3711,3715|false|false|false|C5575035|Well (answer to question)|Well
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3728,3731|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3728,3731|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3728,3731|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3728,3731|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3728,3731|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|3728,3731|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3733,3738|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3767,3773|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3767,3773|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3767,3773|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|SIMPLE_SEGMENT|3774,3783|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3789,3792|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3789,3792|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3797,3810|false|false|false|C0521367|Oropharyngeal|oropharyngeal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3797,3810|false|false|false|C0553694|Disorder of oropharynx|oropharyngeal
Finding|Functional Concept|SIMPLE_SEGMENT|3797,3810|false|false|false|C1522409|Oropharyngeal Route of Administration|oropharyngeal
Finding|Finding|SIMPLE_SEGMENT|3811,3818|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3823,3826|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3823,3826|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3823,3826|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3828,3833|false|false|false|C0024109|Lung|Lungs
Finding|Intellectual Product|SIMPLE_SEGMENT|3835,3840|false|false|false|C1549782|Relational Operator - Equal|Equal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3841,3846|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3841,3846|false|false|false|C0741025|Chest problem|chest
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3841,3851|false|false|false|C5570649|Chest rise|chest rise
Drug|Organic Chemical|SIMPLE_SEGMENT|3847,3851|false|false|false|C0246719|risedronate|rise
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3847,3851|false|false|false|C0246719|risedronate|rise
Finding|Intellectual Product|SIMPLE_SEGMENT|3847,3851|false|false|false|C4321377|Relational and Item-Specific Encoding Task|rise
Finding|Idea or Concept|SIMPLE_SEGMENT|3853,3857|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3858,3861|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3858,3861|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3858,3861|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|3858,3861|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3858,3861|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3858,3861|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3858,3870|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|3862,3870|false|false|false|C0026649|Movement|movement
Finding|Finding|SIMPLE_SEGMENT|3875,3884|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|3875,3884|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Event|Occupational Activity|SIMPLE_SEGMENT|3885,3889|true|false|false|C0043227|Work|work
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3893,3902|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|3893,3902|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|3893,3902|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|3893,3902|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3893,3902|false|false|false|C1160636|respiratory system process|breathing
Finding|Finding|SIMPLE_SEGMENT|3904,3927|false|false|false|C0238844|Decreased breath sounds|Decreased breath sounds
Finding|Body Substance|SIMPLE_SEGMENT|3914,3920|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3914,3927|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3921,3927|false|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3931,3934|false|false|false|C1261077|Structure of left lower lobe of lung|LLL
Finding|Finding|SIMPLE_SEGMENT|3936,3941|false|false|false|C0034642;C0240859|Basilar Rales;Rales|Rales
Finding|Functional Concept|SIMPLE_SEGMENT|3945,3949|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3950,3954|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3950,3954|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3950,3954|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3950,3954|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|3950,3954|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|3950,3954|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Sign or Symptom|SIMPLE_SEGMENT|3960,3967|false|false|false|C0043144|Wheezing|wheezes
Finding|Finding|SIMPLE_SEGMENT|3971,3978|false|false|false|C0035508|Rhonchi|rhonchi
Finding|Finding|SIMPLE_SEGMENT|4007,4014|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|4028,4032|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4037,4044|false|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|SIMPLE_SEGMENT|4045,4051|false|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4060,4067|false|false|false|C0007272|Carotid Arteries|carotid
Drug|Food|SIMPLE_SEGMENT|4068,4074|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4068,4074|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4068,4074|false|false|false|C0034107|Pulse taking|pulses
Finding|Conceptual Entity|SIMPLE_SEGMENT|4083,4089|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|SIMPLE_SEGMENT|4090,4096|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4090,4096|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4090,4096|false|false|false|C0034107|Pulse taking|pulses
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4105,4125|false|false|false|C1706488|Dorsalis pedis pulse|dorsalis pedis pulse
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4120,4125|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|4120,4125|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|4120,4125|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|4120,4125|false|false|false|C0034107|Pulse taking|pulse
Finding|Functional Concept|SIMPLE_SEGMENT|4129,4134|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|SIMPLE_SEGMENT|4136,4142|false|false|false|C1299582|Unable|unable
Finding|Functional Concept|SIMPLE_SEGMENT|4157,4161|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Procedure|Health Care Activity|SIMPLE_SEGMENT|4169,4177|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4169,4177|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4178,4185|false|false|false|C2346961|Bandage Dosage Form|bandage
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4187,4194|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4187,4194|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|4187,4194|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4211,4216|false|false|false|C0021853|Intestines|Bowel
Finding|Finding|SIMPLE_SEGMENT|4211,4223|false|false|false|C0232693|Bowel sounds|Bowel sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4217,4223|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|4224,4231|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4224,4231|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4233,4237|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4254,4263|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4277,4288|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4293,4301|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|SIMPLE_SEGMENT|4305,4313|true|false|false|C0010520|Cyanosis|cyanosis
Finding|Functional Concept|SIMPLE_SEGMENT|4315,4319|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4315,4324|false|false|false|C0230461|Structure of left foot|Left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4320,4324|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|4320,4324|false|false|false|C0555980|Foot problem|foot
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4325,4333|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4325,4333|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|4325,4333|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|4325,4333|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4325,4333|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Activity|SIMPLE_SEGMENT|4334,4339|false|false|false|C1947930|Cleaning (activity)|clean
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4347,4355|false|false|false|C0041834|Erythema|Erythema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4360,4365|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4360,4365|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|4373,4379|false|false|false|C4761388||margin
Procedure|Health Care Activity|SIMPLE_SEGMENT|4383,4391|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4383,4391|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4392,4396|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|4392,4396|false|false|false|C1546778||site
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4416,4422|false|false|false|C0502420|Suture Joint|Suture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4416,4422|false|false|false|C1706068|Suture Dosage Form|Suture
Finding|Intellectual Product|SIMPLE_SEGMENT|4416,4422|false|false|false|C1546803||Suture
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4416,4422|false|false|false|C0009068|Closure by suture|Suture
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4423,4427|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|4423,4427|false|false|false|C1546778||site
Event|Activity|SIMPLE_SEGMENT|4431,4436|false|false|false|C1947930|Cleaning (activity)|clean
Drug|Substance|SIMPLE_SEGMENT|4445,4448|true|false|false|C0444185|Pus specimen|pus
Finding|Body Substance|SIMPLE_SEGMENT|4445,4448|true|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Finding|Intellectual Product|SIMPLE_SEGMENT|4445,4448|true|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Anatomy|Body System|SIMPLE_SEGMENT|4450,4454|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4450,4454|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4450,4454|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|4450,4454|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|4450,4454|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Sign or Symptom|SIMPLE_SEGMENT|4459,4465|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Finding|SIMPLE_SEGMENT|4469,4476|true|false|false|C0221198|Lesion|lesions
Procedure|Health Care Activity|SIMPLE_SEGMENT|4485,4493|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4485,4493|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4494,4498|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|4494,4498|false|false|false|C1546778||site
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4514,4520|false|false|false|C5890614||person
Finding|Intellectual Product|SIMPLE_SEGMENT|4514,4520|false|false|false|C1522390|Person Info|person
Event|Activity|SIMPLE_SEGMENT|4522,4527|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|4522,4527|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4522,4527|false|false|false|C1533810||place
Finding|Finding|SIMPLE_SEGMENT|4533,4537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|4533,4537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|4533,4537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|4559,4565|false|false|false|C1554187|Gender Status - Intact|intact
Procedure|Health Care Activity|SIMPLE_SEGMENT|4588,4597|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4598,4602|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4630,4635|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4630,4635|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4636,4639|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4646,4649|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4646,4649|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4646,4649|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4655,4658|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4655,4658|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4655,4658|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4655,4658|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4664,4667|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4664,4667|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4674,4677|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4674,4677|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4674,4677|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4674,4677|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4681,4684|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4681,4684|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4681,4684|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4681,4684|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4681,4684|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4691,4695|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4721,4724|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4741,4746|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4741,4746|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4759,4765|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4772,4777|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4772,4777|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4772,4777|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4783,4786|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4783,4786|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4889,4894|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4889,4894|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4889,4902|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4889,4902|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4889,4902|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4895,4902|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4895,4902|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4895,4902|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4895,4902|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4895,4902|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4949,4953|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4949,4953|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4949,4953|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4980,4985|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4980,4985|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4986,4989|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|SIMPLE_SEGMENT|4986,4989|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Finding|Gene or Genome|SIMPLE_SEGMENT|4986,4989|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5009,5014|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5009,5014|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Classification|SIMPLE_SEGMENT|5019,5022|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|5019,5022|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5019,5022|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5027,5031|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5027,5031|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5056,5060|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5056,5060|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|5056,5060|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5056,5060|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|5056,5060|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|5056,5060|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5079,5084|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5079,5084|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5079,5092|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|5085,5092|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5085,5092|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5085,5092|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|SIMPLE_SEGMENT|5110,5115|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5110,5115|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5110,5115|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5110,5121|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5116,5121|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5116,5121|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|SIMPLE_SEGMENT|5122,5127|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|SIMPLE_SEGMENT|5135,5140|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|5160,5165|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5160,5165|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5160,5165|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5160,5171|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5166,5171|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|5166,5171|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Finding|Finding|SIMPLE_SEGMENT|5172,5175|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5176,5183|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5176,5183|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5176,5183|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Finding|Finding|SIMPLE_SEGMENT|5184,5187|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5188,5195|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5188,5195|false|false|false|C0033684|Proteins|Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|5188,5195|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5188,5195|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5201,5208|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5201,5208|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5201,5208|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5201,5208|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5201,5208|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5215,5221|false|false|false|C0022634|Ketones|Ketone
Finding|Finding|SIMPLE_SEGMENT|5234,5237|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5246,5249|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|5280,5285|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5280,5285|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5280,5285|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5280,5289|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|SIMPLE_SEGMENT|5286,5289|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5286,5289|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5286,5289|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|5293,5296|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|SIMPLE_SEGMENT|5313,5318|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|5313,5318|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5313,5318|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5313,5318|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5325,5328|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5325,5328|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5325,5328|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|5325,5328|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|5325,5328|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5325,5328|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|5325,5328|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|5325,5328|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5325,5328|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|SIMPLE_SEGMENT|5353,5358|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5353,5358|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5353,5358|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5353,5365|false|false|false|C0455910|Mucus in urine (finding)|URINE Mucous
Finding|Body Substance|SIMPLE_SEGMENT|5359,5365|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|Mucous
Finding|Gene or Genome|SIMPLE_SEGMENT|5366,5370|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Finding|Intellectual Product|SIMPLE_SEGMENT|5383,5391|false|false|false|C1552654|Parameterized Data Type - Interval|INTERVAL
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5392,5396|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5433,5438|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5433,5438|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5439,5442|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5439,5442|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5439,5442|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5439,5442|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5439,5442|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5439,5442|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5439,5442|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5446,5449|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5446,5449|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5446,5449|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5446,5449|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5446,5449|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5446,5449|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5456,5459|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|5456,5459|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Finding|Finding|SIMPLE_SEGMENT|5456,5459|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5456,5459|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5465,5472|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5465,5472|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Finding|Body Substance|SIMPLE_SEGMENT|5492,5501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5492,5501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5492,5501|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5492,5501|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5502,5506|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5534,5539|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5534,5539|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5540,5543|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5548,5551|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5548,5551|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5548,5551|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5558,5561|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5558,5561|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5558,5561|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5558,5561|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5567,5570|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5567,5570|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5578,5581|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5578,5581|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5578,5581|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5578,5581|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5586,5589|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5586,5589|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5586,5589|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5586,5589|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5586,5589|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5595,5599|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5625,5628|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5645,5650|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5645,5650|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5645,5658|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5645,5658|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5645,5658|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5651,5658|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5651,5658|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5651,5658|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5651,5658|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5651,5658|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5705,5709|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5705,5709|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5705,5709|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5734,5739|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5734,5739|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5734,5747|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5740,5747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5740,5747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5740,5747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5740,5747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5740,5747|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5740,5747|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5740,5747|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5780,5785|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5780,5785|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5786,5789|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|SIMPLE_SEGMENT|5786,5789|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Finding|Gene or Genome|SIMPLE_SEGMENT|5786,5789|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Finding|Finding|SIMPLE_SEGMENT|5797,5804|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5797,5804|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Functional Concept|SIMPLE_SEGMENT|5813,5817|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5813,5822|false|false|false|C0230461|Structure of left foot|LEFT FOOT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5818,5822|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|FOOT
Finding|Finding|SIMPLE_SEGMENT|5818,5822|false|false|false|C0555980|Foot problem|FOOT
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5823,5827|false|false|false|C0043309|Roentgen Rays|XRAY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5823,5827|false|false|false|C0043299|Diagnostic radiologic examination|XRAY
Finding|Intellectual Product|SIMPLE_SEGMENT|5834,5844|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5834,5844|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Pathologic Function|SIMPLE_SEGMENT|5869,5879|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5897,5903|false|false|false|C4522154|Distal Resection Margin|distal
Finding|Gene or Genome|SIMPLE_SEGMENT|5919,5924|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5919,5928|false|false|false|C0018534|Hallux structure|great toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5925,5928|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5933,5940|false|false|false|C0333307|Superficial ulcer|erosion
Finding|Pathologic Function|SIMPLE_SEGMENT|5933,5940|false|false|false|C1959609|Erosion lesion|erosion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5958,5962|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5958,5962|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|5958,5962|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5958,5962|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|5958,5962|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|5958,5962|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5970,5976|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5970,5984|false|false|false|C0576464;C3669027|Bone structure of distal phalanx|distal phalanx
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5977,5984|false|false|false|C0222682;C0223792|Phalanx of hand;Phalanx structure|phalanx
Finding|Gene or Genome|SIMPLE_SEGMENT|5993,5998|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5993,6002|false|false|false|C0018534|Hallux structure|great toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5999,6002|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Intellectual Product|SIMPLE_SEGMENT|6062,6070|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6073,6081|false|false|false|C2926606||Findings
Finding|Functional Concept|SIMPLE_SEGMENT|6073,6081|false|false|false|C2607943|findings aspects|Findings
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6110,6123|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Gene or Genome|SIMPLE_SEGMENT|6128,6131|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6128,6131|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|6128,6131|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6128,6145|false|false|false|C0202671|MRI with contrast|MRI with contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6137,6145|false|false|false|C0009924|Contrast Media|contrast
Event|Activity|SIMPLE_SEGMENT|6177,6187|false|false|false|C1516048|Assessed|assessment
Finding|Intellectual Product|SIMPLE_SEGMENT|6177,6187|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6177,6187|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|SIMPLE_SEGMENT|6177,6187|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6217,6225|false|false|false|C2926606||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|6217,6225|false|false|false|C2607943|findings aspects|FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|6237,6242|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6259,6266|false|false|false|C0554756|Doppler studies|Doppler
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6267,6276|false|false|false|C0450448|Waveforms|waveforms
Finding|Functional Concept|SIMPLE_SEGMENT|6294,6299|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6300,6307|false|false|false|C0015811|Femur|femoral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6309,6318|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6339,6347|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|6339,6347|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|6339,6347|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|6350,6356|false|false|false|C0332197|Absent|Absent
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6350,6356|false|false|false|C5237010|Expression Negative|Absent
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6357,6365|false|false|false|C0450448|Waveforms|waveform
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6374,6383|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6384,6390|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6384,6397|false|false|false|C0085427|Tibial Arteries|tibial artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6391,6397|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6391,6397|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|SIMPLE_SEGMENT|6403,6408|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6409,6412|false|false|false|C1328319;C3888326|Ankle brachial pressure index (observable entity)|ABI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6469,6476|false|false|false|C0005847|Blood Vessel|vessels
Finding|Functional Concept|SIMPLE_SEGMENT|6487,6491|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6508,6515|false|false|false|C0554756|Doppler studies|Doppler
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6516,6525|false|false|false|C0450448|Waveforms|waveforms
Finding|Functional Concept|SIMPLE_SEGMENT|6543,6547|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6548,6555|false|false|false|C0015811|Femur|femoral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6560,6569|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6560,6578|false|false|false|C0032649|Structure of popliteal artery|popliteal arteries
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6570,6578|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|6570,6578|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|6570,6578|false|false|false|C0397581|Procedure on artery|arteries
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6592,6601|false|false|false|C0450448|Waveforms|waveforms
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6619,6628|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6629,6635|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6655,6663|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|6655,6663|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|6655,6663|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|6669,6673|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6674,6677|false|false|false|C1328319;C3888326|Ankle brachial pressure index (observable entity)|ABI
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6704,6709|false|false|false|C0232117|Pulse Rate|Pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|6704,6709|false|false|false|C0391850|Physiologic pulse|Pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6704,6709|false|false|false|C1947910|Pulse phenomenon|Pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|6704,6709|false|false|false|C0034107|Pulse taking|Pulse
Finding|Finding|SIMPLE_SEGMENT|6704,6716|false|false|false|C0425580|Pulse volume|Pulse volume
Finding|Intellectual Product|SIMPLE_SEGMENT|6710,6716|false|false|false|C1705102|Volume (publication)|volume
Finding|Functional Concept|SIMPLE_SEGMENT|6774,6779|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6780,6784|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6780,6784|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6786,6791|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6786,6791|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6796,6806|false|false|false|C0025584|Metatarsal bone structure|metatarsal
Finding|Intellectual Product|SIMPLE_SEGMENT|6810,6820|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6810,6820|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Idea or Concept|SIMPLE_SEGMENT|6825,6836|false|false|false|C0750502|Significant|Significant
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6847,6853|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6854,6862|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6854,6876|false|false|false|C0003834|Arterial insufficiency|arterial insufficiency
Finding|Functional Concept|SIMPLE_SEGMENT|6863,6876|false|false|false|C0231179|Insufficiency|insufficiency
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6884,6889|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6884,6889|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6891,6902|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Functional Concept|SIMPLE_SEGMENT|6903,6910|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6906,6910|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6906,6910|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6906,6910|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|6906,6910|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|6906,6910|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Idea or Concept|SIMPLE_SEGMENT|6917,6928|false|false|false|C0750502|Significant|significant
Finding|Functional Concept|SIMPLE_SEGMENT|6936,6941|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6949,6952|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|6974,6984|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6974,6984|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Activity|SIMPLE_SEGMENT|6989,6999|false|false|false|C1707455|Comparison|Comparison
Finding|Functional Concept|SIMPLE_SEGMENT|7021,7027|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7021,7027|true|false|false|C4319952|Change - procedure|change
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7057,7064|false|false|false|C0038293|Sternum|sternal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7057,7070|false|false|false|C0407260|Wiring of sternum|sternal wires
Finding|Intellectual Product|SIMPLE_SEGMENT|7089,7093|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Functional Concept|SIMPLE_SEGMENT|7113,7123|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7113,7129|false|false|false|C0011666;C1305624|Descending aorta|descending aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7124,7129|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|7124,7129|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7155,7160|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7155,7160|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|7155,7160|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Tissue|SIMPLE_SEGMENT|7166,7173|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7166,7173|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|7166,7183|true|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|7174,7183|true|false|false|C0013687|effusion|effusions
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7190,7199|false|false|false|C0032285|Pneumonia|pneumonia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7204,7213|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7204,7213|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7204,7213|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7204,7219|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7214,7219|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7214,7219|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|SIMPLE_SEGMENT|7222,7225|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7222,7225|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|7222,7225|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Functional Concept|SIMPLE_SEGMENT|7226,7230|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7226,7235|false|false|false|C0230461|Structure of left foot|LEFT FOOT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7231,7235|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|FOOT
Finding|Finding|SIMPLE_SEGMENT|7231,7235|false|false|false|C0555980|Foot problem|FOOT
Finding|Intellectual Product|SIMPLE_SEGMENT|7242,7252|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|7242,7252|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|7274,7279|false|false|false|C0002690;C1514517;C4522245;C5848682|Amputation Stumps;Atypical Spitz Nevus;Neoplasm of uncertain behavior of smooth muscle;Prostate Stromal Proliferation of Uncertain Malignant Potential|stump
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7274,7279|false|false|false|C0002690;C1514517;C4522245;C5848682|Amputation Stumps;Atypical Spitz Nevus;Neoplasm of uncertain behavior of smooth muscle;Prostate Stromal Proliferation of Uncertain Malignant Potential|stump
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7280,7284|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7280,7291|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|7280,7291|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|7285,7291|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|7285,7291|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7300,7307|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|plantar
Anatomy|Tissue|SIMPLE_SEGMENT|7308,7311|false|false|false|C0001527|Adipose tissue|fat
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7308,7311|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7308,7311|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Organic Chemical|SIMPLE_SEGMENT|7308,7311|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7308,7311|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Finding|Gene or Genome|SIMPLE_SEGMENT|7308,7311|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Finding|Receptor|SIMPLE_SEGMENT|7308,7311|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7308,7311|false|false|false|C0279453|doxorubicin/fluorouracil/triazinate protocol|fat
Anatomy|Tissue|SIMPLE_SEGMENT|7308,7315|false|false|false|C0935625|Fat pad|fat pad
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|7312,7315|false|false|false|C3669270|Strucure of thick cushion of skin|pad
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7312,7315|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7312,7315|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7312,7315|false|false|false|C2347441|Pad Dosage Form|pad
Finding|Gene or Genome|SIMPLE_SEGMENT|7312,7315|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|pad
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7312,7315|false|false|false|C3814046|PAD Regimen|pad
Finding|Intellectual Product|SIMPLE_SEGMENT|7327,7333|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7334,7343|false|false|false|C0222682;C0223792|Phalanx of hand;Phalanx structure|phalanges
Anatomy|Tissue|SIMPLE_SEGMENT|7372,7378|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|7372,7378|false|false|false|C1547928|Tissue Specimen Code|tissue
Finding|Idea or Concept|SIMPLE_SEGMENT|7384,7392|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7384,7395|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7407,7414|false|false|false|C0000833|Abscess|abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|7407,7414|false|false|false|C1546533||abscess
Finding|Functional Concept|SIMPLE_SEGMENT|7424,7429|false|false|false|C1285542|Has focus|focus
Finding|Finding|SIMPLE_SEGMENT|7433,7436|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|7433,7436|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7440,7446|false|false|false|C1710082|Signal|signal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7452,7457|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7452,7457|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7470,7476|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7478,7484|false|false|false|C0007776;C1176472|Cerebral cortex;Cortex of Organ|cortex
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7478,7484|false|false|false|C0001614;C0595905|Adrenal Cortex Diseases;cortex bone disorders|cortex
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7492,7508|false|false|false|C0459701|First metatarsal structure|first metatarsal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7498,7508|false|false|false|C0025584|Metatarsal bone structure|metatarsal
Event|Activity|SIMPLE_SEGMENT|7548,7558|false|false|false|C1707455|Comparison|comparison
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7548,7564|false|false|false|C0489479;C1579762|Comparison study;comparative study research|comparison study
Procedure|Research Activity|SIMPLE_SEGMENT|7548,7564|false|false|false|C0489479;C1579762|Comparison study;comparative study research|comparison study
Finding|Intellectual Product|SIMPLE_SEGMENT|7559,7564|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|7559,7564|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Functional Concept|SIMPLE_SEGMENT|7569,7574|false|false|false|C1285542|Has focus|focus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7578,7591|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7617,7622|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|7617,7622|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|7617,7622|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7617,7622|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Pathologic Function|SIMPLE_SEGMENT|7617,7629|false|false|false|C0544791|Inflammatory fistula|sinus tracts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7623,7629|false|false|false|C1185740|Tract|tracts
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7644,7648|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7644,7648|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7644,7648|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7644,7648|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7656,7672|false|false|false|C0459701|First metatarsal structure|first metatarsal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7662,7672|false|false|false|C0025584|Metatarsal bone structure|metatarsal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7675,7681|false|false|false|C5889824||status
Finding|Idea or Concept|SIMPLE_SEGMENT|7675,7681|false|false|false|C1546481|What subject filter - Status|status
Finding|Gene or Genome|SIMPLE_SEGMENT|7682,7686|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|7687,7697|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|7687,7697|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7687,7697|false|false|false|C0002688|Amputation|amputation
Drug|Organic Chemical|SIMPLE_SEGMENT|7711,7714|false|false|false|C0065610|maltose tetrapalmitate|MTP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7711,7714|false|false|false|C0065610|maltose tetrapalmitate|MTP
Finding|Gene or Genome|SIMPLE_SEGMENT|7711,7714|false|false|false|C1826328;C3890208|MTTP gene;MTTP wt Allele|MTP
Finding|Functional Concept|SIMPLE_SEGMENT|7733,7740|false|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|7752,7760|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|7752,7760|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body System|SIMPLE_SEGMENT|7773,7777|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7773,7777|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7773,7777|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|7773,7777|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|7773,7777|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|SIMPLE_SEGMENT|7773,7783|false|false|false|C0521464|Edematous skin|skin edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7778,7783|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7778,7783|false|false|false|C0013604|Edema|edema
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7786,7789|false|false|false|C0039985|Plain chest X-ray|CXR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7790,7794|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7790,7804|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC PLACEMENT
Procedure|Health Care Activity|SIMPLE_SEGMENT|7795,7804|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|PLACEMENT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7795,7804|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|PLACEMENT
Finding|Intellectual Product|SIMPLE_SEGMENT|7811,7821|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|7811,7821|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|SIMPLE_SEGMENT|7826,7829|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|7826,7829|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Functional Concept|SIMPLE_SEGMENT|7830,7835|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7836,7840|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Finding|Gene or Genome|SIMPLE_SEGMENT|7846,7849|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7846,7849|false|false|false|C0673828|TIP regimen|tip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7887,7905|false|false|false|C0042459;C4266604|Chest>Vena cava.superior;Superior vena cava structure|superior vena cava
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7896,7900|false|false|false|C0447122|Structure of vein of trunk|vena
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7896,7905|false|false|false|C0042460;C4266402|Chest+Abdomen>Vena cava.superior &or Vena cava.inferior;Vena caval structure|vena cava
Finding|Gene or Genome|SIMPLE_SEGMENT|7901,7905|false|false|false|C1413046|CA5A gene|cava
Finding|Functional Concept|SIMPLE_SEGMENT|7910,7915|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7910,7922|false|false|false|C0225844|Right atrial structure|right atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7916,7922|false|false|false|C0018792|Heart Atrium|atrium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7928,7940|true|false|false|C0032326|Pneumothorax|pneumothorax
Finding|Idea or Concept|SIMPLE_SEGMENT|7943,7948|false|false|false|C1550016|Remote control command - Clear|Clear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7949,7954|false|false|false|C0024109|Lung|lungs
Finding|Functional Concept|SIMPLE_SEGMENT|7957,7966|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|PATHOLOGY
Finding|Pathologic Function|SIMPLE_SEGMENT|7957,7966|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|PATHOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7957,7966|false|false|false|C0919386|Pathology procedure|PATHOLOGY
Procedure|Health Care Activity|SIMPLE_SEGMENT|7978,7986|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|SURGICAL
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7978,7986|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|SURGICAL
Anatomy|Tissue|SIMPLE_SEGMENT|7987,7993|false|false|false|C0040300|Body tissue|TISSUE
Finding|Intellectual Product|SIMPLE_SEGMENT|7987,7993|false|false|false|C1547928|Tissue Specimen Code|TISSUE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8002,8006|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|Bone
Finding|Body Substance|SIMPLE_SEGMENT|8002,8006|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Intellectual Product|SIMPLE_SEGMENT|8002,8006|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Functional Concept|SIMPLE_SEGMENT|8023,8030|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|8032,8042|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|8032,8047|false|false|false|C0332290|Consistent with|consistent with
Finding|Intellectual Product|SIMPLE_SEGMENT|8048,8055|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|8048,8055|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8057,8070|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Idea or Concept|SIMPLE_SEGMENT|8086,8094|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8086,8097|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|SIMPLE_SEGMENT|8098,8103|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8098,8117|true|false|false|C0158371|Acute osteomyelitis|acute osteomyelitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8104,8117|true|false|false|C0029443|Osteomyelitis|osteomyelitis
Procedure|Health Care Activity|SIMPLE_SEGMENT|8121,8129|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|SURGICAL
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8121,8129|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|SURGICAL
Anatomy|Tissue|SIMPLE_SEGMENT|8130,8136|false|false|false|C0040300|Body tissue|TISSUE
Finding|Intellectual Product|SIMPLE_SEGMENT|8130,8136|false|false|false|C1547928|Tissue Specimen Code|TISSUE
Finding|Functional Concept|SIMPLE_SEGMENT|8146,8150|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Finding|Gene or Genome|SIMPLE_SEGMENT|8151,8156|false|false|false|C1424898|RXFP2 gene|GREAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8151,8160|false|false|false|C0018534|Hallux structure|GREAT TOE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8157,8160|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|TOE
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8162,8170|false|false|false|C0015252;C0728940|Excision;removal technique|EXCISION
Finding|Intellectual Product|SIMPLE_SEGMENT|8174,8179|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8174,8193|false|false|false|C0158371|Acute osteomyelitis|Acute osteomyelitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8180,8193|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8204,8208|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|Bone
Finding|Body Substance|SIMPLE_SEGMENT|8204,8208|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Intellectual Product|SIMPLE_SEGMENT|8204,8208|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Functional Concept|SIMPLE_SEGMENT|8225,8232|false|false|false|C0392747|Changing|changes
Anatomy|Body System|SIMPLE_SEGMENT|8236,8240|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8236,8240|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8236,8240|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|8236,8240|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|8236,8240|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Anatomy|Tissue|SIMPLE_SEGMENT|8245,8253|false|false|false|C0222331;C0278403|Subcutaneous Fat;Subcutaneous Tissue|subcutis
Finding|Pathologic Function|SIMPLE_SEGMENT|8259,8269|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Finding|Intellectual Product|SIMPLE_SEGMENT|8274,8279|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|8274,8292|false|false|false|C0333361|Acute inflammation|acute inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|8280,8292|false|false|false|C0021368|Inflammation|inflammation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8296,8311|false|true|false|C0003850;C0004153|Arteriosclerosis;Atherosclerosis|Atherosclerosis
Finding|Finding|SIMPLE_SEGMENT|8313,8319|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8313,8319|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8324,8332|false|false|false|C4489236|Proximal Resection Margin|PROXIMAL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8324,8340|false|false|false|C0576462;C3669035|Bone structure of proximal phalanx|PROXIMAL PHALANX
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8333,8340|false|false|false|C0222682;C0223792|Phalanx of hand;Phalanx structure|PHALANX
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8341,8345|false|false|false|C2987514|Anatomical base|BASE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8341,8345|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|8341,8345|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|8341,8345|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Finding|Gene or Genome|SIMPLE_SEGMENT|8341,8345|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Finding|Idea or Concept|SIMPLE_SEGMENT|8341,8345|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Finding|Finding|SIMPLE_SEGMENT|8346,8352|false|false|false|C4761388||MARGIN
Finding|Functional Concept|SIMPLE_SEGMENT|8354,8358|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8360,8368|false|false|false|C0015252;C0728940|Excision;removal technique|EXCISION
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8372,8376|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|Bone
Finding|Body Substance|SIMPLE_SEGMENT|8372,8376|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Intellectual Product|SIMPLE_SEGMENT|8372,8376|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Functional Concept|SIMPLE_SEGMENT|8393,8400|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|8416,8424|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8416,8427|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|SIMPLE_SEGMENT|8428,8433|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8428,8447|true|false|false|C0158371|Acute osteomyelitis|acute osteomyelitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8434,8447|true|false|false|C0029443|Osteomyelitis|osteomyelitis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8452,8460|false|false|false|C4489236|Proximal Resection Margin|PROXIMAL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8452,8468|false|false|false|C0576462;C3669035|Bone structure of proximal phalanx|PROXIMAL PHALANX
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8461,8468|false|false|false|C0222682;C0223792|Phalanx of hand;Phalanx structure|PHALANX
Finding|Functional Concept|SIMPLE_SEGMENT|8470,8474|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8476,8484|false|false|false|C0015252;C0728940|Excision;removal technique|EXCISION
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8488,8492|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|Bone
Finding|Body Substance|SIMPLE_SEGMENT|8488,8492|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Intellectual Product|SIMPLE_SEGMENT|8488,8492|false|false|false|C1546560;C1550616|Specimen Type - Bone|Bone
Finding|Functional Concept|SIMPLE_SEGMENT|8509,8516|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|8532,8540|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8532,8543|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|SIMPLE_SEGMENT|8544,8549|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8544,8563|true|false|false|C0158371|Acute osteomyelitis|acute osteomyelitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8550,8563|true|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Functional Concept|SIMPLE_SEGMENT|8566,8578|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|8566,8578|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8566,8578|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Anatomy|Tissue|SIMPLE_SEGMENT|8605,8611|false|false|false|C0040300|Body tissue|TISSUE
Finding|Intellectual Product|SIMPLE_SEGMENT|8605,8611|false|false|false|C1547928|Tissue Specimen Code|TISSUE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8617,8625|false|false|false|C4489236|Proximal Resection Margin|PROXIMAL
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8640,8650|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8640,8650|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8640,8650|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8645,8650|false|false|false|C0038128|Stains|STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8645,8650|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|8652,8657|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Conceptual Entity|SIMPLE_SEGMENT|8689,8694|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|8689,8694|false|false|false|C1553496|field - patient encounter|FIELD
Anatomy|Cell|SIMPLE_SEGMENT|8718,8728|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|8718,8728|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|8718,8728|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Conceptual Entity|SIMPLE_SEGMENT|8756,8761|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|8756,8761|false|false|false|C1553496|field - patient encounter|FIELD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|8771,8779|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Finding|Classification|SIMPLE_SEGMENT|8771,8779|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|SIMPLE_SEGMENT|8771,8779|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Anatomy|Tissue|SIMPLE_SEGMENT|8873,8879|false|false|false|C0040300|Body tissue|TISSUE
Finding|Intellectual Product|SIMPLE_SEGMENT|8873,8879|false|false|false|C1547928|Tissue Specimen Code|TISSUE
Finding|Idea or Concept|SIMPLE_SEGMENT|8881,8886|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8899,8904|false|false|false|C0038160|Staphylococcal Infections|STAPH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8912,8916|false|false|false|C0005790|Blood coagulation tests|COAG
Finding|Finding|SIMPLE_SEGMENT|8930,8936|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8930,8936|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|8930,8936|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|8930,8936|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8930,8936|false|false|false|C2911660|Growth action|GROWTH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8948,8962|false|false|false|C0012655|Disease susceptibility|Susceptibility
Finding|Functional Concept|SIMPLE_SEGMENT|8948,8962|false|false|false|C1264642|Susceptibility (property) (qualifier value)|Susceptibility
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8948,8970|false|false|false|C0806957|Microbial susceptibility tests|Susceptibility testing
Finding|Functional Concept|SIMPLE_SEGMENT|8963,8970|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|SIMPLE_SEGMENT|8963,8970|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8984,8991|false|false|false|C1706355|Culture Dose Form|culture
Finding|Functional Concept|SIMPLE_SEGMENT|8984,8991|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|8984,8991|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8984,8991|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9009,9026|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9019,9026|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9019,9026|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9019,9026|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9019,9026|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9028,9033|false|false|false|C1546485|Diagnosis Type - Final|Final
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9071,9080|false|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|SIMPLE_SEGMENT|9076,9080|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|9076,9080|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|9076,9080|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Activity|SIMPLE_SEGMENT|9081,9086|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|9081,9086|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9081,9086|false|false|false|C0444186|Smear test|SMEAR
Finding|Idea or Concept|SIMPLE_SEGMENT|9088,9093|false|false|false|C1546485|Diagnosis Type - Final|Final
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9109,9118|true|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|SIMPLE_SEGMENT|9114,9118|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|9114,9118|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|9114,9118|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Intellectual Product|SIMPLE_SEGMENT|9135,9141|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Event|Activity|SIMPLE_SEGMENT|9142,9147|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|9142,9147|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9142,9147|false|false|false|C0444186|Smear test|SMEAR
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9154,9163|false|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|SIMPLE_SEGMENT|9159,9163|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|9159,9163|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|9159,9163|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9164,9171|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9164,9171|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9164,9171|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9164,9171|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9259,9264|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|9259,9264|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9259,9272|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9265,9272|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9265,9272|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9265,9272|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9265,9272|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9304,9309|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|9304,9316|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9310,9316|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|9310,9316|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|9310,9316|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9325,9330|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|9325,9330|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9325,9338|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9331,9338|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|9331,9338|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9331,9338|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9331,9338|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9340,9347|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|9340,9347|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9340,9347|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|9349,9354|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|9366,9372|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9366,9372|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|9366,9372|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|9366,9372|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9366,9372|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9446,9451|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|9446,9451|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9446,9459|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9452,9459|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9452,9459|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9452,9459|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9452,9459|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9491,9496|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|9491,9503|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9497,9503|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|9497,9503|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|9497,9503|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9512,9517|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|9512,9517|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9512,9525|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9518,9525|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|9518,9525|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9518,9525|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9518,9525|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9527,9534|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|9527,9534|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9527,9534|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|9536,9541|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|9553,9559|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9553,9559|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|9553,9559|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|9553,9559|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9553,9559|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9634,9639|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|9634,9639|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9634,9647|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9640,9647|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9640,9647|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9640,9647|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9640,9647|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9679,9684|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|9679,9691|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9685,9691|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|9685,9691|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|9685,9691|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9700,9705|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|9700,9705|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9700,9713|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9706,9713|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|9706,9713|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9706,9713|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9706,9713|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9715,9722|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|9715,9722|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9715,9722|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|9724,9729|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|9741,9747|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9741,9747|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|9741,9747|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|9741,9747|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9741,9747|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9822,9827|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|9822,9827|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9822,9835|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9828,9835|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|9828,9835|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9828,9835|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9828,9835|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|9867,9872|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|9867,9879|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9873,9879|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|9873,9879|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|9873,9879|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9888,9893|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|9888,9893|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9888,9901|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9894,9901|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|9894,9901|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9894,9901|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9894,9901|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|9903,9910|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|9903,9910|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9903,9910|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|9912,9917|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|9929,9935|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9929,9935|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|9929,9935|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|9929,9935|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9929,9935|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10010,10015|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|10010,10015|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10010,10023|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10016,10023|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|10016,10023|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|10016,10023|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10016,10023|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|10055,10060|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|10055,10067|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10061,10067|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|10061,10067|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|10061,10067|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10076,10081|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|10076,10081|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10076,10089|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10082,10089|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|10082,10089|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|10082,10089|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10082,10089|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|10091,10098|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|10091,10098|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10091,10098|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|10100,10105|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|10117,10123|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10117,10123|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|10117,10123|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|10117,10123|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10117,10123|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10198,10203|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|10198,10203|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10198,10211|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10204,10211|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|10204,10211|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|10204,10211|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10204,10211|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|10243,10248|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|10243,10255|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10249,10255|false|false|false|C4255046||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|10249,10255|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|10249,10255|false|false|false|C0700287|Reporting|REPORT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10264,10269|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|10264,10269|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10264,10277|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10270,10277|false|false|false|C1706355|Culture Dose Form|Culture
Finding|Functional Concept|SIMPLE_SEGMENT|10270,10277|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|10270,10277|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10270,10277|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|SIMPLE_SEGMENT|10279,10286|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|10279,10286|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10279,10286|false|false|false|C1979801|Routine coag|Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|10288,10293|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|10305,10311|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10305,10311|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|10305,10311|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|10305,10311|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10305,10311|true|false|false|C2911660|Growth action|GROWTH
Finding|Intellectual Product|SIMPLE_SEGMENT|10317,10322|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|10323,10331|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10323,10338|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|10323,10338|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Intellectual Product|SIMPLE_SEGMENT|10354,10361|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10403,10406|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Finding|SIMPLE_SEGMENT|10426,10434|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10426,10439|false|false|false|C0206172|Diabetic Foot|diabetic foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10435,10439|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|10435,10439|false|false|false|C0555980|Foot problem|foot
Finding|Body Substance|SIMPLE_SEGMENT|10441,10446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|10441,10446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|10441,10446|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Functional Concept|SIMPLE_SEGMENT|10454,10458|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10459,10465|false|false|false|C0018534|Hallux structure|hallux
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10481,10494|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Procedure|Health Care Activity|SIMPLE_SEGMENT|10511,10519|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10511,10519|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10520,10531|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Finding|Idea or Concept|SIMPLE_SEGMENT|10536,10543|false|false|false|C1550516|Target Awareness - partial|partial
Anatomy|Tissue|SIMPLE_SEGMENT|10544,10550|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|10544,10550|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10555,10559|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|10555,10559|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|10555,10559|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Event|Activity|SIMPLE_SEGMENT|10561,10568|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10561,10568|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10589,10598|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10589,10598|false|false|false|C3714514|Infection|infection
Finding|Functional Concept|SIMPLE_SEGMENT|10629,10633|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10634,10640|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|10641,10651|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|10641,10651|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10641,10651|false|false|false|C0002688|Amputation|amputation
Finding|Finding|SIMPLE_SEGMENT|10677,10682|false|false|false|C3714655|On IV|on IV
Drug|Antibiotic|SIMPLE_SEGMENT|10683,10692|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|10683,10692|false|false|false|C0027324|nafcillin|nafcillin
Finding|Finding|SIMPLE_SEGMENT|10697,10701|false|false|false|C2355591|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|MSSA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10702,10711|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10702,10711|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10717,10721|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|SIMPLE_SEGMENT|10717,10721|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|10717,10721|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|10717,10721|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Idea or Concept|SIMPLE_SEGMENT|10725,10733|false|false|false|C0549178|Continuous|continue
Finding|Idea or Concept|SIMPLE_SEGMENT|10734,10738|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10734,10738|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10734,10738|false|false|false|C1553498|home health encounter|home
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10740,10749|false|false|false|C0574032|Infusion procedures|infusions
Drug|Antibiotic|SIMPLE_SEGMENT|10753,10762|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|10753,10762|false|false|false|C0027324|nafcillin|nafcillin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10812,10825|false|false|false|C0029443|Osteomyelitis|Osteomyelitis
Finding|Functional Concept|SIMPLE_SEGMENT|10829,10833|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10834,10840|false|false|false|C0018534|Hallux structure|hallux
Finding|Finding|SIMPLE_SEGMENT|10849,10857|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10849,10863|false|false|false|C1299632|Skin ulcer due to diabetes mellitus|diabetic ulcer
Finding|Body Substance|SIMPLE_SEGMENT|10858,10863|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|10858,10863|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|10858,10863|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Functional Concept|SIMPLE_SEGMENT|10867,10871|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10873,10879|false|false|false|C0018534|Hallux structure|hallux
Finding|Body Substance|SIMPLE_SEGMENT|10881,10888|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10881,10888|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10881,10888|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10899,10906|false|false|false|C1550516|Target Awareness - partial|partial
Finding|Functional Concept|SIMPLE_SEGMENT|10907,10911|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10912,10918|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|10919,10929|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|10919,10929|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10919,10929|false|false|false|C0002688|Amputation|amputation
Finding|Finding|SIMPLE_SEGMENT|10976,10981|false|false|false|C3714655|On IV|on IV
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10982,10992|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|10982,10992|false|false|false|C0042313|vancomycin|Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10982,10992|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Organic Chemical|SIMPLE_SEGMENT|10994,11000|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10994,11000|false|false|false|C0699678|Flagyl|Flagyl
Drug|Antibiotic|SIMPLE_SEGMENT|11007,11015|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|11007,11015|false|false|false|C0055003|cefepime|cefepime
Finding|Idea or Concept|SIMPLE_SEGMENT|11017,11024|false|false|false|C1555582|Initial (abbreviation)|Initial
Procedure|Health Care Activity|SIMPLE_SEGMENT|11025,11033|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11025,11033|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Finding|Idea or Concept|SIMPLE_SEGMENT|11034,11042|false|false|false|C0010453|Culture (Anthropological)|cultures
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|11053,11061|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|SIMPLE_SEGMENT|11053,11061|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|11053,11061|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|11053,11065|false|false|false|C1446409|Positive|positive for
Finding|Finding|SIMPLE_SEGMENT|11067,11071|false|false|false|C2355591|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|MSSA
Drug|Antibiotic|SIMPLE_SEGMENT|11094,11103|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|11094,11103|false|false|false|C0027324|nafcillin|nafcillin
Finding|Body Substance|SIMPLE_SEGMENT|11105,11112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11105,11112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11105,11112|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|11130,11138|false|false|false|C0277797|Apyrexial|afebrile
Finding|Functional Concept|SIMPLE_SEGMENT|11148,11152|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11148,11157|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11153,11157|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|11153,11157|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11176,11184|false|false|false|C0041834|Erythema|erythema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11186,11191|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|11186,11191|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11194,11198|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11194,11198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11194,11198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|11208,11213|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|11208,11213|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|11208,11213|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Finding|SIMPLE_SEGMENT|11230,11234|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|SIMPLE_SEGMENT|11246,11253|false|false|false|C2699424|Concern|concern
Finding|Intellectual Product|SIMPLE_SEGMENT|11259,11263|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11264,11272|false|false|false|C0003842|Arteries|arterial
Anatomy|Tissue|SIMPLE_SEGMENT|11264,11278|false|false|false|C2335890|Portion of arterial blood|arterial blood
Finding|Body Substance|SIMPLE_SEGMENT|11264,11278|false|false|false|C0229665;C1550611|Arterial blood;Specimen Type - Blood arterial|arterial blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11273,11278|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|11273,11278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Physiologic Function|SIMPLE_SEGMENT|11273,11283|false|false|false|C0005775;C0232338|Blood Circulation;Blood flow|blood flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11279,11283|false|false|false|C0806140|Flow|flow
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11321,11329|false|false|false|C0003842|Arteries|arterial
Procedure|Research Activity|SIMPLE_SEGMENT|11330,11337|false|false|false|C0947630|Scientific Study|studies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11351,11356|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|11351,11356|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11351,11368|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11357,11368|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Research Activity|SIMPLE_SEGMENT|11374,11381|false|false|false|C0947630|Scientific Study|studies
Finding|Intellectual Product|SIMPLE_SEGMENT|11390,11394|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|11395,11410|false|false|false|C0333482|atherosclerotic|atherosclerotic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11411,11418|false|false|false|C0012634|Disease|disease
Finding|Functional Concept|SIMPLE_SEGMENT|11426,11430|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11426,11434|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11431,11434|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11439,11443|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|11439,11443|false|false|false|C0555980|Foot problem|foot
Finding|Finding|SIMPLE_SEGMENT|11450,11456|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11450,11456|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|SIMPLE_SEGMENT|11457,11472|false|false|false|C0333482|atherosclerotic|atherosclerotic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11473,11480|false|false|false|C0012634|Disease|disease
Finding|Functional Concept|SIMPLE_SEGMENT|11488,11493|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11488,11497|false|false|false|C0230415;C0230442|Right lower extremity;Structure of right lower leg|right leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11494,11497|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11502,11506|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|11502,11506|false|false|false|C0555980|Foot problem|foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11509,11517|false|false|false|C0005847|Blood Vessel|Vascular
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11509,11525|false|false|false|C0042381|Vascular Surgical Procedures|Vascular surgery
Finding|Finding|SIMPLE_SEGMENT|11518,11525|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|11518,11525|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|11518,11525|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11518,11525|false|false|false|C0543467|Operative Surgical Procedures|surgery
Procedure|Health Care Activity|SIMPLE_SEGMENT|11554,11566|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11554,11566|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11599,11607|false|false|false|C0005847|Blood Vessel|vascular
Procedure|Health Care Activity|SIMPLE_SEGMENT|11608,11620|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11608,11620|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Finding|SIMPLE_SEGMENT|11655,11662|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|11655,11662|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|11655,11662|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11655,11662|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Body Substance|SIMPLE_SEGMENT|11668,11675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11668,11675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11668,11675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|11733,11737|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11738,11744|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|11745,11755|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|11745,11755|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11745,11755|false|false|false|C0002688|Amputation|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|11771,11779|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Finding|Conceptual Entity|SIMPLE_SEGMENT|11780,11791|false|false|false|C2986411|Improvement|improvement
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11801,11806|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|11801,11806|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|SIMPLE_SEGMENT|11801,11811|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11801,11817|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|SIMPLE_SEGMENT|11807,11811|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|11807,11811|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11807,11817|false|false|false|C0007584|Cell Count|cell count
Finding|Functional Concept|SIMPLE_SEGMENT|11848,11857|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|11848,11857|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11848,11857|false|false|false|C0919386|Pathology procedure|pathology
Finding|Intellectual Product|SIMPLE_SEGMENT|11848,11864|false|false|false|C0807321|Pathology report|pathology report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11858,11864|false|false|false|C4255046||report
Finding|Intellectual Product|SIMPLE_SEGMENT|11858,11864|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|11858,11864|false|false|false|C0700287|Reporting|report
Event|Activity|SIMPLE_SEGMENT|11872,11877|false|false|false|C1947930|Cleaning (activity)|clean
Finding|Body Substance|SIMPLE_SEGMENT|11897,11904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11897,11904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11897,11904|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11923,11932|false|false|false|C2984058|Have Pain|have pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11928,11932|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11928,11932|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11928,11932|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11959,11967|false|false|false|C0041834|Erythema|erythema
Finding|Finding|SIMPLE_SEGMENT|11972,11980|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|11972,11980|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Procedure|Health Care Activity|SIMPLE_SEGMENT|11988,11996|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11988,11996|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11997,12001|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|11997,12001|false|false|false|C1546778||site
Finding|Gene or Genome|SIMPLE_SEGMENT|12006,12009|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12006,12009|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|12006,12009|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Functional Concept|SIMPLE_SEGMENT|12018,12022|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12018,12027|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12023,12027|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|12023,12027|false|false|false|C0555980|Foot problem|foot
Procedure|Health Care Activity|SIMPLE_SEGMENT|12074,12082|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12074,12082|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12074,12087|false|false|false|C0038925|Surgical Flaps|surgical flap
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12083,12087|false|false|false|C0038925|Surgical Flaps|flap
Finding|Gene or Genome|SIMPLE_SEGMENT|12083,12087|false|false|false|C1412362|ALOX5AP gene|flap
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12094,12099|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|12094,12099|false|false|false|C0013604|Edema|edema
Finding|Conceptual Entity|SIMPLE_SEGMENT|12126,12130|false|false|false|C1427618;C1705203|Spot (mark);THEMIS gene|spot
Finding|Gene or Genome|SIMPLE_SEGMENT|12126,12130|false|false|false|C1427618;C1705203|Spot (mark);THEMIS gene|spot
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12139,12143|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|12139,12143|false|false|false|C1546778||site
Finding|Finding|SIMPLE_SEGMENT|12151,12158|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|12151,12158|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|12151,12158|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12151,12158|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|SIMPLE_SEGMENT|12174,12179|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|12174,12179|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12183,12190|true|false|false|C0000833|Abscess|abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|12183,12190|true|false|false|C1546533||abscess
Drug|Substance|SIMPLE_SEGMENT|12194,12199|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|12194,12199|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|SIMPLE_SEGMENT|12201,12211|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|12201,12211|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|12201,12211|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|12201,12211|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Body Substance|SIMPLE_SEGMENT|12232,12239|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12232,12239|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12232,12239|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12257,12262|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Procedure|Health Care Activity|SIMPLE_SEGMENT|12264,12272|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12264,12272|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Finding|Finding|SIMPLE_SEGMENT|12264,12285|false|false|false|C0549433|Surgical intervention (finding)|surgical intervention
Procedure|Health Care Activity|SIMPLE_SEGMENT|12273,12285|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12273,12285|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Finding|SIMPLE_SEGMENT|12300,12305|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|12300,12305|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|12306,12312|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|12306,12312|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|12306,12315|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|12306,12315|false|false|false|C1522577|follow-up|follow-up
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12327,12331|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12332,12336|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|12332,12336|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|12332,12336|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|SIMPLE_SEGMENT|12332,12336|false|false|false|C1546701|line source specimen code|line
Finding|Functional Concept|SIMPLE_SEGMENT|12355,12360|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12355,12364|false|false|false|C0230346;C4048756|Right arm;Right upper arm structure|right arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12361,12364|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|12361,12364|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|12361,12364|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12361,12364|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|12361,12364|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12361,12364|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12385,12389|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|SIMPLE_SEGMENT|12385,12389|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|12385,12389|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|12385,12389|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|12408,12412|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Antibiotic|SIMPLE_SEGMENT|12427,12436|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|12427,12436|false|false|false|C0027324|nafcillin|nafcillin
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|12453,12458|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|12453,12458|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|12453,12458|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|12453,12458|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12487,12495|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|12487,12495|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|12487,12495|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|12487,12495|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12487,12495|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Functional Concept|SIMPLE_SEGMENT|12496,12503|false|false|false|C0392747|Changing|changes
Finding|Functional Concept|SIMPLE_SEGMENT|12507,12511|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12507,12516|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12512,12516|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|12512,12516|false|false|false|C0555980|Foot problem|foot
Procedure|Health Care Activity|SIMPLE_SEGMENT|12517,12525|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12517,12525|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12526,12530|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|12526,12530|false|false|false|C1546778||site
Drug|Organic Chemical|SIMPLE_SEGMENT|12532,12540|false|false|false|C0699524|Betadine|Betadine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12532,12540|false|false|false|C0699524|Betadine|Betadine
Drug|Organic Chemical|SIMPLE_SEGMENT|12584,12589|false|false|false|C3815497|Cough (guaifenesin)|Cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12584,12589|false|false|false|C3815497|Cough (guaifenesin)|Cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|12584,12589|false|false|false|C0010200|Coughing|Cough
Finding|Body Substance|SIMPLE_SEGMENT|12611,12618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12611,12618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12611,12618|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|12629,12634|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12629,12634|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|12629,12634|false|false|false|C0010200|Coughing|cough
Finding|Pathologic Function|SIMPLE_SEGMENT|12688,12699|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Finding|SIMPLE_SEGMENT|12707,12714|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|12707,12714|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|12707,12714|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12707,12714|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|SIMPLE_SEGMENT|12737,12742|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Functional Concept|SIMPLE_SEGMENT|12746,12750|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|12746,12750|false|false|false|C0582103|Medical Examination|exam
Finding|Idea or Concept|SIMPLE_SEGMENT|12757,12762|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Sign or Symptom|SIMPLE_SEGMENT|12769,12777|false|false|false|C0010200|Coughing|coughing
Finding|Functional Concept|SIMPLE_SEGMENT|12781,12787|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12788,12793|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12788,12793|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12788,12799|false|false|false|C0039985|Plain chest X-ray|chest x-ray
Finding|Functional Concept|SIMPLE_SEGMENT|12794,12799|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|SIMPLE_SEGMENT|12794,12799|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|12794,12799|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12794,12799|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Finding|Classification|SIMPLE_SEGMENT|12804,12812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|12804,12812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|12804,12812|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|12804,12816|false|false|false|C0205160|Negative|negative for
Finding|Intellectual Product|SIMPLE_SEGMENT|12821,12826|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12828,12843|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12828,12843|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Event|Activity|SIMPLE_SEGMENT|12861,12871|false|false|false|C1707455|Comparison|comparison
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12884,12889|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12884,12889|false|false|false|C0741025|Chest problem|chest
Finding|Functional Concept|SIMPLE_SEGMENT|12891,12896|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|SIMPLE_SEGMENT|12891,12896|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|12891,12896|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12891,12896|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Finding|Idea or Concept|SIMPLE_SEGMENT|12909,12917|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Functional Concept|SIMPLE_SEGMENT|12937,12944|true|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|12960,12964|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12960,12964|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12960,12964|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|12965,12970|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12965,12970|false|false|false|C0699992|Lasix|Lasix
Finding|Body Substance|SIMPLE_SEGMENT|12974,12983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12974,12983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12974,12983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12974,12983|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12987,12999|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Body Substance|SIMPLE_SEGMENT|13001,13008|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13001,13008|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13001,13008|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13011,13028|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Procedure|Health Care Activity|SIMPLE_SEGMENT|13045,13054|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13070,13075|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|13070,13075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13070,13085|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Finding|Finding|SIMPLE_SEGMENT|13076,13085|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13076,13085|false|false|false|C0033095||pressures
Finding|Finding|SIMPLE_SEGMENT|13091,13094|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|13091,13094|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13100,13108|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13110,13115|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|13110,13115|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13110,13125|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Finding|Finding|SIMPLE_SEGMENT|13116,13125|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13116,13125|false|false|false|C0033095||pressures
Finding|Finding|SIMPLE_SEGMENT|13137,13143|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|13137,13143|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13151,13157|false|true|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Finding|Mental Process|SIMPLE_SEGMENT|13166,13173|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13181,13194|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Finding|SIMPLE_SEGMENT|13204,13212|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13204,13217|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13204,13223|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13213,13217|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|13213,13217|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13213,13223|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|13218,13223|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|13218,13223|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|13218,13223|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13242,13253|false|false|false|C0011079;C3245462|Debridement;Sterile maggot wound debridement|debridement
Finding|Body Substance|SIMPLE_SEGMENT|13255,13262|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13255,13262|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13255,13262|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13265,13270|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|13265,13270|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13265,13280|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Finding|Finding|SIMPLE_SEGMENT|13271,13280|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13271,13280|false|false|false|C0033095||pressures
Finding|Functional Concept|SIMPLE_SEGMENT|13281,13289|false|false|false|C0442805|Increase|increase
Drug|Organic Chemical|SIMPLE_SEGMENT|13324,13332|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13324,13332|false|false|false|C0126174|losartan|losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|13337,13347|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13337,13347|false|false|false|C0016860|furosemide|furosemide
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13362,13367|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|13362,13367|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13362,13376|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|13362,13376|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|13362,13376|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|SIMPLE_SEGMENT|13368,13376|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|13368,13376|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13368,13376|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13368,13376|false|false|false|C0033095||pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13411,13419|false|false|false|C0039155|Systole|systolic
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13429,13439|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|13429,13439|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|13429,13439|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13429,13439|false|false|false|C0201975|Creatinine measurement|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|13481,13489|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13481,13489|false|false|false|C0126174|losartan|losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|13494,13504|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13494,13504|false|false|false|C0016860|furosemide|furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|13510,13520|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13510,13520|false|false|false|C0025859|metoprolol|metoprolol
Finding|Finding|SIMPLE_SEGMENT|13549,13559|false|false|false|C0449381|Observation parameter|parameters
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13586,13594|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13595,13600|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|13595,13600|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13602,13610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|13602,13610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13602,13610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13602,13610|false|false|false|C0033095||pressure
Finding|Finding|SIMPLE_SEGMENT|13664,13676|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Drug|Organic Chemical|SIMPLE_SEGMENT|13704,13712|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13704,13712|false|false|false|C0126174|losartan|losartan
Finding|Idea or Concept|SIMPLE_SEGMENT|13727,13735|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Body Substance|SIMPLE_SEGMENT|13755,13762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13755,13762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13755,13762|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|13778,13783|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13778,13783|false|false|false|C0699992|Lasix|Lasix
Finding|Body Substance|SIMPLE_SEGMENT|13790,13799|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13790,13799|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13790,13799|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13790,13799|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|13809,13817|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|SIMPLE_SEGMENT|13821,13826|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13821,13840|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute Kidney Injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|13821,13840|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute Kidney Injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13827,13833|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13827,13833|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|13827,13833|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13827,13833|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13827,13833|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|13827,13840|false|false|false|C0160420|Injury of kidney|Kidney Injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|13834,13840|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|Injury
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13846,13854|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|13846,13854|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13855,13865|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|13855,13865|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|13855,13865|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13855,13865|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Mental Process|SIMPLE_SEGMENT|13902,13909|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13913,13919|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Drug|Organic Chemical|SIMPLE_SEGMENT|13936,13944|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13936,13944|false|false|false|C0126174|losartan|losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|13950,13960|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13950,13960|false|false|false|C0016860|furosemide|furosemide
Finding|Finding|SIMPLE_SEGMENT|13966,13977|false|false|false|C0020649|Hypotension|hypotension
Drug|Substance|SIMPLE_SEGMENT|13994,14000|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|SIMPLE_SEGMENT|13994,14000|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13994,14000|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Organic Chemical|SIMPLE_SEGMENT|14018,14026|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14018,14026|false|false|false|C0126174|losartan|losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|14031,14041|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14031,14041|false|false|false|C0016860|furosemide|furosemide
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14047,14057|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|14047,14057|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|14047,14057|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14047,14057|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Functional Concept|SIMPLE_SEGMENT|14091,14099|false|false|false|C1879489|Measures (attribute)|measures
Finding|Body Substance|SIMPLE_SEGMENT|14109,14118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14109,14118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14109,14118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14109,14118|false|false|false|C0030685|Patient Discharge|discharge
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14156,14164|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|14156,14164|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Intellectual Product|SIMPLE_SEGMENT|14167,14174|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|14167,14174|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14198,14206|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14198,14215|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14198,14222|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes Mellitus Type 2
Finding|Gene or Genome|SIMPLE_SEGMENT|14216,14220|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|14216,14220|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|14216,14222|false|false|false|C0441730|Type 2|Type 2
Procedure|Health Care Activity|SIMPLE_SEGMENT|14229,14238|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|14229,14247|false|false|false|C0030673|Patient Admission|admission, patient
Finding|Body Substance|SIMPLE_SEGMENT|14240,14247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14240,14247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|14240,14247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14271,14275|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|14271,14275|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|14271,14275|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14276,14283|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|14276,14283|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14276,14283|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|14276,14283|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14276,14283|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14295,14301|false|false|false|C0876064|Lantus|Lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14295,14301|false|false|false|C0876064|Lantus|Lantus
Finding|Idea or Concept|SIMPLE_SEGMENT|14302,14311|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|14302,14311|false|false|false|C1555324|inpatient encounter|inpatient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14340,14347|false|false|false|C0528249|Humalog|Humalog
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14340,14347|false|false|false|C0528249|Humalog|Humalog
Finding|Idea or Concept|SIMPLE_SEGMENT|14348,14357|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|14348,14357|false|false|false|C1555324|inpatient encounter|inpatient
Finding|Finding|SIMPLE_SEGMENT|14376,14383|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14378,14383|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Body Substance|SIMPLE_SEGMENT|14392,14399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14392,14399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|14392,14399|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14402,14407|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|14402,14407|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|14402,14414|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|14408,14414|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14408,14414|false|false|false|C0242209|Sugars|sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14408,14414|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Idea or Concept|SIMPLE_SEGMENT|14451,14460|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|14451,14460|false|false|false|C1555324|inpatient encounter|inpatient
Event|Occupational Activity|SIMPLE_SEGMENT|14462,14469|false|false|false|C0043227|Work|Working
Finding|Idea or Concept|SIMPLE_SEGMENT|14462,14469|false|false|false|C1563351|Diagnosis Type - Working|Working
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14483,14491|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Procedure|Health Care Activity|SIMPLE_SEGMENT|14492,14499|false|false|false|C0009818|Consultation|consult
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14522,14529|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|14522,14529|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14522,14529|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|14522,14529|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14522,14529|false|false|false|C0202098|Insulin measurement|insulin
Finding|Body Substance|SIMPLE_SEGMENT|14580,14587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14580,14587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|14580,14587|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14603,14609|false|false|false|C3892970|Toujeo|Toujeo
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14603,14609|false|false|false|C3892970|Toujeo|Toujeo
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14640,14645|false|false|false|C1998602|Meal (occasion for eating)|meals
Finding|Finding|SIMPLE_SEGMENT|14649,14653|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|14670,14678|false|false|false|C3153996|Tradjenta|Trajenta
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14670,14678|false|false|false|C3153996|Tradjenta|Trajenta
Drug|Organic Chemical|SIMPLE_SEGMENT|14684,14693|false|false|false|C3848669|Jardiance|Jardiance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14684,14693|false|false|false|C3848669|Jardiance|Jardiance
Event|Occupational Activity|SIMPLE_SEGMENT|14697,14701|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|14697,14701|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|SIMPLE_SEGMENT|14697,14708|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14702,14708|false|false|false|C5889824||STATUS
Finding|Idea or Concept|SIMPLE_SEGMENT|14702,14708|false|false|false|C1546481|What subject filter - Status|STATUS
Event|Activity|SIMPLE_SEGMENT|14727,14734|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|14727,14734|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|14727,14734|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|14727,14734|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|14727,14734|false|false|false|C0392367|Physical contact|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|14769,14781|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Body Substance|SIMPLE_SEGMENT|14813,14820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|14813,14820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|14813,14820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|14827,14836|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14827,14836|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14827,14836|false|false|false|C0524222|Oxycodone measurement|oxycodone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14854,14858|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|14854,14858|false|false|false|C0555980|Foot problem|foot
Finding|Sign or Symptom|SIMPLE_SEGMENT|14854,14863|false|false|false|C0016512;C2016948|Foot pain;soft tissue pain in foot|foot pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14859,14863|false|true|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|14859,14863|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|14859,14863|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|14874,14881|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|14874,14881|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|14874,14881|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14874,14881|false|false|false|C0543467|Operative Surgical Procedures|surgery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14922,14925|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14922,14925|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14922,14925|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14922,14925|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|14922,14925|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|14922,14925|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|14922,14925|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14922,14925|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|14922,14925|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|14922,14925|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Activity|SIMPLE_SEGMENT|14926,14937|false|false|false|C0003629|Appointments|appointment
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14971,14975|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|14971,14975|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|14971,14975|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14971,14986|false|false|false|C0002766|Pain management (procedure)|pain management
Event|Occupational Activity|SIMPLE_SEGMENT|14976,14986|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|14976,14986|false|false|false|C0376636|Disease Management|management
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14993,15006|false|false|false|C0029443|Osteomyelitis|Osteomyelitis
Finding|Finding|SIMPLE_SEGMENT|15008,15016|false|false|false|C0439663|Infected|infected
Finding|Finding|SIMPLE_SEGMENT|15017,15025|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15017,15030|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15017,15036|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15026,15030|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|15026,15030|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15026,15036|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|15031,15036|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|15031,15036|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|15031,15036|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Procedure|Health Care Activity|SIMPLE_SEGMENT|15038,15046|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15038,15046|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15038,15053|false|false|false|C0229985|Surgical margins|Surgical margin
Finding|Finding|SIMPLE_SEGMENT|15047,15053|false|false|false|C4761388||margin
Finding|Functional Concept|SIMPLE_SEGMENT|15066,15070|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15071,15077|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|15078,15088|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|15078,15088|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15078,15088|false|false|false|C0002688|Amputation|amputation
Finding|Classification|SIMPLE_SEGMENT|15100,15108|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|15100,15108|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|15100,15108|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|15100,15112|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15114,15127|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Finding|Body Substance|SIMPLE_SEGMENT|15129,15136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|15129,15136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|15129,15136|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|15153,15157|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Antibiotic|SIMPLE_SEGMENT|15168,15177|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|15168,15177|false|false|false|C0027324|nafcillin|nafcillin
Finding|Idea or Concept|SIMPLE_SEGMENT|15183,15190|false|false|false|C0549178|Continuous|ongoing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15191,15195|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15191,15202|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|15191,15202|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15191,15212|false|false|false|C0149778|Soft Tissue Infection|soft tissue infection
Anatomy|Tissue|SIMPLE_SEGMENT|15196,15202|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|15196,15202|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15203,15212|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|15203,15212|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|SIMPLE_SEGMENT|15264,15275|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Conceptual Entity|SIMPLE_SEGMENT|15286,15296|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|15286,15296|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Drug|Antibiotic|SIMPLE_SEGMENT|15329,15338|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|15329,15338|false|false|false|C0027324|nafcillin|nafcillin
Finding|Molecular Function|SIMPLE_SEGMENT|15359,15363|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Finding|Intellectual Product|SIMPLE_SEGMENT|15365,15369|false|false|false|C1720092|Once - dosing instruction fragment|Once
Drug|Antibiotic|SIMPLE_SEGMENT|15383,15393|false|false|false|C0003232|Antibiotics|antibiotic
Finding|Functional Concept|SIMPLE_SEGMENT|15411,15416|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15411,15420|false|false|false|C0230346;C4048756|Right arm;Right upper arm structure|right arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15417,15420|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|15417,15420|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|15417,15420|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15417,15420|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|15417,15420|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15417,15420|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15421,15425|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15426,15430|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|15426,15430|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|15426,15430|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|SIMPLE_SEGMENT|15426,15430|false|false|false|C1546701|line source specimen code|line
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|15449,15454|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|15449,15454|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|15449,15454|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|15449,15454|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15482,15490|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|15482,15490|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|15482,15490|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|15482,15490|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15482,15490|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Functional Concept|SIMPLE_SEGMENT|15492,15499|false|false|false|C0392747|Changing|changes
Finding|Functional Concept|SIMPLE_SEGMENT|15503,15507|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15503,15512|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15508,15512|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|15508,15512|false|false|false|C0555980|Foot problem|foot
Procedure|Health Care Activity|SIMPLE_SEGMENT|15513,15521|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15513,15521|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15522,15526|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|15522,15526|false|false|false|C1546778||site
Drug|Organic Chemical|SIMPLE_SEGMENT|15528,15536|false|false|false|C0699524|Betadine|Betadine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15528,15536|false|false|false|C0699524|Betadine|Betadine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15582,15590|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15582,15599|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15582,15606|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes mellitus type 2
Finding|Gene or Genome|SIMPLE_SEGMENT|15600,15604|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|15600,15604|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Classification|SIMPLE_SEGMENT|15600,15606|false|false|false|C0441730|Type 2|type 2
Finding|Body Substance|SIMPLE_SEGMENT|15608,15615|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|15608,15615|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|15608,15615|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15618,15623|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15618,15623|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|15618,15630|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|15624,15630|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15624,15630|false|false|false|C0242209|Sugars|sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15624,15630|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|15680,15688|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15680,15693|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15680,15699|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15689,15693|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|15689,15693|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15689,15699|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|15694,15699|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|15694,15699|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|15694,15699|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15721,15726|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|15721,15726|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|15721,15733|true|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|15727,15733|true|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15727,15733|true|false|false|C0242209|Sugars|sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15727,15733|true|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|15742,15746|true|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|SIMPLE_SEGMENT|15762,15766|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|15762,15766|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|15762,15766|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|15778,15783|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|15778,15783|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|15784,15790|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|15784,15790|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|15784,15793|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|15784,15793|false|false|false|C1522577|follow-up|follow-up
Finding|Finding|SIMPLE_SEGMENT|15810,15818|false|false|false|C0241863|Diabetic|diabetic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15820,15830|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|15820,15830|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15820,15838|false|false|false|C0237125|Medication Regimen|medication regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|15831,15838|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15831,15838|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15881,15887|false|false|false|C3892970|Toujeo|Toujeo
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15881,15887|false|false|false|C3892970|Toujeo|Toujeo
Finding|Idea or Concept|SIMPLE_SEGMENT|15900,15904|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|15900,15904|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|15900,15904|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|15934,15942|false|false|false|C3153996|Tradjenta|Trajenta
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15934,15942|false|false|false|C3153996|Tradjenta|Trajenta
Drug|Organic Chemical|SIMPLE_SEGMENT|15948,15957|false|false|false|C3848669|Jardiance|Jardiance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15948,15957|false|false|false|C3848669|Jardiance|Jardiance
Finding|Finding|SIMPLE_SEGMENT|15963,15968|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|15963,15968|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|15969,15975|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|15969,15975|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|15969,15978|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|15969,15978|false|false|false|C1522577|follow-up|follow-up
Finding|Body Substance|SIMPLE_SEGMENT|16036,16043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16036,16043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|16036,16043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|16046,16050|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|16046,16054|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Drug|Organic Chemical|SIMPLE_SEGMENT|16056,16065|false|false|false|C3848669|Jardiance|Jardiance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16056,16065|false|false|false|C3848669|Jardiance|Jardiance
Finding|Conceptual Entity|SIMPLE_SEGMENT|16072,16079|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|16072,16079|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|16072,16079|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|16072,16082|false|false|false|C0262926|Medical History|history of
Drug|Organic Chemical|SIMPLE_SEGMENT|16103,16108|false|false|false|C3815497|Cough (guaifenesin)|Cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16103,16108|false|false|false|C3815497|Cough (guaifenesin)|Cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|16103,16108|false|false|false|C0010200|Coughing|Cough
Finding|Body Substance|SIMPLE_SEGMENT|16110,16117|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16110,16117|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|16110,16117|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|16143,16148|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16143,16148|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|16143,16148|false|false|false|C0010200|Coughing|cough
Finding|Idea or Concept|SIMPLE_SEGMENT|16159,16167|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|SIMPLE_SEGMENT|16172,16180|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16185,16197|true|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|SIMPLE_SEGMENT|16185,16197|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|16199,16202|true|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|SIMPLE_SEGMENT|16206,16211|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|16206,16211|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Tissue|SIMPLE_SEGMENT|16215,16222|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16215,16222|true|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|16224,16232|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|16224,16232|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|16224,16232|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16236,16249|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Pathologic Function|SIMPLE_SEGMENT|16266,16277|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Organism Function|SIMPLE_SEGMENT|16290,16296|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|SIMPLE_SEGMENT|16290,16296|false|false|false|C2347804|Clinical Trial Period|period
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16303,16307|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|16303,16307|false|false|false|C0555980|Foot problem|foot
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16303,16315|false|false|false|C0188413|Operative procedure on foot|foot surgery
Finding|Finding|SIMPLE_SEGMENT|16308,16315|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|16308,16315|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|16308,16315|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16308,16315|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|16372,16376|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|16372,16376|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|16372,16376|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|16377,16382|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16377,16382|false|false|false|C0699992|Lasix|Lasix
Finding|Classification|SIMPLE_SEGMENT|16386,16396|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|16386,16396|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Intellectual Product|SIMPLE_SEGMENT|16415,16419|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Classification|SIMPLE_SEGMENT|16428,16438|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|16428,16438|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|SIMPLE_SEGMENT|16439,16444|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16439,16444|false|false|false|C0699992|Lasix|Lasix
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16483,16495|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Body Substance|SIMPLE_SEGMENT|16497,16504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16497,16504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|16497,16504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16535,16539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|16535,16539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|16535,16539|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16541,16552|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16541,16552|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|16541,16552|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|SIMPLE_SEGMENT|16571,16580|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|16571,16580|false|false|false|C1555324|inpatient encounter|inpatient
Finding|Pathologic Function|SIMPLE_SEGMENT|16593,16604|false|false|false|C0857353|Hypotensive|hypotensive
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16642,16659|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16680,16685|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|16680,16685|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|16680,16694|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|16680,16694|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|16680,16694|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|SIMPLE_SEGMENT|16686,16694|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|16686,16694|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|16686,16694|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|16686,16694|false|false|false|C0033095||pressure
Finding|Functional Concept|SIMPLE_SEGMENT|16724,16729|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|SIMPLE_SEGMENT|16731,16738|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16731,16738|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Finding|SIMPLE_SEGMENT|16743,16750|false|false|false|C4036057|Too low|too low
Finding|Finding|SIMPLE_SEGMENT|16747,16750|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|16747,16750|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Organic Chemical|SIMPLE_SEGMENT|16776,16786|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16776,16786|false|false|false|C0016860|furosemide|furosemide
Finding|Body Substance|SIMPLE_SEGMENT|16798,16807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|16798,16807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|16798,16807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|16798,16807|false|false|false|C0030685|Patient Discharge|Discharge
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16808,16818|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|16808,16818|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|16808,16818|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|16808,16818|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Body Substance|SIMPLE_SEGMENT|16839,16846|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16839,16846|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|16839,16846|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|16860,16866|false|false|false|C5202796|Intensity and Distress 1|slight
Drug|Biologically Active Substance|SIMPLE_SEGMENT|16875,16885|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|16875,16885|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|16875,16885|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|16875,16885|false|false|false|C0201975|Creatinine measurement|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|16903,16911|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16903,16911|false|false|false|C0126174|losartan|losartan
Finding|Body Substance|SIMPLE_SEGMENT|16921,16928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|16921,16928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|16921,16928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|16940,16944|false|false|false|C0587081|Laboratory test finding|labs
Drug|Antibiotic|SIMPLE_SEGMENT|16961,16971|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16973,16982|false|false|false|C0574032|Infusion procedures|infusions
Drug|Organic Chemical|SIMPLE_SEGMENT|17000,17004|false|false|false|C0246719|risedronate|rise
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17000,17004|false|false|false|C0246719|risedronate|rise
Finding|Intellectual Product|SIMPLE_SEGMENT|17000,17004|false|false|false|C4321377|Relational and Item-Specific Encoding Task|rise
Drug|Antibiotic|SIMPLE_SEGMENT|17020,17029|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|17020,17029|false|false|false|C0027324|nafcillin|nafcillin
Drug|Antibiotic|SIMPLE_SEGMENT|17060,17070|false|false|false|C0003232|Antibiotics|antibiotic
Drug|Antibiotic|SIMPLE_SEGMENT|17074,17083|false|false|false|C0007546|cefazolin|cefazolin
Drug|Organic Chemical|SIMPLE_SEGMENT|17074,17083|false|false|false|C0007546|cefazolin|cefazolin
Event|Occupational Activity|SIMPLE_SEGMENT|17087,17091|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|17087,17091|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|SIMPLE_SEGMENT|17087,17098|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17092,17098|false|false|false|C5889824||STATUS
Finding|Idea or Concept|SIMPLE_SEGMENT|17092,17098|false|false|false|C1546481|What subject filter - Status|STATUS
Event|Activity|SIMPLE_SEGMENT|17117,17124|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|17117,17124|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|17117,17124|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|17117,17124|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|17117,17124|false|false|false|C0392367|Physical contact|CONTACT
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|17180,17187|false|false|false|C1704241|complex (molecular entity)|complex
Finding|Body Substance|SIMPLE_SEGMENT|17188,17197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|17188,17197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|17188,17197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|17188,17197|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17201,17212|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17201,17212|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|17201,17212|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|17201,17225|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|17216,17225|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17244,17254|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|17244,17254|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|17244,17259|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|17255,17259|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|17276,17284|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17276,17284|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|17276,17284|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|17276,17284|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|17276,17284|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|17289,17302|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17289,17302|false|false|false|C2974540|canagliflozin|canagliflozin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|17310,17314|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17310,17314|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|17310,17314|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|17310,17314|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|17325,17338|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17325,17338|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|17358,17361|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17362,17368|false|false|false|C2926611||angina
Finding|Finding|SIMPLE_SEGMENT|17362,17368|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|17362,17368|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Drug|Organic Chemical|SIMPLE_SEGMENT|17373,17383|false|false|false|C0244821|ropinirole|rOPINIRole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17373,17383|false|false|false|C0244821|ropinirole|rOPINIRole
Finding|Sign or Symptom|SIMPLE_SEGMENT|17398,17406|false|false|false|C0085631;C3887611|Agitation;Restlessness|restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17398,17410|false|false|false|C0035258|Restless Legs Syndrome|restless leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17398,17419|false|true|false|C0035258|Restless Legs Syndrome|restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|17407,17410|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|17411,17419|false|false|false|C0039082|Syndrome|syndrome
Drug|Organic Chemical|SIMPLE_SEGMENT|17424,17433|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17424,17433|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|SIMPLE_SEGMENT|17447,17450|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17451,17459|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|17451,17459|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|SIMPLE_SEGMENT|17464,17476|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17464,17476|false|false|false|C0081876|pantoprazole|Pantoprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|17486,17489|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|17486,17489|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|17486,17489|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|17486,17489|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|17494,17504|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17494,17504|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Gene or Genome|SIMPLE_SEGMENT|17519,17522|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Finding|SIMPLE_SEGMENT|17523,17539|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|Neuropathic pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|17523,17539|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|Neuropathic pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17535,17539|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|17535,17539|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|17535,17539|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|17544,17556|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17544,17556|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|17574,17585|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17574,17585|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|17574,17596|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17574,17596|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|17586,17596|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|17614,17617|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|17614,17617|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|17614,17617|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|17614,17617|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|17622,17633|false|false|false|C2746078|linagliptin|linaGLIPtin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17622,17633|false|false|false|C2746078|linagliptin|linaGLIPtin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|17639,17643|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17639,17643|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|17639,17643|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|17639,17643|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|17655,17663|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17655,17663|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|17655,17673|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17655,17673|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|17664,17673|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|17664,17673|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|17664,17673|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|17664,17673|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17664,17673|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|17664,17673|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17664,17673|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|17694,17703|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17694,17703|false|false|false|C0030049|oxycodone|OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17694,17703|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|17705,17718|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17705,17718|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17705,17718|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17733,17736|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|17744,17747|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17748,17752|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|17748,17752|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|17748,17752|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|17756,17762|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|17756,17762|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Organic Chemical|SIMPLE_SEGMENT|17768,17777|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17768,17777|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17768,17777|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17781,17786|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|SIMPLE_SEGMENT|17781,17786|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|17789,17793|false|false|false|C4308013|PTCH1 protein, human|PTCH
Finding|Gene or Genome|SIMPLE_SEGMENT|17789,17793|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|SIMPLE_SEGMENT|17789,17793|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Drug|Organic Chemical|SIMPLE_SEGMENT|17806,17816|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17806,17816|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|17837,17847|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17837,17847|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|17837,17857|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17837,17857|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|17848,17857|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|17882,17891|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17882,17891|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|17882,17899|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17882,17899|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|17892,17899|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|17892,17899|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17892,17899|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|17917,17927|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|17917,17927|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|SIMPLE_SEGMENT|17932,17935|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|17941,17948|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17941,17948|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|17941,17951|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17941,17951|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Organic Chemical|SIMPLE_SEGMENT|17973,17986|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|17973,17986|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Clinical Drug|SIMPLE_SEGMENT|17973,17994|false|false|false|C0360349||MetronidAZOLE Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17987,17994|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|17987,17994|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|17999,18002|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|17999,18002|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Substance|SIMPLE_SEGMENT|17999,18002|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|17999,18002|false|false|false|C5977403|Blood group antibody screen.GEL|Gel
Finding|Gene or Genome|SIMPLE_SEGMENT|18005,18009|false|false|false|C1858559|APPL1 gene|Appl
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|18019,18026|false|false|false|C0035854|Rosacea|Rosacea
Drug|Antibiotic|SIMPLE_SEGMENT|18032,18040|false|false|false|C0028741|nystatin|nystatin
Drug|Organic Chemical|SIMPLE_SEGMENT|18032,18040|false|false|false|C0028741|nystatin|nystatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18059,18066|false|false|false|C1710439|Topical Dosage Form|topical
Finding|Functional Concept|SIMPLE_SEGMENT|18059,18066|false|false|false|C1522168|Topical Route of Administration|topical
Finding|Gene or Genome|SIMPLE_SEGMENT|18073,18076|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|SIMPLE_SEGMENT|18081,18090|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|18081,18090|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|18081,18090|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|18081,18090|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|18081,18102|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18091,18102|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18091,18102|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|18091,18102|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|18108,18121|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18108,18121|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18108,18121|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|18142,18155|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18142,18155|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18142,18155|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18165,18171|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|18175,18183|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18178,18183|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18178,18183|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|18184,18189|false|false|false|C1720374|Every - dosing instruction fragment|Every
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18203,18207|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|18203,18207|false|false|false|C0555980|Foot problem|foot
Finding|Sign or Symptom|SIMPLE_SEGMENT|18203,18212|false|false|false|C0016512;C2016948|Foot pain;soft tissue pain in foot|foot pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18208,18212|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|18208,18212|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|18208,18212|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18223,18229|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|18230,18237|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|18246,18255|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18246,18255|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|SIMPLE_SEGMENT|18271,18274|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|18275,18287|false|false|false|C0009806|Constipation|Constipation
Finding|Functional Concept|SIMPLE_SEGMENT|18290,18296|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|Second
Finding|Idea or Concept|SIMPLE_SEGMENT|18290,18296|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|Second
Finding|Intellectual Product|SIMPLE_SEGMENT|18290,18296|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|Second
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18297,18301|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|18297,18301|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|18297,18301|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|18297,18301|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|SIMPLE_SEGMENT|18307,18316|false|false|false|C0005632|bisacodyl|bisacodyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18307,18316|false|false|false|C0005632|bisacodyl|bisacodyl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18324,18330|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|18334,18342|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18337,18342|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18337,18342|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|18350,18353|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|18350,18353|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Sign or Symptom|SIMPLE_SEGMENT|18369,18381|false|false|false|C0009806|Constipation|constipation
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18392,18398|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|18399,18406|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|18415,18423|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18415,18423|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|18415,18430|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18415,18430|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18424,18430|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|18424,18430|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18424,18430|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|18424,18430|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18424,18430|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|18441,18444|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|18441,18444|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18441,18444|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|18441,18444|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|18450,18458|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18450,18458|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|18450,18465|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18450,18465|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18459,18465|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|18459,18465|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18459,18465|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|18459,18465|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18459,18465|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18475,18482|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|18475,18482|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18475,18482|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|18486,18494|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18489,18494|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18489,18494|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|18503,18506|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|18503,18506|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18518,18525|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|18518,18525|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18518,18525|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|SIMPLE_SEGMENT|18526,18533|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|SIMPLE_SEGMENT|18542,18551|false|false|false|C0027324|nafcillin|Nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|18542,18551|false|false|false|C0027324|nafcillin|Nafcillin
Drug|Antibiotic|SIMPLE_SEGMENT|18568,18577|false|false|false|C0027324|nafcillin|nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|18568,18577|false|false|false|C0027324|nafcillin|nafcillin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18581,18589|false|false|false|C0017725|glucose|dextrose
Drug|Organic Chemical|SIMPLE_SEGMENT|18581,18589|false|false|false|C0017725|glucose|dextrose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18581,18589|false|false|false|C0017725|glucose|dextrose
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18581,18589|false|false|false|C2034479|intravenous infusion of intravenous dextrose|dextrose
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|18594,18597|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18594,18597|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18594,18597|false|false|false|C0279238;C1702221;C3887694|OSM protein, human;Recombinant Oncostatin M;ovine sialomucin|osm
Finding|Gene or Genome|SIMPLE_SEGMENT|18594,18597|false|false|false|C1335093;C1427709|CCM2 gene;OSM gene|osm
Finding|Intellectual Product|SIMPLE_SEGMENT|18619,18624|false|false|false|C1720374|Every - dosing instruction fragment|Every
Finding|Functional Concept|SIMPLE_SEGMENT|18647,18658|false|false|false|C1522726|Intravenous Route of Administration|Intravenous
Finding|Intellectual Product|SIMPLE_SEGMENT|18659,18662|false|false|false|C1552710|Bag Data Type|Bag
Finding|Idea or Concept|SIMPLE_SEGMENT|18663,18670|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|18679,18688|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18679,18688|false|false|false|C0030049|oxycodone|OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18679,18688|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|SIMPLE_SEGMENT|18690,18699|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|18690,18699|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18690,18707|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Finding|Functional Concept|SIMPLE_SEGMENT|18700,18707|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|18700,18707|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|18700,18707|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|18721,18724|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18725,18729|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|18725,18729|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|18725,18729|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|18733,18741|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|18733,18741|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Organic Chemical|SIMPLE_SEGMENT|18747,18756|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18747,18756|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|18747,18756|false|false|false|C0524222|Oxycodone measurement|oxycodone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18764,18771|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|18764,18771|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18764,18771|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|18775,18783|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18778,18783|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18778,18783|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|SIMPLE_SEGMENT|18818,18824|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|18818,18824|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18825,18829|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|18825,18829|false|false|false|C0555980|Foot problem|foot
Finding|Sign or Symptom|SIMPLE_SEGMENT|18825,18834|false|true|false|C0016512;C2016948|Foot pain;soft tissue pain in foot|foot pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|18830,18834|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|18830,18834|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|18830,18834|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|18846,18853|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|18846,18853|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18846,18853|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|SIMPLE_SEGMENT|18854,18861|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|18870,18875|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18870,18875|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|18886,18889|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|18886,18889|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18886,18889|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|18886,18889|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|18890,18893|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|18894,18906|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|18915,18919|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|18915,18919|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|18915,18919|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|18915,18919|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|SIMPLE_SEGMENT|18925,18935|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18925,18935|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Organic Chemical|SIMPLE_SEGMENT|18937,18942|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|18937,18942|false|false|false|C3489575|sennosides, USP|senna
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|18953,18959|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|18960,18968|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|18963,18968|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|18963,18968|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|18977,18980|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|18977,18980|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Sign or Symptom|SIMPLE_SEGMENT|18996,19008|false|false|false|C0009806|Constipation|constipation
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19019,19025|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|19026,19033|false|false|false|C0807726|refill|Refills
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|19059,19068|false|false|false|C2698559|Breakfast|Breakfast
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|19086,19091|false|false|false|C2697949|Lunch|Lunch
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|19109,19115|false|false|false|C4048877|Dinner|Dinner
Drug|Organic Chemical|SIMPLE_SEGMENT|19121,19130|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19121,19130|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|19121,19138|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19121,19138|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|19131,19138|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|19131,19138|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19131,19138|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|19156,19166|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|19156,19166|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|SIMPLE_SEGMENT|19171,19174|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|19181,19188|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19181,19188|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|19181,19191|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19181,19191|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Organic Chemical|SIMPLE_SEGMENT|19215,19227|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19215,19227|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|19248,19261|false|false|false|C2974540|canagliflozin|canagliflozin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19248,19261|false|false|false|C2974540|canagliflozin|canagliflozin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|19269,19273|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19269,19273|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|19269,19273|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|19269,19273|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|19287,19298|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19287,19298|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|19287,19309|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19287,19309|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|19299,19309|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|19327,19330|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19327,19330|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|19327,19330|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|19327,19330|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|19338,19348|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19338,19348|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|19371,19381|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19371,19381|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Gene or Genome|SIMPLE_SEGMENT|19396,19399|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Finding|SIMPLE_SEGMENT|19400,19416|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|Neuropathic pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|19400,19416|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|Neuropathic pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|19412,19416|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|19412,19416|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|19412,19416|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|19424,19433|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19424,19433|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19424,19433|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19437,19442|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|SIMPLE_SEGMENT|19437,19442|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19445,19449|false|false|false|C4308013|PTCH1 protein, human|PTCH
Finding|Gene or Genome|SIMPLE_SEGMENT|19445,19449|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|SIMPLE_SEGMENT|19445,19449|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Drug|Organic Chemical|SIMPLE_SEGMENT|19464,19475|false|false|false|C2746078|linagliptin|linaGLIPtin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19464,19475|false|false|false|C2746078|linagliptin|linaGLIPtin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|19481,19485|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19481,19485|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|19481,19485|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|19481,19485|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|19499,19507|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19499,19507|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|19499,19517|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19499,19517|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|19508,19517|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|19508,19517|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|19508,19517|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|19508,19517|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19508,19517|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|19508,19517|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19508,19517|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|19540,19550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19540,19550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|19540,19560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19540,19560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|19551,19560|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|19587,19600|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19587,19600|false|false|false|C0025872|metronidazole|MetronidAZOLE
Drug|Clinical Drug|SIMPLE_SEGMENT|19587,19608|false|false|false|C0360349||MetronidAZOLE Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19601,19608|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|SIMPLE_SEGMENT|19601,19608|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19613,19616|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|19613,19616|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Drug|Substance|SIMPLE_SEGMENT|19613,19616|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|Gel
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19613,19616|false|false|false|C5977403|Blood group antibody screen.GEL|Gel
Finding|Gene or Genome|SIMPLE_SEGMENT|19619,19623|false|false|false|C1858559|APPL1 gene|Appl
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|19633,19640|false|false|false|C0035854|Rosacea|Rosacea
Drug|Organic Chemical|SIMPLE_SEGMENT|19648,19661|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19648,19661|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|19681,19684|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|19685,19691|false|false|false|C2926611||angina
Finding|Finding|SIMPLE_SEGMENT|19685,19691|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|19685,19691|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Drug|Antibiotic|SIMPLE_SEGMENT|19699,19707|false|false|false|C0028741|nystatin|nystatin
Drug|Organic Chemical|SIMPLE_SEGMENT|19699,19707|false|false|false|C0028741|nystatin|nystatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19726,19733|false|false|false|C1710439|Topical Dosage Form|topical
Finding|Functional Concept|SIMPLE_SEGMENT|19726,19733|false|false|false|C1522168|Topical Route of Administration|topical
Finding|Gene or Genome|SIMPLE_SEGMENT|19740,19743|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|19751,19760|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19751,19760|false|false|false|C0030049|oxycodone|OxyCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19751,19760|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|19762,19775|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19762,19775|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19762,19775|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|19790,19793|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Gene or Genome|SIMPLE_SEGMENT|19801,19804|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|19805,19809|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|19805,19809|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|19805,19809|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|19813,19819|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|19813,19819|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Organic Chemical|SIMPLE_SEGMENT|19827,19839|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19827,19839|false|false|false|C0081876|pantoprazole|Pantoprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|19849,19852|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19849,19852|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|19849,19852|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|19849,19852|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|19860,19870|false|false|false|C0244821|ropinirole|rOPINIRole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19860,19870|false|false|false|C0244821|ropinirole|rOPINIRole
Finding|Sign or Symptom|SIMPLE_SEGMENT|19885,19893|false|false|false|C0085631;C3887611|Agitation;Restlessness|restless
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|19885,19897|false|false|false|C0035258|Restless Legs Syndrome|restless leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|19885,19906|false|true|false|C0035258|Restless Legs Syndrome|restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|19894,19897|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|19898,19906|false|false|false|C0039082|Syndrome|syndrome
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19933,19940|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|19933,19940|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19933,19940|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|19933,19940|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19933,19940|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19942,19949|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|19942,19949|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19942,19949|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|19942,19949|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|19942,19949|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19942,19958|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Hormone|SIMPLE_SEGMENT|19942,19958|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19942,19958|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|19950,19958|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|19950,19958|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|19950,19958|false|false|false|C0907402|insulin glargine|glargine
Finding|Functional Concept|SIMPLE_SEGMENT|19982,19994|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|SIMPLE_SEGMENT|20022,20031|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|20022,20031|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|SIMPLE_SEGMENT|20045,20048|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|20049,20057|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|20049,20057|false|false|false|C0917801|Sleeplessness|insomnia
Finding|Classification|SIMPLE_SEGMENT|20063,20073|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|20063,20073|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|SIMPLE_SEGMENT|20074,20077|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|SIMPLE_SEGMENT|20074,20077|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Occupational Activity|SIMPLE_SEGMENT|20078,20082|false|false|false|C0043227|Work|Work
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20083,20086|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|20083,20086|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Finding|Gene or Genome|SIMPLE_SEGMENT|20083,20086|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|20083,20086|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|20083,20086|false|false|false|C5575277|Icd Regimen|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|20083,20089|false|false|false|C1137110|International Statistical Classification of Diseases and Related Health Problems, Tenth Revision (ICD-10)|ICD-10
Finding|Gene or Genome|SIMPLE_SEGMENT|20134,20137|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Finding|Intellectual Product|SIMPLE_SEGMENT|20134,20137|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20134,20142|false|false|false|C0022885|Laboratory Procedures|LAB TEST
Anatomy|Body Location or Region|SIMPLE_SEGMENT|20138,20142|false|false|false|C4318744|Test - temporal region|TEST
Finding|Functional Concept|SIMPLE_SEGMENT|20138,20142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Finding|Intellectual Product|SIMPLE_SEGMENT|20138,20142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|20138,20142|false|false|false|C0456984|Test Result|TEST
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20138,20142|false|false|false|C0022885|Laboratory Procedures|TEST
Anatomy|Cell Component|SIMPLE_SEGMENT|20144,20147|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20144,20147|false|false|false|C0009555|Complete Blood Count|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20144,20165|false|false|false|C0545131|complete blood count with differential|CBC with differential
Finding|Idea or Concept|SIMPLE_SEGMENT|20153,20165|false|false|false|C1549478|Amount type - Differential|differential
Drug|Biologically Active Substance|SIMPLE_SEGMENT|20167,20170|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|20167,20170|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20167,20170|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|20176,20179|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|20176,20179|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|20176,20179|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|20176,20179|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|20176,20179|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|SIMPLE_SEGMENT|20176,20179|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|20181,20184|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|20181,20184|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|20181,20184|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|20181,20184|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|20181,20184|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|20181,20184|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|20181,20184|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|20198,20201|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|20198,20201|false|false|false|C1663627|ALK protein, human|ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|20198,20201|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|20198,20201|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|20198,20206|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|20198,20206|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20198,20206|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Finding|Gene or Genome|SIMPLE_SEGMENT|20208,20211|false|false|false|C1414461;C1704489;C1706235|ESR1 gene;ESR1 wt Allele;Extended Rotated Sidebent|ESR
Finding|Pathologic Function|SIMPLE_SEGMENT|20208,20211|false|false|false|C1414461;C1704489;C1706235|ESR1 gene;ESR1 wt Allele;Extended Rotated Sidebent|ESR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|20208,20211|false|false|false|C0013845;C1176468|Electron Spin Resonance Spectroscopy;Erythrocyte sedimentation rate measurement|ESR
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|20213,20216|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|SIMPLE_SEGMENT|20213,20216|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Finding|Gene or Genome|SIMPLE_SEGMENT|20213,20216|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Finding|Idea or Concept|SIMPLE_SEGMENT|20224,20227|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Intellectual Product|SIMPLE_SEGMENT|20224,20227|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Idea or Concept|SIMPLE_SEGMENT|20259,20262|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Intellectual Product|SIMPLE_SEGMENT|20259,20262|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20313,20322|false|false|false|C0945731||DIAGNOSIS
Finding|Classification|SIMPLE_SEGMENT|20313,20322|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|20313,20322|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|20313,20322|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|20324,20328|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|20329,20335|false|false|false|C0018534|Hallux structure|hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|20336,20346|false|false|false|C0332840|Amputated structure (morphologic abnormality)|amputation
Finding|Intellectual Product|SIMPLE_SEGMENT|20336,20346|false|false|false|C1546539|Amputation Specimen Code|amputation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|20336,20346|false|false|false|C0002688|Amputation|amputation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20347,20350|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|20347,20350|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Finding|Gene or Genome|SIMPLE_SEGMENT|20347,20350|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|20347,20350|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|20347,20350|false|false|false|C5575277|Icd Regimen|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|20347,20353|false|false|false|C1137110|International Statistical Classification of Diseases and Related Health Problems, Tenth Revision (ICD-10)|ICD-10
Finding|Idea or Concept|SIMPLE_SEGMENT|20364,20368|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Finding|Body Substance|SIMPLE_SEGMENT|20387,20396|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|20387,20396|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|20387,20396|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|20387,20396|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20387,20408|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|20387,20408|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20397,20408|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|20397,20408|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|20410,20414|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|20410,20414|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|20410,20414|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|20420,20427|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|20420,20427|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|SIMPLE_SEGMENT|20430,20438|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|SIMPLE_SEGMENT|20446,20455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|20446,20455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|20446,20455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|20446,20455|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|20446,20465|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20456,20465|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|20456,20465|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|20456,20465|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|20456,20465|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20467,20484|false|false|false|C0801658||PRIMARY DIAGNOSIS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20475,20484|false|false|false|C0945731||DIAGNOSIS
Finding|Classification|SIMPLE_SEGMENT|20475,20484|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|20475,20484|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|20475,20484|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20503,20516|false|false|false|C0029443|Osteomyelitis|Osteomyelitis
Finding|Functional Concept|SIMPLE_SEGMENT|20520,20524|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|20525,20531|false|false|false|C0018534|Hallux structure|hallux
Disorder|Neoplastic Process|SIMPLE_SEGMENT|20533,20542|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|SIMPLE_SEGMENT|20533,20542|false|false|false|C1522484|metastatic qualifier|SECONDARY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|20543,20552|false|false|false|C0011900|Diagnosis|DIAGNOSES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20573,20585|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Gene or Genome|SIMPLE_SEGMENT|20586,20590|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|20586,20590|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|SIMPLE_SEGMENT|20586,20592|false|false|false|C0441730|Type 2|Type 2
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20586,20601|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20586,20610|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type 2 Diabetes Mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20593,20601|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20593,20610|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Finding|Body Substance|SIMPLE_SEGMENT|20614,20623|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|20614,20623|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|20614,20623|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|20614,20623|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20624,20633|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20624,20633|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|20624,20633|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|20635,20641|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20635,20648|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|20635,20648|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20642,20648|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|20642,20648|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|20650,20655|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|20660,20668|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20670,20692|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|20670,20692|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|20679,20692|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|20679,20692|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20694,20699|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|20694,20699|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|20694,20699|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|20694,20699|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|20694,20699|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|20694,20699|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|20704,20715|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|20717,20725|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|20717,20725|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|20717,20725|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20726,20732|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|20726,20732|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|20734,20744|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|20734,20744|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|20734,20744|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|20734,20744|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|20747,20758|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|20747,20758|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|20763,20772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|20763,20772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|20763,20772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|20763,20772|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20763,20785|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|20763,20785|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|20763,20785|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|20773,20785|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|20773,20785|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|20787,20791|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|SIMPLE_SEGMENT|20811,20819|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|20811,20819|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|20827,20831|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|20827,20831|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|20827,20831|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|20827,20834|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|SIMPLE_SEGMENT|20867,20875|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Finding|SIMPLE_SEGMENT|20887,20895|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20887,20900|false|false|false|C0206172|Diabetic Foot|diabetic foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20887,20906|false|false|false|C1456868|Diabetic foot ulcer|diabetic foot ulcer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|20896,20900|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|20896,20900|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20896,20906|false|false|false|C0085119|Foot Ulcer|foot ulcer
Finding|Body Substance|SIMPLE_SEGMENT|20901,20906|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Intellectual Product|SIMPLE_SEGMENT|20901,20906|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Pathologic Function|SIMPLE_SEGMENT|20901,20906|false|false|false|C0041582;C1547940;C1550672|Specimen Type - Ulcer;Ulcer|ulcer
Finding|Functional Concept|SIMPLE_SEGMENT|20915,20919|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|20920,20923|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Finding|Finding|SIMPLE_SEGMENT|20939,20947|false|false|false|C0439663|Infected|infected
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|20966,20975|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|20966,20975|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|20984,20988|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|20984,20988|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|20984,20988|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Functional Concept|SIMPLE_SEGMENT|21032,21036|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|21037,21040|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|21071,21074|false|false|false|C4522181|Brachial Amyotrophic Diplegia|bad
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|21071,21074|false|false|false|C1530798|BAD protein, human|bad
Drug|Biologically Active Substance|SIMPLE_SEGMENT|21071,21074|false|false|false|C1530798|BAD protein, human|bad
Finding|Gene or Genome|SIMPLE_SEGMENT|21071,21074|false|false|false|C1366450|BAD gene|bad
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|21075,21079|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|21075,21079|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|21075,21079|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|21081,21090|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|21081,21090|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|SIMPLE_SEGMENT|21114,21125|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|21140,21149|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|21140,21149|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|SIMPLE_SEGMENT|21170,21174|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|21170,21174|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|21170,21174|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|21175,21180|false|false|false|C3714655|On IV|on IV
Drug|Antibiotic|SIMPLE_SEGMENT|21181,21192|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Activity|SIMPLE_SEGMENT|21223,21228|false|false|false|C1706081||LEAVE
Finding|Functional Concept|SIMPLE_SEGMENT|21223,21228|false|false|false|C5401409|Leave from Employment|LEAVE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|21259,21270|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|21259,21270|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|21259,21270|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|SIMPLE_SEGMENT|21298,21302|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|21298,21302|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|21298,21302|false|false|false|C1553498|home health encounter|home
Drug|Antibiotic|SIMPLE_SEGMENT|21311,21321|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21311,21330|false|false|false|C0199779|Injection of antibiotic|antibiotic infusion
Finding|Functional Concept|SIMPLE_SEGMENT|21322,21330|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21322,21330|false|false|false|C0574032|Infusion procedures|infusion
Finding|Molecular Function|SIMPLE_SEGMENT|21331,21335|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Procedure|Educational Activity|SIMPLE_SEGMENT|21390,21395|false|false|false|C0039401|Education (procedure)|teach
Drug|Antibiotic|SIMPLE_SEGMENT|21445,21456|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Molecular Function|SIMPLE_SEGMENT|21469,21473|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Finding|Finding|SIMPLE_SEGMENT|21507,21515|false|false|false|C0241863|Diabetic|diabetic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|21516,21526|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|21516,21526|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21516,21534|false|false|false|C0237125|Medication Regimen|medication regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|21527,21534|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21527,21534|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Finding|SIMPLE_SEGMENT|21589,21594|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|21589,21594|false|false|false|C0587267;C3810854|Close;Closed|close
Drug|Organic Chemical|SIMPLE_SEGMENT|21610,21616|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|21610,21616|false|false|false|C0242209|Sugars|sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|21610,21616|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|21617,21624|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|21620,21624|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|21620,21624|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|21620,21624|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|21637,21643|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|21637,21643|false|false|false|C0242209|Sugars|sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|21637,21643|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|21644,21651|false|false|false|C4264481|4 times|4 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|21646,21651|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|21654,21657|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|21654,21657|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|21662,21665|false|false|false|C0228228|lateral occipital gyrus (human only)|log
Finding|Intellectual Product|SIMPLE_SEGMENT|21662,21665|false|false|false|C1708728|Event Log|log
Event|Activity|SIMPLE_SEGMENT|21723,21734|false|false|false|C0003629|Appointments|appointment
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|21783,21793|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|21783,21793|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21783,21801|false|false|false|C0237125|Medication Regimen|medication regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|21794,21801|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21794,21801|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Antibiotic|SIMPLE_SEGMENT|21909,21919|false|false|false|C0003232|Antibiotics|antibiotic
Finding|Intellectual Product|SIMPLE_SEGMENT|21920,21927|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|21920,21927|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Finding|SIMPLE_SEGMENT|22014,22018|false|false|false|C5575035|Well (answer to question)|well
Event|Activity|SIMPLE_SEGMENT|22030,22034|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|22030,22034|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|22030,22034|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|22030,22039|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|22030,22039|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|22042,22050|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|22051,22063|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|22051,22063|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

