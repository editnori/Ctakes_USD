 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
CARDIOTHORACIC|152,166
<EOL>|166,167
<EOL>|168,169
Allergies|169,178
:|178,179
<EOL>|180,181
IV|181,183
Dye|184,187
,|187,188
Iodine|189,195
Containing|196,206
Contrast|207,215
Media|216,221
/|222,223
Oxycodone|224,233
/|234,235
<EOL>|236,237
cilostazol|237,247
/|248,249
Varenicline|250,261
<EOL>|261,262
<EOL>|263,264
Attending|264,273
:|273,274
_|275,276
_|276,277
_|277,278
.|278,279
<EOL>|279,280
<EOL>|281,282
Chief|282,287
Complaint|288,297
:|297,298
<EOL>|298,299
Shortness|299,308
of|309,311
breath|312,318
<EOL>|318,319
<EOL>|320,321
Major|321,326
Surgical|327,335
or|336,338
Invasive|339,347
Procedure|348,357
:|357,358
<EOL>|358,359
Intubation|359,369
&|370,371
Mechanical|372,382
Ventilation|383,394
(|395,396
Extubated|396,405
)|405,406
<EOL>|406,407
Temporary|407,416
Pacer|417,422
Placement|423,432
<EOL>|432,433
CVL|433,436
Insertion|437,446
<EOL>|446,447
<EOL>|447,448
<EOL>|449,450
History|450,457
of|458,460
Present|461,468
Illness|469,476
:|476,477
<EOL>|477,478
_|478,479
_|479,480
_|480,481
with|482,486
COPD|487,491
who|492,495
has|496,499
been|500,504
admitted|505,513
9|514,515
times|516,521
since|522,527
_|528,529
_|529,530
_|530,531
for|532,535
<EOL>|536,537
dyspnea|537,544
,|544,545
CAD|546,549
,|549,550
atrial|551,557
fibrillation|558,570
on|571,573
apixaban|574,582
who|583,586
presented|587,596
with|597,601
<EOL>|602,603
shortness|603,612
of|613,615
breath|616,622
since|623,628
being|629,634
discharged|635,645
on|646,648
_|649,650
_|650,651
_|651,652
.|652,653
She|654,657
was|658,661
<EOL>|662,663
discharged|663,673
home|674,678
with|679,683
services|684,692
.|692,693
<EOL>|695,696
<EOL>|697,698
Mrs.|698,702
_|703,704
_|704,705
_|705,706
has|707,710
significant|711,722
COPD|723,727
,|727,728
with|729,733
recent|734,740
PFTs|741,745
on|746,748
_|749,750
_|750,751
_|751,752
<EOL>|753,754
showing|754,761
severely|762,770
reduced|771,778
FEV1|779,783
and|784,787
moderately|788,798
reduced|799,806
FEV1|807,811
/|811,812
FVC|812,815
.|815,816
<EOL>|817,818
She|818,821
was|822,825
generally|826,835
feeling|836,843
better|844,850
since|851,856
discharged|857,867
on|868,870
_|871,872
_|872,873
_|873,874
,|874,875
<EOL>|876,877
continuing|877,887
her|888,891
prednisone|892,902
(|903,904
at|904,906
40mg|907,911
today|912,917
)|917,918
until|919,924
the|925,928
day|929,932
prior|933,938
to|939,941
<EOL>|942,943
presentation|943,955
.|955,956
She|957,960
subsequently|961,973
began|974,979
to|980,982
become|983,989
short|990,995
of|996,998
breath|999,1005
,|1005,1006
<EOL>|1007,1008
especially|1008,1018
with|1019,1023
exertion|1024,1032
,|1032,1033
and|1034,1037
developed|1038,1047
a|1048,1049
cough|1050,1055
productive|1056,1066
of|1067,1069
<EOL>|1070,1071
brown|1071,1076
sputum|1077,1083
.|1083,1084
No|1085,1087
fever|1088,1093
,|1093,1094
chills|1095,1101
,|1101,1102
nausea|1103,1109
,|1109,1110
vomiting|1111,1119
,|1119,1120
diarrhea|1121,1129
.|1129,1130
She|1131,1134
<EOL>|1135,1136
sleeps|1136,1142
with|1143,1147
three|1148,1153
pillows|1154,1161
laying|1162,1168
on|1169,1171
her|1172,1175
side|1176,1180
,|1180,1181
which|1182,1187
is|1188,1190
stable|1191,1197
.|1197,1198
<EOL>|1199,1200
Her|1200,1203
secondary|1204,1213
concern|1214,1221
is|1222,1224
that|1225,1229
she|1230,1233
is|1234,1236
having|1237,1243
trouble|1244,1251
walking|1252,1259
due|1260,1263
<EOL>|1264,1265
to|1265,1267
pain|1268,1272
in|1273,1275
her|1276,1279
R|1280,1281
-|1281,1282
hip|1282,1285
to|1286,1288
R|1289,1290
-|1290,1291
thigh|1291,1296
with|1297,1301
weight|1302,1308
bearing|1309,1316
.|1316,1317
This|1318,1322
was|1323,1326
<EOL>|1327,1328
new|1328,1331
.|1331,1332
No|1333,1335
falls|1336,1341
or|1342,1344
trauma|1345,1351
.|1351,1352
No|1353,1355
loss|1356,1360
of|1361,1363
sensation|1364,1373
,|1373,1374
numbness|1375,1383
,|1383,1384
<EOL>|1385,1386
weakness|1386,1394
,|1394,1395
urinary|1396,1403
or|1404,1406
fecal|1407,1412
incontinence|1413,1425
or|1426,1428
difficulty|1429,1439
urinating|1440,1449
.|1449,1450
<EOL>|1451,1452
<EOL>|1453,1454
<EOL>|1455,1456
In|1456,1458
the|1459,1462
ED|1463,1465
,|1465,1466
initial|1467,1474
vital|1475,1480
signs|1481,1486
were|1487,1491
:|1491,1492
99.0|1493,1497
80|1498,1500
116|1501,1504
/|1504,1505
66|1505,1507
24|1508,1510
98|1511,1513
%|1513,1514
Nasal|1515,1520
<EOL>|1521,1522
Cannula|1522,1529
<EOL>|1531,1532
-|1533,1534
Exam|1535,1539
was|1540,1543
notable|1544,1551
for|1552,1555
:|1555,1556
diffuse|1557,1564
ronchi|1565,1571
worst|1572,1577
in|1578,1580
the|1581,1584
RLL|1585,1588
,|1588,1589
<EOL>|1590,1591
tripoding|1591,1600
<EOL>|1602,1603
-|1604,1605
Labs|1606,1610
were|1611,1615
notable|1616,1623
for|1624,1627
:|1627,1628
flu|1629,1632
swab|1633,1637
negative|1638,1646
,|1646,1647
WBC|1648,1651
7.5|1652,1655
with|1656,1660
left|1661,1665
<EOL>|1666,1667
shift|1667,1672
,|1672,1673
CBC|1674,1677
otherwise|1678,1687
WNL|1688,1691
,|1691,1692
BNP|1693,1696
425|1697,1700
,|1700,1701
lactate|1702,1709
3.0|1710,1713
,|1713,1714
U|1715,1716
/|1716,1717
A|1717,1718
cloudy|1719,1725
with|1726,1730
<EOL>|1731,1732
30|1732,1734
protein|1735,1742
but|1743,1746
otherwise|1747,1756
negative|1757,1765
,|1765,1766
BUN|1767,1770
/|1770,1771
Cr|1771,1773
_|1774,1775
_|1775,1776
_|1776,1777
<EOL>|1779,1780
-|1781,1782
Imaging|1783,1790
:|1790,1791
CXR|1792,1795
with|1796,1800
mild|1801,1805
bibasilar|1806,1815
atelectasis|1816,1827
,|1827,1828
though|1829,1835
ED|1836,1838
<EOL>|1839,1840
physicians|1840,1850
concerned|1851,1860
for|1861,1864
pneumonia|1865,1874
on|1875,1877
lateral|1878,1885
view|1886,1890
<EOL>|1892,1893
-|1894,1895
The|1896,1899
patient|1900,1907
was|1908,1911
given|1912,1917
:|1917,1918
1g|1919,1921
Vancomycin|1922,1932
,|1932,1933
2g|1934,1936
cefepime|1937,1945
,|1945,1946
500|1947,1950
mg|1951,1953
PO|1954,1956
<EOL>|1957,1958
azithromycin|1958,1970
,|1970,1971
1|1972,1973
duoneb|1974,1980
,|1980,1981
20|1982,1984
mg|1985,1987
prednisone|1988,1998
(|1999,2000
total|2000,2005
60|2006,2008
mg|2009,2011
that|2012,2016
day|2017,2020
)|2020,2021
<EOL>|2023,2024
<EOL>|2024,2025
-|2026,2027
Consults|2028,2036
:|2036,2037
none|2038,2042
<EOL>|2044,2045
Vitals|2046,2052
prior|2053,2058
to|2059,2061
transfer|2062,2070
were|2071,2075
:|2075,2076
98.2|2077,2081
87|2082,2084
148|2085,2088
/|2088,2089
76|2089,2091
18|2092,2094
92|2095,2097
%|2097,2098
RA|2099,2101
<EOL>|2103,2104
<EOL>|2105,2106
Upon|2106,2110
arrival|2111,2118
to|2119,2121
the|2122,2125
floor|2126,2131
,|2131,2132
Mrs.|2133,2137
_|2138,2139
_|2139,2140
_|2140,2141
stated|2142,2148
her|2149,2152
breathing|2153,2162
<EOL>|2163,2164
was|2164,2167
slightly|2168,2176
better|2177,2183
,|2183,2184
but|2185,2188
she|2189,2192
continued|2193,2202
to|2203,2205
have|2206,2210
shortness|2211,2220
of|2221,2223
<EOL>|2224,2225
breath|2225,2231
.|2231,2232
She|2233,2236
felt|2237,2241
as|2242,2244
though|2245,2251
her|2252,2255
ears|2256,2260
are|2261,2264
clogged|2265,2272
up|2273,2275
,|2275,2276
and|2277,2280
this|2281,2285
was|2286,2289
<EOL>|2290,2291
her|2291,2294
as|2295,2297
well|2298,2302
.|2302,2303
She|2304,2307
stated|2308,2314
she|2315,2318
has|2319,2322
been|2323,2327
taking|2328,2334
all|2335,2338
her|2339,2342
medications|2343,2354
<EOL>|2355,2356
as|2356,2358
prescribed|2359,2369
.|2369,2370
<EOL>|2372,2373
<EOL>|2374,2375
Past|2375,2379
Medical|2380,2387
History|2388,2395
:|2395,2396
<EOL>|2396,2397
-|2397,2398
COPD|2399,2403
/|2403,2404
Asthma|2404,2410
on|2411,2413
home|2414,2418
2L|2419,2421
O2|2422,2424
<EOL>|2424,2425
-|2425,2426
Atypical|2427,2435
Chest|2436,2441
Pain|2442,2446
<EOL>|2446,2447
-|2447,2448
Hypertension|2449,2461
<EOL>|2461,2462
-|2462,2463
Hyperlipidemia|2464,2478
<EOL>|2478,2479
-|2479,2480
Osteroarthritis|2481,2496
<EOL>|2496,2497
-|2497,2498
Atrial|2499,2505
Fibrillation|2506,2518
on|2519,2521
Apixaban|2522,2530
<EOL>|2530,2531
-|2531,2532
Anxiety|2533,2540
<EOL>|2540,2541
-|2541,2542
Cervical|2543,2551
Radiculitis|2552,2563
<EOL>|2563,2564
-|2564,2565
Cervical|2566,2574
Spondylosis|2575,2586
<EOL>|2586,2587
-|2587,2588
Coronary|2589,2597
Artery|2598,2604
Disease|2605,2612
<EOL>|2612,2613
-|2613,2614
Headache|2615,2623
<EOL>|2623,2624
-|2624,2625
Herpes|2626,2632
Zoster|2633,2639
<EOL>|2639,2640
-|2640,2641
GI|2642,2644
Bleeding|2645,2653
<EOL>|2653,2654
-|2654,2655
Peripheral|2656,2666
Vascular|2667,2675
Disease|2676,2683
s|2684,2685
/|2685,2686
p|2686,2687
bilateral|2688,2697
iliac|2698,2703
stents|2704,2710
<EOL>|2710,2711
-|2711,2712
s|2713,2714
/|2714,2715
p|2715,2716
hip|2717,2720
replacement|2721,2732
<EOL>|2732,2733
<EOL>|2734,2735
Social|2735,2741
History|2742,2749
:|2749,2750
<EOL>|2750,2751
_|2751,2752
_|2752,2753
_|2753,2754
<EOL>|2754,2755
Family|2755,2761
History|2762,2769
:|2769,2770
<EOL>|2770,2771
Mother|2771,2777
with|2778,2782
asthma|2783,2789
and|2790,2793
hypertension|2794,2806
.|2806,2807
Father|2808,2814
with|2815,2819
colon|2820,2825
cancer|2826,2832
.|2832,2833
<EOL>|2834,2835
Brother|2835,2842
with|2843,2847
leukemia|2848,2856
.|2856,2857
<EOL>|2857,2858
<EOL>|2858,2859
<EOL>|2860,2861
Physical|2861,2869
Exam|2870,2874
:|2874,2875
<EOL>|2875,2876
PHYSICAL|2876,2884
EXAMINATION|2885,2896
ON|2897,2899
ADMISSION|2900,2909
:|2909,2910
<EOL>|2910,2911
=|2911,2912
=|2912,2913
=|2913,2914
=|2914,2915
=|2915,2916
=|2916,2917
=|2917,2918
=|2918,2919
=|2919,2920
=|2920,2921
=|2921,2922
=|2922,2923
=|2923,2924
=|2924,2925
=|2925,2926
=|2926,2927
=|2927,2928
=|2928,2929
=|2929,2930
=|2930,2931
=|2931,2932
=|2932,2933
=|2933,2934
=|2934,2935
=|2935,2936
=|2936,2937
=|2937,2938
=|2938,2939
=|2939,2940
=|2940,2941
=|2941,2942
=|2942,2943
=|2943,2944
=|2944,2945
<EOL>|2945,2946
VITALS|2947,2953
:|2953,2954
98.4|2955,2959
140|2960,2963
/|2963,2964
83|2964,2966
77|2967,2969
22|2970,2972
94|2973,2975
%|2975,2976
RA|2977,2979
<EOL>|2981,2982
GENERAL|2983,2990
:|2990,2991
breathing|2992,3001
somewhat|3002,3010
heavily|3011,3018
with|3019,3023
audible|3024,3031
wheeze|3032,3038
<EOL>|3040,3041
HEENT|3042,3047
-|3048,3049
no|3050,3052
pallor|3053,3059
or|3060,3062
icterus|3063,3070
,|3070,3071
no|3072,3074
oropharyngeal|3075,3088
lesion|3089,3095
,|3095,3096
no|3097,3099
sinus|3100,3105
<EOL>|3106,3107
tenderness|3107,3117
<EOL>|3119,3120
NECK|3121,3125
:|3125,3126
Supple|3127,3133
,|3133,3134
JVP|3135,3138
flat|3139,3143
<EOL>|3145,3146
CARDIAC|3147,3154
:|3154,3155
RRR|3156,3159
,|3159,3160
unable|3161,3167
to|3168,3170
appreciate|3171,3181
any|3182,3185
m|3186,3187
/|3187,3188
r|3188,3189
/|3189,3190
g|3190,3191
due|3192,3195
to|3196,3198
breathing|3199,3208
<EOL>|3210,3211
PULMONARY|3212,3221
:|3221,3222
diffuse|3223,3230
wheezes|3231,3238
and|3239,3242
ronchi|3243,3249
<EOL>|3251,3252
ABDOMEN|3253,3260
:|3260,3261
NT|3262,3264
/|3264,3265
ND|3265,3267
,|3267,3268
+|3269,3270
BS|3270,3272
<EOL>|3274,3275
EXTREMITIES|3276,3287
:|3287,3288
1|3289,3290
+|3290,3291
lower|3292,3297
extremity|3298,3307
edema|3308,3313
up|3314,3316
shins|3317,3322
,|3322,3323
patient|3324,3331
is|3332,3334
<EOL>|3335,3336
sitting|3336,3343
_|3344,3345
_|3345,3346
_|3346,3347
style|3348,3353
and|3354,3357
I|3358,3359
do|3360,3362
not|3363,3366
appreciate|3367,3377
tenderness|3378,3388
at|3389,3391
the|3392,3395
R|3396,3397
<EOL>|3398,3399
hip|3399,3402
<EOL>|3404,3405
SKIN|3406,3410
:|3410,3411
Without|3412,3419
rash|3420,3424
.|3424,3425
<EOL>|3427,3428
NEUROLOGIC|3429,3439
:|3439,3440
A|3441,3442
&|3442,3443
Ox3|3443,3446
,|3446,3447
moving|3448,3454
all|3455,3458
extremities|3459,3470
with|3471,3475
purpose|3476,3483
<EOL>|3485,3486
<EOL>|3487,3488
PHYSICAL|3488,3496
EXAMINATION|3497,3508
ON|3509,3511
DISCHARGE|3512,3521
:|3521,3522
<EOL>|3522,3523
=|3523,3524
=|3524,3525
=|3525,3526
=|3526,3527
=|3527,3528
=|3528,3529
=|3529,3530
=|3530,3531
=|3531,3532
=|3532,3533
=|3533,3534
=|3534,3535
=|3535,3536
=|3536,3537
=|3537,3538
=|3538,3539
=|3539,3540
=|3540,3541
=|3541,3542
=|3542,3543
=|3543,3544
=|3544,3545
=|3545,3546
=|3546,3547
=|3547,3548
=|3548,3549
=|3549,3550
=|3550,3551
=|3551,3552
=|3552,3553
=|3553,3554
=|3554,3555
=|3555,3556
=|3556,3557
<EOL>|3557,3558
HR|3559,3561
and|3562,3565
RR|3566,3568
went|3569,3573
to|3574,3576
zero|3577,3581
on|3582,3584
continuous|3585,3595
telemetry|3596,3605
.|3605,3606
Patient|3607,3614
did|3615,3618
not|3619,3622
<EOL>|3623,3624
respond|3624,3631
to|3632,3634
vocal|3635,3640
or|3641,3643
tactile|3644,3651
stimuli|3652,3659
.|3659,3660
Pupils|3661,3667
were|3668,3672
non-reactive|3673,3685
to|3686,3688
<EOL>|3689,3690
light|3690,3695
.|3695,3696
She|3697,3700
had|3701,3704
no|3705,3707
heart|3708,3713
or|3714,3716
lung|3717,3721
sounds|3722,3728
for|3729,3732
>|3733,3734
1|3735,3736
minute|3737,3743
on|3744,3746
<EOL>|3747,3748
auscultation|3748,3760
.|3760,3761
She|3762,3765
was|3766,3769
pronounced|3770,3780
dead|3781,3785
at|3786,3788
0515|3789,3793
.|3793,3794
Family|3795,3801
was|3802,3805
<EOL>|3806,3807
notified|3807,3815
,|3815,3816
they|3817,3821
had|3822,3825
previously|3826,3836
declined|3837,3845
an|3846,3848
autopsy|3849,3856
.|3856,3857
<EOL>|3858,3859
<EOL>|3860,3861
Pertinent|3861,3870
Results|3871,3878
:|3878,3879
<EOL>|3879,3880
LABS|3880,3884
ON|3885,3887
ADMISSION|3888,3897
:|3897,3898
<EOL>|3898,3899
=|3899,3900
=|3900,3901
=|3901,3902
=|3902,3903
=|3903,3904
=|3904,3905
=|3905,3906
=|3906,3907
=|3907,3908
=|3908,3909
=|3909,3910
=|3910,3911
=|3911,3912
=|3912,3913
=|3913,3914
=|3914,3915
=|3915,3916
=|3916,3917
<EOL>|3917,3918
_|3918,3919
_|3919,3920
_|3920,3921
04|3922,3924
:|3924,3925
38PM|3925,3929
BLOOD|3930,3935
WBC|3936,3939
-|3939,3940
7.5|3940,3943
RBC|3944,3947
-|3947,3948
4|3948,3949
.|3949,3950
39|3950,3952
Hgb|3953,3956
-|3956,3957
12.3|3957,3961
Hct|3962,3965
-|3965,3966
38.6|3966,3970
MCV|3971,3974
-|3974,3975
88|3975,3977
<EOL>|3978,3979
MCH|3979,3982
-|3982,3983
28.0|3983,3987
MCHC|3988,3992
-|3992,3993
31|3993,3995
.|3995,3996
9|3996,3997
*|3997,3998
RDW|3999,4002
-|4002,4003
18|4003,4005
.|4005,4006
0|4006,4007
*|4007,4008
RDWSD|4009,4014
-|4014,4015
56|4015,4017
.|4017,4018
9|4018,4019
*|4019,4020
Plt|4021,4024
_|4025,4026
_|4026,4027
_|4027,4028
<EOL>|4028,4029
_|4029,4030
_|4030,4031
_|4031,4032
04|4033,4035
:|4035,4036
38PM|4036,4040
BLOOD|4041,4046
Neuts|4047,4052
-|4052,4053
92|4053,4055
.|4055,4056
1|4056,4057
*|4057,4058
Lymphs|4059,4065
-|4065,4066
3|4066,4067
.|4067,4068
9|4068,4069
*|4069,4070
Monos|4071,4076
-|4076,4077
3|4077,4078
.|4078,4079
5|4079,4080
*|4080,4081
<EOL>|4082,4083
Eos|4083,4086
-|4086,4087
0|4087,4088
.|4088,4089
0|4089,4090
*|4090,4091
Baso|4092,4096
-|4096,4097
0.0|4097,4100
Im|4101,4103
_|4104,4105
_|4105,4106
_|4106,4107
AbsNeut|4108,4115
-|4115,4116
6|4116,4117
.|4117,4118
91|4118,4120
*|4120,4121
AbsLymp|4122,4129
-|4129,4130
0|4130,4131
.|4131,4132
29|4132,4134
*|4134,4135
<EOL>|4136,4137
AbsMono|4137,4144
-|4144,4145
0|4145,4146
.|4146,4147
26|4147,4149
AbsEos|4150,4156
-|4156,4157
0|4157,4158
.|4158,4159
00|4159,4161
*|4161,4162
AbsBaso|4163,4170
-|4170,4171
0|4171,4172
.|4172,4173
00|4173,4175
*|4175,4176
<EOL>|4176,4177
_|4177,4178
_|4178,4179
_|4179,4180
04|4181,4183
:|4183,4184
38PM|4184,4188
BLOOD|4189,4194
Plt|4195,4198
_|4199,4200
_|4200,4201
_|4201,4202
<EOL>|4202,4203
_|4203,4204
_|4204,4205
_|4205,4206
04|4207,4209
:|4209,4210
38PM|4210,4214
BLOOD|4215,4220
Glucose|4221,4228
-|4228,4229
143|4229,4232
*|4232,4233
UreaN|4234,4239
-|4239,4240
20|4240,4242
Creat|4243,4248
-|4248,4249
1.1|4249,4252
Na|4253,4255
-|4255,4256
135|4256,4259
<EOL>|4260,4261
K|4261,4262
-|4262,4263
3.5|4263,4266
Cl|4267,4269
-|4269,4270
91|4270,4272
*|4272,4273
HCO3|4274,4278
-|4278,4279
29|4279,4281
AnGap|4282,4287
-|4287,4288
19|4288,4290
<EOL>|4290,4291
_|4291,4292
_|4292,4293
_|4293,4294
04|4295,4297
:|4297,4298
38PM|4298,4302
BLOOD|4303,4308
ALT|4309,4312
-|4312,4313
50|4313,4315
*|4315,4316
AST|4317,4320
-|4320,4321
41|4321,4323
*|4323,4324
AlkPhos|4325,4332
-|4332,4333
73|4333,4335
TotBili|4336,4343
-|4343,4344
0.3|4344,4347
<EOL>|4347,4348
_|4348,4349
_|4349,4350
_|4350,4351
04|4352,4354
:|4354,4355
38PM|4355,4359
BLOOD|4360,4365
proBNP|4366,4372
-|4372,4373
425|4373,4376
<EOL>|4376,4377
_|4377,4378
_|4378,4379
_|4379,4380
04|4381,4383
:|4383,4384
38PM|4384,4388
BLOOD|4389,4394
Albumin|4395,4402
-|4402,4403
4.4|4403,4406
Calcium|4407,4414
-|4414,4415
10.3|4415,4419
Phos|4420,4424
-|4424,4425
3.6|4425,4428
Mg|4429,4431
-|4431,4432
2.0|4432,4435
<EOL>|4435,4436
_|4436,4437
_|4437,4438
_|4438,4439
10|4440,4442
:|4442,4443
40AM|4443,4447
BLOOD|4448,4453
_|4454,4455
_|4455,4456
_|4456,4457
pO2|4458,4461
-|4461,4462
130|4462,4465
*|4465,4466
pCO2|4467,4471
-|4471,4472
41|4472,4474
pH|4475,4477
-|4477,4478
7.42|4478,4482
<EOL>|4483,4484
calTCO2|4484,4491
-|4491,4492
28|4492,4494
Base|4495,4499
XS|4500,4502
-|4502,4503
2|4503,4504
Comment|4505,4512
-|4512,4513
GREEN|4513,4518
TOP|4519,4522
<EOL>|4522,4523
_|4523,4524
_|4524,4525
_|4525,4526
04|4527,4529
:|4529,4530
44PM|4530,4534
BLOOD|4535,4540
Lactate|4541,4548
-|4548,4549
3|4549,4550
.|4550,4551
0|4551,4552
*|4552,4553
<EOL>|4553,4554
<EOL>|4554,4555
LABS|4555,4559
ON|4560,4562
DISCHARGE|4563,4572
:|4572,4573
<EOL>|4573,4574
=|4574,4575
=|4575,4576
=|4576,4577
=|4577,4578
=|4578,4579
=|4579,4580
=|4580,4581
=|4581,4582
=|4582,4583
=|4583,4584
=|4584,4585
=|4585,4586
=|4586,4587
=|4587,4588
=|4588,4589
=|4589,4590
=|4590,4591
=|4591,4592
<EOL>|4592,4593
_|4593,4594
_|4594,4595
_|4595,4596
04|4597,4599
:|4599,4600
15AM|4600,4604
BLOOD|4605,4610
WBC|4611,4614
-|4614,4615
13|4615,4617
.|4617,4618
4|4618,4619
*|4619,4620
RBC|4621,4624
-|4624,4625
2|4625,4626
.|4626,4627
42|4627,4629
*|4629,4630
Hgb|4631,4634
-|4634,4635
7|4635,4636
.|4636,4637
0|4637,4638
*|4638,4639
Hct|4640,4643
-|4643,4644
22|4644,4646
.|4646,4647
9|4647,4648
*|4648,4649
<EOL>|4650,4651
MCV|4651,4654
-|4654,4655
95|4655,4657
MCH|4658,4661
-|4661,4662
28.9|4662,4666
MCHC|4667,4671
-|4671,4672
30|4672,4674
.|4674,4675
6|4675,4676
*|4676,4677
RDW|4678,4681
-|4681,4682
17|4682,4684
.|4684,4685
5|4685,4686
*|4686,4687
RDWSD|4688,4693
-|4693,4694
56|4694,4696
.|4696,4697
8|4697,4698
*|4698,4699
Plt|4700,4703
_|4704,4705
_|4705,4706
_|4706,4707
<EOL>|4707,4708
_|4708,4709
_|4709,4710
_|4710,4711
04|4712,4714
:|4714,4715
15AM|4715,4719
BLOOD|4720,4725
Glucose|4726,4733
-|4733,4734
94|4734,4736
UreaN|4737,4742
-|4742,4743
15|4743,4745
Creat|4746,4751
-|4751,4752
0.6|4752,4755
Na|4756,4758
-|4758,4759
138|4759,4762
<EOL>|4763,4764
K|4764,4765
-|4765,4766
4.2|4766,4769
Cl|4770,4772
-|4772,4773
97|4773,4775
HCO3|4776,4780
-|4780,4781
37|4781,4783
*|4783,4784
AnGap|4785,4790
-|4790,4791
8|4791,4792
<EOL>|4792,4793
_|4793,4794
_|4794,4795
_|4795,4796
04|4797,4799
:|4799,4800
15AM|4800,4804
BLOOD|4805,4810
Calcium|4811,4818
-|4818,4819
8|4819,4820
.|4820,4821
3|4821,4822
*|4822,4823
Phos|4824,4828
-|4828,4829
3.0|4829,4832
Mg|4833,4835
-|4835,4836
2.0|4836,4839
<EOL>|4839,4840
<EOL>|4840,4841
SELECT|4841,4847
IMAGING|4848,4855
:|4855,4856
<EOL>|4856,4857
=|4857,4858
=|4858,4859
=|4859,4860
=|4860,4861
=|4861,4862
=|4862,4863
=|4863,4864
=|4864,4865
=|4865,4866
=|4866,4867
=|4867,4868
=|4868,4869
=|4869,4870
=|4870,4871
=|4871,4872
<EOL>|4872,4873
_|4873,4874
_|4874,4875
_|4875,4876
CXR|4877,4880
:|4880,4881
<EOL>|4883,4884
COMPARISON|4884,4894
:|4894,4895
_|4896,4897
_|4897,4898
_|4898,4899
<EOL>|4901,4902
FINDINGS|4902,4910
:|4910,4911
<EOL>|4913,4914
Heart|4915,4920
size|4921,4925
is|4926,4928
mildly|4929,4935
enlarged|4936,4944
.|4944,4945
There|4946,4951
is|4952,4954
mild|4955,4959
unfolding|4960,4969
of|4970,4972
the|4973,4976
<EOL>|4977,4978
thoracic|4978,4986
aorta|4987,4992
.|4992,4993
Cardiomediastinal|4994,5011
silhouette|5012,5022
and|5023,5026
hilar|5027,5032
contours|5033,5041
<EOL>|5042,5043
are|5043,5046
otherwise|5047,5056
unremarkable|5057,5069
.|5069,5070
There|5071,5076
is|5077,5079
mild|5080,5084
bibasilar|5085,5094
atelectasis|5095,5106
.|5106,5107
<EOL>|5108,5109
Lungs|5109,5114
are|5115,5118
otherwise|5119,5128
clear|5129,5134
.|5134,5135
Pleural|5136,5143
surfaces|5144,5152
are|5153,5156
clear|5157,5162
without|5163,5170
<EOL>|5171,5172
effusion|5172,5180
or|5181,5183
pneumothorax|5184,5196
.|5196,5197
Focus|5198,5203
of|5204,5206
air|5207,5210
seen|5211,5215
under|5216,5221
the|5222,5225
right|5226,5231
<EOL>|5232,5233
hemidiaphragm|5233,5246
,|5246,5247
likely|5248,5254
represents|5255,5265
colonic|5266,5273
interposition|5274,5287
.|5287,5288
<EOL>|5290,5291
IMPRESSION|5291,5301
:|5301,5302
No|5302,5304
acute|5305,5310
cardiopulmonary|5311,5326
abnormality|5327,5338
.|5338,5339
<EOL>|5341,5342
<EOL>|5342,5343
_|5343,5344
_|5344,5345
_|5345,5346
RUE|5347,5350
U|5351,5352
/|5352,5353
S|5353,5354
:|5354,5355
<EOL>|5355,5356
IMPRESSION|5357,5367
:|5367,5368
4|5369,5370
cm|5371,5373
acute|5374,5379
deep|5380,5384
vein|5385,5389
thrombosis|5390,5400
noted|5401,5406
within|5407,5413
the|5414,5417
<EOL>|5418,5419
mid|5419,5422
right|5423,5428
brachial|5429,5437
vein|5438,5442
as|5443,5445
detailed|5446,5454
above|5455,5460
.|5460,5461
<EOL>|5462,5463
<EOL>|5463,5464
_|5464,5465
_|5465,5466
_|5466,5467
CXR|5468,5471
:|5471,5472
<EOL>|5472,5473
IMPRESSION|5474,5484
:|5484,5485
The|5486,5489
endotracheal|5490,5502
tube|5503,5507
tip|5508,5511
is|5512,5514
6|5515,5516
cm|5517,5519
above|5520,5525
the|5526,5529
carina|5530,5536
.|5536,5537
<EOL>|5538,5539
Nasogastric|5540,5551
tube|5552,5556
tip|5557,5560
is|5561,5563
beyond|5564,5570
the|5571,5574
GE|5575,5577
junction|5578,5586
and|5587,5590
off|5591,5594
the|5595,5598
edge|5599,5603
<EOL>|5604,5605
of|5605,5607
the|5608,5611
film|5612,5616
.|5616,5617
A|5619,5620
left|5621,5625
central|5626,5633
line|5634,5638
is|5639,5641
present|5642,5649
in|5650,5652
the|5653,5656
tip|5657,5660
is|5661,5663
in|5664,5666
<EOL>|5667,5668
the|5668,5671
mid|5672,5675
SVC|5676,5679
.|5679,5680
A|5682,5683
pacemaker|5684,5693
is|5694,5696
noted|5697,5702
on|5703,5705
the|5706,5709
right|5710,5715
in|5716,5718
the|5719,5722
lead|5723,5727
<EOL>|5728,5729
projects|5729,5737
over|5738,5742
the|5743,5746
right|5747,5752
ventricle|5753,5762
.|5762,5763
There|5765,5770
is|5771,5773
probable|5774,5782
scarring|5783,5791
<EOL>|5792,5793
in|5793,5795
both|5796,5800
lung|5801,5805
apices|5806,5812
.|5812,5813
There|5815,5820
are|5821,5824
no|5825,5827
new|5828,5831
areas|5832,5837
of|5838,5840
consolidation|5841,5854
.|5854,5855
<EOL>|5857,5858
There|5858,5863
is|5864,5866
upper|5867,5872
zone|5873,5877
redistribution|5878,5892
and|5893,5896
cardiomegaly|5897,5909
suggesting|5910,5920
<EOL>|5921,5922
pulmonary|5922,5931
venous|5932,5938
hypertension|5939,5951
.|5951,5952
There|5953,5958
is|5959,5961
no|5962,5964
pneumothorax|5965,5977
.|5977,5978
<EOL>|5979,5980
<EOL>|5981,5982
Brief|5982,5987
Hospital|5988,5996
Course|5997,6003
:|6003,6004
<EOL>|6004,6005
_|6005,6006
_|6006,6007
_|6007,6008
hx|6009,6011
severe|6012,6018
COPD|6019,6023
,|6023,6024
AFib|6025,6029
,|6029,6030
CAD|6031,6034
,|6034,6035
HTN|6036,6039
,|6039,6040
HLD|6041,6044
,|6044,6045
recent|6046,6052
hospitalizations|6053,6069
<EOL>|6070,6071
for|6071,6074
recurrent|6075,6084
COPD|6085,6089
exacerbations|6090,6103
over|6104,6108
the|6109,6112
last|6113,6117
several|6118,6125
months|6126,6132
,|6132,6133
<EOL>|6134,6135
who|6135,6138
presented|6139,6148
with|6149,6153
dyspnea|6154,6161
and|6162,6165
increased|6166,6175
wheezing|6176,6184
secondary|6185,6194
to|6195,6197
<EOL>|6198,6199
severe|6199,6205
COPD|6206,6210
.|6210,6211
<EOL>|6212,6213
<EOL>|6213,6214
She|6214,6217
was|6218,6221
treated|6222,6229
for|6230,6233
her|6234,6237
COPD|6238,6242
with|6243,6247
nebulizers|6248,6258
and|6259,6262
steroids|6263,6271
,|6271,6272
but|6273,6276
<EOL>|6277,6278
continued|6278,6287
to|6288,6290
decline|6291,6298
eventually|6299,6309
suffering|6310,6319
a|6320,6321
PEA|6322,6325
arrest|6326,6332
thought|6333,6340
<EOL>|6341,6342
due|6342,6345
to|6346,6348
hypoxemia|6349,6358
requiring|6359,6368
endotracheal|6369,6381
intubation|6382,6392
and|6393,6396
<EOL>|6397,6398
mechanical|6398,6408
ventilation|6409,6420
.|6420,6421
A|6422,6423
temporary|6424,6433
pacemaker|6434,6443
was|6444,6447
placed|6448,6454
for|6455,6458
<EOL>|6459,6460
periods|6460,6467
of|6468,6470
bradycardia|6471,6482
that|6483,6487
may|6488,6491
also|6492,6496
have|6497,6501
contributed|6502,6513
to|6514,6516
her|6517,6520
PEA|6521,6524
<EOL>|6525,6526
arrest|6526,6532
(|6533,6534
versus|6534,6540
being|6541,6546
a|6547,6548
manifestation|6549,6562
of|6563,6565
severe|6566,6572
hypoxemia|6573,6582
/|6582,6583
severe|6583,6589
<EOL>|6590,6591
hypercarbia|6591,6602
preceding|6603,6612
her|6613,6616
arrest|6617,6623
)|6623,6624
.|6624,6625
She|6626,6629
made|6630,6634
a|6635,6636
cognitive|6637,6646
recovery|6647,6655
<EOL>|6656,6657
but|6657,6660
was|6661,6664
unable|6665,6671
to|6672,6674
be|6675,6677
successfully|6678,6690
weaned|6691,6697
from|6698,6702
her|6703,6706
ventilator|6707,6717
.|6717,6718
<EOL>|6719,6720
She|6720,6723
had|6724,6727
capacity|6728,6736
and|6737,6740
was|6741,6744
able|6745,6749
to|6750,6752
make|6753,6757
it|6758,6760
understand|6761,6771
that|6772,6776
she|6777,6780
did|6781,6784
<EOL>|6785,6786
not|6786,6789
wish|6790,6794
:|6794,6795
continued|6796,6805
intubation|6806,6816
&|6817,6818
mechanical|6819,6829
ventilation|6830,6841
;|6841,6842
<EOL>|6843,6844
re-intubation|6844,6857
and|6858,6861
mechanical|6862,6872
ventilation|6873,6884
once|6885,6889
extubated|6890,6899
;|6899,6900
or|6901,6903
,|6903,6904
<EOL>|6905,6906
positive|6906,6914
non-invasive|6915,6927
pressure|6928,6936
ventilation|6937,6948
.|6948,6949
After|6950,6955
extensive|6956,6965
<EOL>|6966,6967
discussions|6967,6978
with|6979,6983
her|6984,6987
and|6988,6991
her|6992,6995
family|6996,7002
,|7002,7003
she|7004,7007
was|7008,7011
transitioned|7012,7024
to|7025,7027
<EOL>|7028,7029
DNR|7029,7032
/|7032,7033
DNI|7033,7036
and|7037,7040
comfort|7041,7048
-|7048,7049
oriented|7049,7057
care|7058,7062
.|7062,7063
She|7064,7067
was|7068,7071
extubated|7072,7081
to|7082,7084
spend|7085,7090
<EOL>|7091,7092
quality|7092,7099
time|7100,7104
with|7105,7109
her|7110,7113
family|7114,7120
before|7121,7127
passing|7128,7135
from|7136,7140
respiratory|7141,7152
<EOL>|7153,7154
failure|7154,7161
on|7162,7164
the|7165,7168
morning|7169,7176
of|7177,7179
_|7180,7181
_|7181,7182
_|7182,7183
at|7184,7186
0515|7187,7191
.|7191,7192
Autopsy|7193,7200
was|7201,7204
declined|7205,7213
<EOL>|7214,7215
by|7215,7217
family|7218,7224
.|7224,7225
<EOL>|7225,7226
<EOL>|7226,7227
She|7227,7230
was|7231,7234
incidentally|7235,7247
found|7248,7253
to|7254,7256
have|7257,7261
a|7262,7263
RUE|7264,7267
DVT|7268,7271
that|7272,7276
was|7277,7280
treated|7281,7288
<EOL>|7289,7290
with|7290,7294
heparin|7295,7302
gtt|7303,7306
(|7307,7308
which|7308,7313
was|7314,7317
also|7318,7322
used|7323,7327
for|7328,7331
anticoagulation|7332,7347
for|7348,7351
<EOL>|7352,7353
her|7353,7356
atrial|7357,7363
fibrillation|7364,7376
;|7376,7377
she|7378,7381
was|7382,7385
temporarily|7386,7397
transitioned|7398,7410
to|7411,7413
<EOL>|7414,7415
argatroban|7415,7425
for|7426,7429
concern|7430,7437
of|7438,7440
HIT|7441,7444
,|7444,7445
but|7446,7449
PF4|7450,7453
antibodies|7454,7464
returned|7465,7473
at|7474,7476
<EOL>|7477,7478
very|7478,7482
low|7483,7486
OD|7487,7489
,|7489,7490
making|7491,7497
this|7498,7502
diagnosis|7503,7512
unlikely|7513,7521
)|7521,7522
.|7522,7523
She|7524,7527
was|7528,7531
also|7532,7536
<EOL>|7537,7538
treated|7538,7545
for|7546,7549
an|7550,7552
acute|7553,7558
sinusitis|7559,7568
with|7569,7573
Augmentin|7574,7583
during|7584,7590
her|7591,7594
<EOL>|7595,7596
hospital|7596,7604
stay|7605,7609
.|7609,7610
<EOL>|7611,7612
<EOL>|7613,7614
Medications|7614,7625
on|7626,7628
Admission|7629,7638
:|7638,7639
<EOL>|7639,7640
The|7640,7643
Preadmission|7644,7656
Medication|7657,7667
list|7668,7672
is|7673,7675
accurate|7676,7684
and|7685,7688
complete|7689,7697
.|7697,7698
<EOL>|7698,7699
1.|7699,7701
Acetaminophen|7702,7715
325|7716,7719
mg|7720,7722
PO|7723,7725
Q4H|7726,7729
:|7729,7730
PRN|7730,7733
Pain|7734,7738
<EOL>|7739,7740
2.|7740,7742
Calcitrate|7743,7753
-|7753,7754
Vitamin|7754,7761
D|7762,7763
(|7764,7765
calcium|7765,7772
citrate|7773,7780
-|7780,7781
vitamin|7781,7788
D3|7789,7791
)|7791,7792
315|7793,7796
mg|7797,7799
-|7800,7801
<EOL>|7802,7803
200|7803,7806
units|7807,7812
oral|7814,7818
DAILY|7819,7824
<EOL>|7825,7826
3.|7826,7828
Tiotropium|7829,7839
Bromide|7840,7847
1|7848,7849
CAP|7850,7853
IH|7854,7856
DAILY|7857,7862
<EOL>|7863,7864
4.|7864,7866
Theophylline|7867,7879
SR|7880,7882
300|7883,7886
mg|7887,7889
PO|7890,7892
BID|7893,7896
<EOL>|7897,7898
5.|7898,7900
Sulfameth|7901,7910
/|7910,7911
Trimethoprim|7911,7923
SS|7924,7926
1|7927,7928
TAB|7929,7932
PO|7933,7935
DAILY|7936,7941
prophylaxis|7942,7953
for|7954,7957
long|7958,7962
<EOL>|7963,7964
term|7964,7968
steroid|7969,7976
use|7977,7980
<EOL>|7981,7982
6.|7982,7984
Ranitidine|7985,7995
300|7996,7999
mg|8000,8002
PO|8003,8005
DAILY|8006,8011
<EOL>|8012,8013
7.|8013,8015
PredniSONE|8016,8026
40|8027,8029
mg|8030,8032
PO|8033,8035
DAILY|8036,8041
<EOL>|8042,8043
8.|8043,8045
Lorazepam|8046,8055
0.5|8056,8059
mg|8060,8062
PO|8063,8065
Q8H|8066,8069
:|8069,8070
PRN|8070,8073
Insomnia|8074,8082
,|8082,8083
anxiety|8084,8091
,|8091,8092
vertigo|8093,8100
<EOL>|8101,8102
9.|8102,8104
Latanoprost|8105,8116
0.005|8117,8122
%|8122,8123
Ophth|8124,8129
.|8129,8130
Soln.|8131,8136
1|8137,8138
DROP|8139,8143
BOTH|8144,8148
EYES|8149,8153
QHS|8154,8157
<EOL>|8158,8159
10.|8159,8162
Isosorbide|8163,8173
Mononitrate|8174,8185
(|8186,8187
Extended|8187,8195
Release|8196,8203
)|8203,8204
240|8205,8208
mg|8209,8211
PO|8212,8214
DAILY|8215,8220
<EOL>|8221,8222
11.|8222,8225
Ipratropium|8226,8237
Bromide|8238,8245
Neb|8246,8249
1|8250,8251
NEB|8252,8255
IH|8256,8258
Q6H|8259,8262
Wheezing|8263,8271
<EOL>|8272,8273
12.|8273,8276
Hydrochlorothiazide|8277,8296
50|8297,8299
mg|8300,8302
PO|8303,8305
DAILY|8306,8311
<EOL>|8312,8313
13.|8313,8316
Guaifenesin|8317,8328
_|8329,8330
_|8330,8331
_|8331,8332
mL|8333,8335
PO|8336,8338
Q4H|8339,8342
:|8342,8343
PRN|8343,8346
cough|8347,8352
<EOL>|8353,8354
14.|8354,8357
Fluticasone|8358,8369
-|8369,8370
Salmeterol|8370,8380
Diskus|8381,8387
(|8388,8389
500|8389,8392
/|8392,8393
50|8393,8395
)|8395,8396
1|8398,8399
INH|8400,8403
IH|8404,8406
BID|8407,8410
<EOL>|8411,8412
15.|8412,8415
Fluticasone|8416,8427
Propionate|8428,8438
NASAL|8439,8444
2|8445,8446
SPRY|8447,8451
NU|8452,8454
DAILY|8455,8460
:|8460,8461
PRN|8461,8464
allergies|8465,8474
<EOL>|8475,8476
16|8476,8478
.|8478,8479
Ferrous|8480,8487
Sulfate|8488,8495
325|8496,8499
mg|8500,8502
PO|8503,8505
DAILY|8506,8511
<EOL>|8512,8513
17.|8513,8516
Dorzolamide|8517,8528
2|8529,8530
%|8530,8531
Ophth|8532,8537
.|8537,8538
Soln.|8539,8544
1|8545,8546
DROP|8547,8551
BOTH|8552,8556
EYES|8557,8561
BID|8562,8565
<EOL>|8566,8567
18.|8567,8570
albuterol|8571,8580
sulfate|8581,8588
90|8589,8591
mcg|8592,8595
/|8595,8596
actuation|8596,8605
inhalation|8606,8616
Q4H|8617,8620
<EOL>|8621,8622
19|8622,8624
.|8624,8625
Apixaban|8626,8634
5|8635,8636
mg|8637,8639
PO|8640,8642
BID|8643,8646
<EOL>|8647,8648
20|8648,8650
.|8650,8651
Aspirin|8652,8659
81|8660,8662
mg|8663,8665
PO|8666,8668
DAILY|8669,8674
<EOL>|8675,8676
21|8676,8678
.|8678,8679
Atorvastatin|8680,8692
10|8693,8695
mg|8696,8698
PO|8699,8701
QPM|8702,8705
<EOL>|8706,8707
22.|8707,8710
Diltiazem|8711,8720
Extended|8721,8729
-|8729,8730
Release|8730,8737
240|8738,8741
mg|8742,8744
PO|8745,8747
BID|8748,8751
<EOL>|8752,8753
23|8753,8755
.|8755,8756
Docusate|8757,8765
Sodium|8766,8772
100|8773,8776
mg|8777,8779
PO|8780,8782
BID|8783,8786
<EOL>|8787,8788
24|8788,8790
.|8790,8791
Sodium|8792,8798
Chloride|8799,8807
Nasal|8808,8813
_|8814,8815
_|8815,8816
_|8816,8817
SPRY|8818,8822
NU|8823,8825
QID|8826,8829
:|8829,8830
PRN|8830,8833
nasal|8834,8839
discomfort|8840,8850
<EOL>|8851,8852
25|8852,8854
.|8854,8855
Morphine|8856,8864
Sulfate|8865,8872
(|8873,8874
Oral|8874,8878
Solution|8879,8887
)|8887,8888
2|8889,8890
mg|8891,8893
/|8893,8894
mL|8894,8896
5|8897,8898
mg|8899,8901
PO|8902,8904
Q4H|8905,8908
:|8908,8909
PRN|8909,8912
<EOL>|8913,8914
shortness|8914,8923
of|8924,8926
breath|8927,8933
<EOL>|8934,8935
26|8935,8937
.|8937,8938
Budesonide|8939,8949
Nasal|8950,8955
Inhaler|8956,8963
180|8964,8967
mcg|8968,8971
Other|8972,8977
DAILY|8978,8983
<EOL>|8984,8985
<EOL>|8985,8986
<EOL>|8987,8988
Discharge|8988,8997
Medications|8998,9009
:|9009,9010
<EOL>|9010,9011
None|9011,9015
.|9015,9016
<EOL>|9016,9017
<EOL>|9018,9019
Discharge|9019,9028
Disposition|9029,9040
:|9040,9041
<EOL>|9041,9042
Expired|9042,9049
<EOL>|9049,9050
<EOL>|9051,9052
Discharge|9052,9061
Diagnosis|9062,9071
:|9071,9072
<EOL>|9072,9073
PRIMARY|9073,9080
DIAGNOSES|9081,9090
:|9090,9091
<EOL>|9091,9092
s|9092,9093
/|9093,9094
p|9094,9095
PEA|9096,9099
Arrest|9100,9106
<EOL>|9107,9108
Respiratory|9108,9119
Failure|9120,9127
<EOL>|9127,9128
COPD|9128,9132
<EOL>|9132,9133
Sinusitis|9133,9142
<EOL>|9142,9143
RUE|9143,9146
DVT|9147,9150
<EOL>|9150,9151
<EOL>|9151,9152
SECONDARY|9152,9161
DIAGNOSES|9162,9171
:|9171,9172
<EOL>|9172,9173
Atrial|9173,9179
fibrillation|9180,9192
<EOL>|9192,9193
Hypertension|9193,9205
<EOL>|9205,9206
CAD|9206,9209
<EOL>|9209,9210
<EOL>|9211,9212
Discharge|9212,9221
Condition|9222,9231
:|9231,9232
<EOL>|9232,9233
Deceased|9233,9241
.|9241,9242
<EOL>|9243,9244
<EOL>|9245,9246
Discharge|9246,9255
Instructions|9256,9268
:|9268,9269
<EOL>|9269,9270
N|9270,9271
/|9271,9272
A|9272,9273
<EOL>|9273,9274
<EOL>|9275,9276
Followup|9276,9284
Instructions|9285,9297
:|9297,9298
<EOL>|9298,9299
_|9299,9300
_|9300,9301
_|9301,9302
<EOL>|9302,9303

