CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Robotics|Subject|false|false||roboticnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Structure of ileal conduit|Disorder|false|false||ileal conduitnull|Ileal conduit procedure|Procedure|false|false||ileal conduitnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Surgical construction|Procedure|false|false||creationnull|Creation|Event|false|false||creationnull|Postoperative Period|Time|false|false||postopnull|Course|Time|false|false||coursenull|Bacteremia|Finding|false|false||bacteremianull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Drugs used in migraine prophylaxis|Drug|false|false||prophylacticnull|Prophylactic behavior|Finding|false|false||prophylacticnull|Condoms, Male|Device|false|false||prophylacticnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|day|Time|false|false||daysnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Initially|Time|false|false||initiallynull|Urology service|Entity|false|false||Urology servicenull|Urology|Title|false|false||Urologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Robotics|Subject|false|false||roboticnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|null|Procedure|false|false||exenterationnull|ileum|Anatomy|false|false||ilealnull|Conduit implant|Device|false|false||conduitnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Drugs used in migraine prophylaxis|Drug|false|false||prophylacticnull|Prophylactic behavior|Finding|false|false||prophylacticnull|Condoms, Male|Device|false|false||prophylacticnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|1 Month|Time|false|false||1 monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Ileus|Disorder|false|false||ileus
null|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileusnull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|TAPBP protein, human|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|TAPBP protein, human|Drug|false|false||TPNnull|TAPBP wt Allele|Finding|false|false||TPN
null|TAPBP gene|Finding|false|false||TPNnull|Parenteral Nutrition, Total|Procedure|false|false||TPNnull|Citrobacter|Entity|false|false||Citrobacternull|C-Terminal Telopeptide Type 1 Collagen, human|Drug|false|false||CTX
null|cyclophosphamide|Drug|false|false||CTX
null|cyclophosphamide|Drug|false|false||CTX
null|Crotoxin|Drug|false|false||CTX
null|Crotoxin|Drug|false|false||CTX
null|Crotoxin|Drug|false|false||CTX
null|C-Terminal Telopeptide Type 1 Collagen, human|Drug|false|false||CTXnull|Xanthomatosis, Cerebrotendinous|Disorder|false|false||CTXnull|CYP27A1 wt Allele|Finding|false|false||CTX
null|CYP27A1 gene|Finding|false|false||CTXnull|Intraabdominal Route of Administration|Finding|false|false||intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Burning Mouth Syndrome|Disorder|false|false||BMsnull|Cipro|Drug|false|false||cipro
null|Cipro|Drug|false|false||cipronull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|Bactrim|Drug|false|false||Bactrim
null|Bactrim|Drug|false|false||Bactrimnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Bilateral|Modifier|false|false||bilateralnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Deep vein thrombosis of lower limb|Disorder|false|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Duplication (finding)|Finding|false|false||duplicatednull|Duplicate|Modifier|false|false||duplicatednull|Middle|Modifier|false|false||midnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Femoral vein|Anatomy|false|false||femoral veinsnull|Femur|Anatomy|false|false||femoralnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||dailynull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Daily|Time|false|false||dailynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Improvement|Finding|false|false||improvementnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Assisted Living Facilities|Device|false|false||assisted living facilitynull|Assisted Living Facilities|Entity|false|false||assisted living facilitynull|Assisted Living|Procedure|false|false||assisted livingnull|Assisted (qualifier value)|Modifier|false|false||assistednull|Living|Finding|false|false||living
null|Household composition|Finding|false|false||living
null|Alive|Finding|false|false||livingnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Block Dosage Form|Drug|false|false||blocknull|Fixed Block|Finding|false|false||block
null|Obstruction|Finding|false|false||block
null|Blocking|Finding|false|false||blocknull|Geographic Block|Entity|false|false||blocknull|Block (unit of presentation)|LabModifier|false|false||block
null|Block Dosing Unit|LabModifier|false|false||block
null|Block (unit of measure)|LabModifier|false|false||blocknull|Catch - Finding of sensory dimension of pain|Finding|false|false||catchnull|Breath|Finding|false|false||breathnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Unable|Finding|false|false||unablenull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Step (specific stage)|Finding|false|false||stepsnull|STEPS to Enhance Physical Activity|Procedure|false|false||stepsnull|More|LabModifier|false|false||morenull|Difficult (qualifier value)|Finding|false|false||difficultnull|Bedroom|Device|false|false||bedroomnull|Bathroom|Device|false|false||bathroom
null|Toilet Facilities|Device|false|false||bathroomnull|Referral category - Ambulatory|Finding|false|false||ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||ambulatory
null|Ambulatory|Finding|false|false||ambulatory
null|Level of Care - Ambulatory|Finding|false|false||ambulatorynull|ambulatory encounter|Procedure|false|false||ambulatorynull|Specialty Type - Ambulatory|Title|false|false||ambulatorynull|Saturated|Phenomenon|false|false||saturationnull|Associated with|Modifier|false|false||associatednull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Pallor of skin|Finding|false|false||pallornull|Increased sweating|Finding|false|false||diaphoresisnull|Associated with|Modifier|false|false||associatednull|Swelling of lower limb|Finding|false|false||leg swellingnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Thigh structure|Anatomy|false|false||thighsnull|Feelings|Finding|false|false||feelnull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Associated with|Modifier|false|false||associatednull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Inspiration (function)|Finding|false|false||inspirationnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Skin rash|Finding|false|false||rashes
null|Exanthema|Finding|false|false||rashesnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Lightheadedness|Finding|false|false||lightheadednessnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Oxygen nasal cannula|Device|false|false||Nasal Cannula
null|Nasal Cannula|Device|false|false||Nasal Cannulanull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Specimen Type - Cannula|Finding|false|false||Cannula
null|null|Finding|false|false||Cannulanull|Body Parts - Cannula|Anatomy|false|false||Cannulanull|Cannula device|Device|false|false||Cannulanull|Calamus <grasshoppers>|Entity|false|false||Cannulanull|physical examination (physical finding)|Finding|false|false||physical examnull|Physical Examination|Procedure|false|false||physical examnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Benign neoplasm of the lip|Disorder|false|false||lip
null|Lymphoid interstitial pneumonia|Disorder|false|false||lipnull|SMG1 wt Allele|Finding|false|false||lip
null|SMG1 gene|Finding|false|false||lipnull|Lip structure|Anatomy|false|false||lipnull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Unable to speak (finding)|Finding|false|false||unable to speak
null|Unable to Speak at All|Finding|false|false||unable to speaknull|Unable|Finding|false|false||unablenull|Speak - language ability|Finding|false|false||speak
null|Speaking (function)|Finding|false|false||speak
null|Does speak|Finding|false|false||speaknull|Full|Modifier|false|false||fullnull|Sentence|Finding|false|false||sentencesnull|Dyspnea|Finding|false|false||short of breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|Urostomy bag|Device|false|false||urostomy pouchnull|Urostomy procedure|Procedure|false|false||urostomynull|Urological stoma|Anatomy|false|false||urostomynull|Abdominal skin pouch|Anatomy|false|false||pouchnull|Pouch - device|Device|false|false||pouchnull|Pouch (unit of presentation)|LabModifier|false|false||pouch
null|Pouch Dosing Unit|LabModifier|false|false||pouchnull|Structure of right lower quadrant of abdomen|Anatomy|false|false||RLQnull|Right lower quadrant|Modifier|false|false||RLQnull|Surgical Stoma|Anatomy|false|false||stomanull|Pink color|Modifier|false|false||pinknull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Laboratory test finding|Lab|false|false||labsnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Primed lymphocyte test|Procedure|false|false||pltnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Leukocytes|Anatomy|false|false||WBCnull|Bacteria|Entity|false|false||bactnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epinull|Exocrine pancreatic insufficiency|Disorder|false|false||epinull|Eysenck personality inventory|Finding|false|false||epi
null|TFPI wt Allele|Finding|false|false||epi
null|TFPI gene|Finding|false|false||epinull|Electronic Portal Imaging|Procedure|false|false||epi
null|Echo-Planar Imaging|Procedure|false|false||epinull|Neg - answer|Finding|false|false||negnull|Negative - qualifier|Modifier|false|false||negnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Extensive|Modifier|false|false||Extensivenull|Pulmonary Embolism|Finding|false|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Right pulmonary artery|Anatomy|false|false||right main pulmonary artery
null|Right pulmonary arterial tree|Anatomy|false|false||right main pulmonary arterynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Main|Modifier|false|false||main
null|Primary|Modifier|false|false||mainnull|Pulmonary artery structure|Anatomy|false|false||pulmonary arterynull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Segmental|Modifier|false|false||segmentalnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Structure of lobe of lung|Anatomy|false|false||lobe pulmonarynull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Right side of heart|Anatomy|false|false||right heartnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Muscle strain|Disorder|true|false||strainnull|Nature of Abnormal Testing - Strain|Finding|true|false||strain
null|Straining (finding)|Finding|true|false||strain
null|strain symptom|Finding|true|false||strain
null|Emotional Strain|Finding|true|false||strainnull|Organism Strain|Entity|true|false||strainnull|Microbiological strain|Modifier|false|false||strainnull|Smaller|Modifier|false|false||smallernull|Small|LabModifier|false|false||smallernull|Pulmonary Embolism|Finding|false|false||pulmonary embolinull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolus|Finding|false|false||embolinull|Segmental|Modifier|false|false||segmentalnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|lobe|Anatomy|false|false||lobesnull|Several|LabModifier|false|false||Severalnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Largest|LabModifier|false|false||largestnull|Structure of middle lobe of right lung|Anatomy|false|false||right middle lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of middle lobe of right lung|Anatomy|false|false||middle lobenull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Suspicious for Malignancy|Finding|false|false||suspicious for malignancynull|Suspicious|Modifier|false|false||suspiciousnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|PET/CT scan|Procedure|false|false||PET-CTnull|Tomography, Emission-Computed|Procedure|false|false||PET
null|Positron-Emission Tomography|Procedure|false|false||PETnull|Pet Animal|Entity|false|false||PETnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Mass in breast|Finding|false|false||breast nodulesnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Correlation|Modifier|false|false||correlationnull|Mammography, Female|Procedure|false|false||mammography
null|Mammography|Procedure|false|false||mammographynull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|Frequently|Time|false|false||frequentnull|Atrial Premature Complexes|Disorder|false|false||PACnull|Atrial Premature Complex by ECG Finding|Finding|false|false||PAC
null|PACC1 gene|Finding|false|false||PACnull|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||PAC
null|CAP Regimen|Procedure|false|false||PACnull|protein aggregate center|Anatomy|false|false||PACnull|P1 Bacteriophage Artificial Chromosomes|Device|false|false||PACnull|Political action committee|Entity|false|false||PACnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|ciprofloxacin hydrochloride|Drug|false|false||Ciprofloxacin HCl
null|ciprofloxacin hydrochloride|Drug|false|false||Ciprofloxacin HClnull|ciprofloxacin|Drug|false|false||Ciprofloxacin
null|ciprofloxacin|Drug|false|false||Ciprofloxacinnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Transfer - product ownership|Finding|false|false||Transfer
null|Transfer Technique|Finding|false|false||Transfer
null|ActClass - transfer|Finding|false|false||Transfer
null|null|Finding|false|false||Transfernull|Transfer (immobility management)|Procedure|false|false||Transfernull|Oxygen nasal cannula|Device|false|false||Nasal Cannula
null|Nasal Cannula|Device|false|false||Nasal Cannulanull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Specimen Type - Cannula|Finding|false|false||Cannula
null|null|Finding|false|false||Cannulanull|Body Parts - Cannula|Anatomy|false|false||Cannulanull|Cannula device|Device|false|false||Cannulanull|Calamus <grasshoppers>|Entity|false|false||Cannulanull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Exertion|Finding|false|false||exertionnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Palpitations|Finding|true|false||palpitationsnull|Lightheadedness|Finding|false|false||lightheadednessnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Reactive Oxygen Species|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|Reactive Oxygen Species|Drug|false|false||ROSnull|ROS1 wt Allele|Finding|false|false||ROS
null|ROS1 gene|Finding|false|false||ROSnull|Review of systems (procedure)|Procedure|false|false||ROSnull|rostral sulcus|Anatomy|false|false||ROSnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Cholecystectomy, Laparoscopic|Procedure|false|false||laparoscopic cholecystectomynull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Cholecystectomy procedure|Procedure|false|false||cholecystectomynull|Structure of left knee region|Anatomy|false|false||left knee
null|Structure of left knee|Anatomy|false|false||left kneenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Laminectomy|Procedure|false|false||laminectomynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Robot Device|Device|false|false||Robot
null|null|Device|false|false||Robotnull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Bilateral|Modifier|false|false||bilateralnull|Pelvic lymph node group|Anatomy|false|false||pelvic lymph nodenull|Pelvis|Anatomy|false|false||pelvicnull|lymph nodes|Anatomy|false|false||lymph nodenull|Lymph|Finding|false|false||lymphnull|Dissecting hemorrhage|Finding|false|false||dissectionnull|Tissue Dissection|Procedure|false|false||dissectionnull|Robot Device|Device|false|false||Robot
null|null|Device|false|false||Robotnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Bilateral oophorectomy|Procedure|false|false||bilateral oophorectomynull|Bilateral|Modifier|false|false||bilateralnull|Ovariectomy|Procedure|false|false||oophorectomynull|Enlarged uterus|Finding|false|false||large uterusnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Neoplasm of uncertain or unknown behavior of uterus|Disorder|false|false||uterus
null|Uterine Diseases|Disorder|false|false||uterusnull|examination of uterus|Procedure|false|false||uterusnull|Pelvis>Uterus|Anatomy|false|false||uterus
null|Mouse Uterus|Anatomy|false|false||uterus
null|Uterus|Anatomy|false|false||uterusnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|gram|LabModifier|false|false||gramsnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Fibroid Tumor|Disorder|false|false||fibroidnull|Laparoscopic radical cystectomy|Procedure|false|false||Laparoscopic radical cystectomynull|Laparoscopy|Procedure|false|false||Laparoscopicnull|Laparoscopic approach|Modifier|false|false||Laparoscopicnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Reconstruction of vagina|Procedure|false|false||vaginal reconstructionnull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Optical Image Reconstruction|Procedure|false|false||reconstruction
null|Reconstructive Surgical Procedures|Procedure|false|false||reconstructionnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Negative|Finding|false|false||Negative fornull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Malignant neoplasm of urinary bladder|Disorder|false|false||bladder CAnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Term (lexical)|Finding|false|false||wordnull|Sentence|Finding|false|false||sentencesnull|Benign neoplasm of the lip|Disorder|false|false||lip
null|Lymphoid interstitial pneumonia|Disorder|false|false||lipnull|SMG1 wt Allele|Finding|false|false||lip
null|SMG1 gene|Finding|false|false||lipnull|Lip structure|Anatomy|false|false||lipnull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Eye|Anatomy|false|false||Eyesnull|null|Attribute|false|false||Eyesnull|Anicteric|Finding|false|false||anictericnull|ENT problem|Finding|false|false||ENT
null|NT5E gene|Finding|false|false||ENT
null|NT5E wt Allele|Finding|false|false||ENTnull|Structure of entorhinal cortex|Anatomy|false|false||ENT
null|Ear, nose and throat|Anatomy|false|false||ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|MAS1L gene|Finding|true|false||MRGnull|Full|Modifier|false|false||fullnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Compression Stockings|Device|false|false||compression stockings
null|Support stockings - garment|Device|false|false||compression stockingsnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Stocking (hosiery)|Device|false|false||stockings
null|Socks|Device|false|false||stockingsnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Jugular venous engorgement|Finding|true|false||JVDnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Exertion|Finding|false|false||effortnull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Lung|Anatomy|false|false||lungsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Auscultation|Procedure|false|false||auscultationnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Urostomy Site|Finding|false|false||Urostomy sitenull|Urostomy procedure|Procedure|false|false||Urostomynull|Urological stoma|Anatomy|false|false||Urostomynull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Infected|Finding|false|false||infectednull|Medullary sponge kidney|Disorder|false|false||MSK
null|Medullary sponge kidney|Disorder|false|false||MSKnull|SIK1 gene|Finding|false|false||MSKnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Kyphosis deformity of spine|Disorder|true|false||kyphosis
null|Acquired kyphosis|Disorder|true|false||kyphosis
null|Congenital kyphosis|Disorder|true|false||kyphosisnull|kyphosis|Finding|true|false||kyphosisnull|Palpable|Modifier|false|false||palpablenull|Synovitis|Disorder|true|false||synovitisnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Visible|Modifier|false|false||visiblenull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|jaundice|Finding|true|false||jaundice
null|Icterus|Finding|true|false||jaundice
null|yellow skin or eyes (symptom)|Finding|true|false||jaundicenull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Facial Paresis|Disorder|true|false||facial droopnull|Unilateral facial palsy|Finding|true|false||facial droopnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|Full|Modifier|false|false||Fullnull|Concept model range (foundation metadata concept)|Finding|false|false||rangenull|Sample Range|LabModifier|false|false||range
null|Range|LabModifier|false|false||rangenull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Lying in bed|Modifier|false|false||Lying in bednull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|apparent|Finding|true|false||apparentnull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Anicteric|Finding|false|false||Anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Cardiovascular system|Anatomy|false|false||Cardiovascular
null|Cardiovascular|Anatomy|false|false||Cardiovascularnull|Right sided|Modifier|false|false||right sided
null|Right|Modifier|false|false||right sidednull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Chronic obstructive pulmonary disease of horses|Disorder|true|false||heavenull|Systolic Murmurs|Finding|false|false||systolic murmurnull|Systole|Finding|false|false||systolicnull|Heart murmur|Finding|false|false||murmurnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Lung diseases|Disorder|false|false||Lungnull|Lung Problem|Finding|false|false||Lungnull|Chest>Lung|Anatomy|false|false||Lung
null|Lung|Anatomy|false|false||Lungnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Auscultation|Procedure|false|false||auscultationnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Wheezing|Finding|false|false||wheezingnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Urostomy procedure|Procedure|false|false||urostomynull|Urological stoma|Anatomy|false|false||urostomynull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Structure of left lower leg|Anatomy|false|false||left leg
null|Left lower extremity|Anatomy|false|false||left legnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower extremity>Lower leg|Anatomy|false|false||lower leg
null|Leg|Anatomy|false|false||lower legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Laboratory test finding|Lab|false|false||LABSnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||labsnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Laboratory test finding|Lab|false|false||labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood iron measurement|Procedure|false|false||BLOOD Ironnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Bacterial|Modifier|false|false||BACTERIALnull|Colony (cells or organisms)|Anatomy|false|false||COLONYnull|colonies (qualifier value)|LabModifier|false|false||COLONYnull|null|Modifier|false|false||TYPESnull|Consistent with|Finding|false|false||CONSISTENTnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Specimen Type - Genital|Finding|false|false||GENITAL
null|null|Finding|false|false||GENITALnull|Genital system|Anatomy|false|false||GENITAL
null|Genitalia|Anatomy|false|false||GENITALnull|Contamination|Finding|false|false||CONTAMINATIONnull|adulteration|Phenomenon|false|false||CONTAMINATIONnull|Specimen Reject Reason - Contamination|Modifier|false|false||CONTAMINATIONnull|Enterococcus|Entity|false|false||ENTEROCOCCUS SPnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|cfu/mL|LabModifier|false|false||CFU/mLnull|Colony-forming unit|LabModifier|false|false||CFUnull|per milliliter|LabModifier|false|false||/mLnull|Predominate|Modifier|false|false||PREDOMINATINGnull|Organism|Entity|false|false||ORGANISMnull|Interprets|Finding|false|false||INTERPRETnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|Enterococcus|Entity|false|false||ENTEROCOCCUS SPnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|ampicillin|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillin|Drug|false|false||AMPICILLINnull|nitrofurantoin|Drug|false|false||NITROFURANTOIN
null|nitrofurantoin|Drug|false|false||NITROFURANTOINnull|Tetracycline Antibiotics|Drug|false|false||TETRACYCLINE
null|Tetracycline Antibiotics|Drug|false|false||TETRACYCLINE
null|tetracycline|Drug|false|false||TETRACYCLINE
null|tetracycline|Drug|false|false||TETRACYCLINEnull|Tetracyclines causing adverse effects in therapeutic use|Disorder|false|false||TETRACYCLINEnull|vancomycin|Drug|false|false||VANCOMYCIN
null|vancomycin|Drug|false|false||VANCOMYCINnull|Vancomycin measurement|Procedure|false|false||VANCOMYCINnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Hilar|Modifier|false|false||Hilarnull|Congestion|Finding|false|false||congestionnull|Immune thrombocytopenic purpura|Disorder|false|false||franknull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Pneumonia|Disorder|false|false||pneumonianull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Extensive|Modifier|false|false||Extensivenull|Pulmonary Embolism|Finding|false|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Right pulmonary artery|Anatomy|false|false||right main pulmonary artery
null|Right pulmonary arterial tree|Anatomy|false|false||right main pulmonary arterynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Main|Modifier|false|false||main
null|Primary|Modifier|false|false||mainnull|Pulmonary artery structure|Anatomy|false|false||pulmonary arterynull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Segmental|Modifier|false|false||segmentalnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Structure of lobe of lung|Anatomy|false|false||lobe pulmonarynull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Right side of heart|Anatomy|false|false||right heartnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Muscle strain|Disorder|true|false||strainnull|Nature of Abnormal Testing - Strain|Finding|true|false||strain
null|Straining (finding)|Finding|true|false||strain
null|strain symptom|Finding|true|false||strain
null|Emotional Strain|Finding|true|false||strainnull|Organism Strain|Entity|true|false||strainnull|Microbiological strain|Modifier|false|false||strainnull|Smaller|Modifier|false|false||smallernull|Small|LabModifier|false|false||smallernull|Pulmonary Embolism|Finding|false|false||pulmonary embolinull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolus|Finding|false|false||embolinull|Segmental|Modifier|false|false||segmentalnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|lobe|Anatomy|false|false||lobesnull|Several|LabModifier|false|false||Severalnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Largest|LabModifier|false|false||largestnull|Structure of middle lobe of right lung|Anatomy|false|false||right middle lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of middle lobe of right lung|Anatomy|false|false||middle lobenull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Suspicious for Malignancy|Finding|false|false||suspicious for malignancynull|Suspicious|Modifier|false|false||suspiciousnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|PET/CT scan|Procedure|false|false||PET-CTnull|Tomography, Emission-Computed|Procedure|false|false||PET
null|Positron-Emission Tomography|Procedure|false|false||PETnull|Pet Animal|Entity|false|false||PETnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Mass in breast|Finding|false|false||breast nodulesnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Correlation|Modifier|false|false||correlationnull|Mammography, Female|Procedure|false|false||mammography
null|Mammography|Procedure|false|false||mammographynull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Deep vein thrombosis of lower limb|Disorder|false|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Occlusive thrombus|Disorder|false|false||occlusive thrombusnull|Occluded|Finding|false|false||occlusivenull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Femoral vein|Anatomy|false|false||femoral veinnull|Femur|Anatomy|false|false||femoralnull|Veins|Anatomy|false|false||veinnull|Middle|Modifier|false|false||midnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Femoral vein|Anatomy|false|false||femoral veinnull|Femur|Anatomy|false|false||femoralnull|Veins|Anatomy|false|false||veinnull|Additional|Finding|false|false||additionalnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Structure of profunda femoris vein|Anatomy|false|false||deep femoral veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Femoral vein|Anatomy|false|false||femoral veinnull|Femur|Anatomy|false|false||femoralnull|Veins|Anatomy|false|false||veinnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Femur|Anatomy|false|false||femoralnull|Structure of popliteal vein|Anatomy|false|false||popliteal veinsnull|popliteal|Anatomy|false|false||poplitealnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Bilateral|Modifier|false|false||bilateralnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Procedure on vein|Procedure|true|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|false|false||thrombosisnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Conclusion|Finding|false|false||Conclusionsnull|Left atrial structure|Anatomy|false|false||left atriumnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false||atriumnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Heart Atrium|Anatomy|false|false||atrialnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mmHgnull|Wall of left ventricle|Anatomy|false|false||Left ventricular wallnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|cardiac evaluation of ventricular wall thickness|Finding|false|false||ventricular wall thicknessnull|Wall of ventricle|Anatomy|false|false||ventricular wallnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Thick|Modifier|false|false||thicknessnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Doppler studies|Procedure|false|false||Dopplernull|Observation parameter|Finding|false|false||parametersnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Grade|Finding|false|false||with Gradenull|Grade 1 (qualifier value)|Finding|false|false||Grade I
null|Tumor grade G1|Finding|false|false||Grade I
null|Clavien-Dindo Grade I|Finding|false|false||Grade Inull|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Diastolic dysfunction|Finding|false|false||diastolic dysfunctionnull|Diastole|Attribute|false|false||diastolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|AORTIC VALVE DISEASE 3|Disorder|true|false||aortic valve stenosis
null|Stenosis of aorta|Disorder|true|false||aortic valve stenosisnull|Aortic Valve Stenosis|Finding|true|false||aortic valve stenosisnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|true|false||stenosisnull|Stenosis <Pimeliinae>|Entity|true|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Plain chest X-ray|Procedure|false|false||CXRnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Plain x-ray|Procedure|false|false||radiographsnull|heart size|Finding|false|false||Heart sizenull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pleural Diseases|Disorder|true|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Congenital Abnormality|Disorder|false|false||abnormalitynull|Abnormality|Finding|false|false||abnormalitynull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Central lymph|Finding|false|false||central lymphnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|Lymphadenopathy|Disorder|false|false||lymph node enlargementnull|Swollen Lymph Node|Finding|false|false||lymph node enlargementnull|lymph nodes|Anatomy|false|false||lymph nodenull|Lymph|Finding|false|false||lymphnull|Enlargement (morphologic abnormality)|Disorder|false|false||enlargementnull|Hypertrophy|Finding|false|false||enlargementnull|Enlargement procedure|Procedure|false|false||enlargementnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Robotics|Subject|false|false||roboticnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Bacteremia|Finding|false|false||bacteremianull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Current (present time)|Time|false|false||currentlynull|Daily|Time|false|false||dailynull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Due to|Finding|false|false||due tonull|Due to|Finding|false|false||due
null|Due|Finding|false|false||duenull|Undertreatment|Procedure|false|false||undertreatmentnull|Known|Modifier|false|false||knownnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Drugs used in migraine prophylaxis|Drug|false|false||prophylacticnull|Prophylactic behavior|Finding|false|false||prophylacticnull|Condoms, Male|Device|false|false||prophylacticnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Charge Type Reason - Treatment Failure|Finding|false|false||treatment failure
null|treatment failure|Finding|false|false||treatment failure
null|Absent response to treatment|Finding|false|false||treatment failurenull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Inspiratory Vital Capacity Test|Procedure|false|false||IVCnull|lamina IVC|Anatomy|false|false||IVCnull|filter information process|Finding|false|false||filter
null|Specimen Type - Filter|Finding|false|false||filter
null|null|Finding|false|false||filter
null|Filter (function)|Finding|false|false||filternull|Filter - medical device|Device|false|false||filter
null|Optical filter|Device|false|false||filter
null|Filters|Device|false|false||filternull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Right side of heart|Anatomy|false|false||right heartnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Muscle strain|Disorder|true|false||strainnull|Nature of Abnormal Testing - Strain|Finding|true|false||strain
null|Straining (finding)|Finding|true|false||strain
null|strain symptom|Finding|true|false||strain
null|Emotional Strain|Finding|true|false||strainnull|Organism Strain|Entity|true|false||strainnull|Microbiological strain|Modifier|false|false||strainnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Right side of heart|Anatomy|false|false||right heartnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Muscle strain|Disorder|true|false||strainnull|Nature of Abnormal Testing - Strain|Finding|true|false||strain
null|Straining (finding)|Finding|true|false||strain
null|strain symptom|Finding|true|false||strain
null|Emotional Strain|Finding|true|false||strainnull|Organism Strain|Entity|true|false||strainnull|Microbiological strain|Modifier|false|false||strainnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Thrombosis|Finding|false|false||thrombosisnull|clotrimazole|Drug|false|false||CLOT
null|clotrimazole|Drug|false|false||CLOTnull|Blood Clot|Finding|false|false||CLOTnull|Clinical Trials|Procedure|false|false||trialnull|Symptomatic|Finding|false|false||symptomaticnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Dietary Supplementation|Procedure|false|false||supplementationnull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Multiple Pulmonary Nodules|Finding|false|false||Pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Known|Modifier|false|false||Knownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Malignant neoplasm of lung|Disorder|false|false||lung malignancynull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|ETV3 wt Allele|Finding|false|false||mets
null|ETV3 gene|Finding|false|false||metsnull|Electrical Current|Phenomenon|false|false||Currentnull|Current (present time)|Time|false|false||Currentnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Still|Disorder|false|false||stillnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false||thoracicnull|Chest|Anatomy|false|false||thoracicnull|Team|Subject|false|false||teamnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Primary Care Provider - Provider role|Finding|false|false||primary care providernull|null|Attribute|false|false||primary care providernull|Primary care provider|Subject|false|false||primary care providernull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|Enterococcus|Entity|false|false||Enterococcalnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Leukocytes|Anatomy|false|false||WBCnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Urostomy procedure|Procedure|false|false||urostomynull|Urological stoma|Anatomy|false|false||urostomynull|Enterococcus|Entity|false|false||Enterococcusnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|On IV|Finding|false|false||on IVnull|ampicillin|Drug|false|false||Ampicillin
null|ampicillins|Drug|false|false||Ampicillin
null|ampicillins|Drug|false|false||Ampicillin
null|ampicillin|Drug|false|false||Ampicillinnull|Macrobid|Drug|false|false||macrobid
null|Macrobid|Drug|false|false||macrobidnull|Leukocytosis|Disorder|false|false||Leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||Leukocytosisnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Day 7|Finding|false|false||day 7null|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|true|false||bleedingnull|Hemolysis (biological function)|Finding|true|false||hemolysis
null|null|Finding|true|false||hemolysis
null|Hemolysis (finding)|Finding|true|false||hemolysis
null|Hemolysis (disorder)|Finding|true|false||hemolysisnull|Specimen Reject Reason - Hemolysis|Modifier|false|false||hemolysisnull|Lowest|Modifier|false|false||nadirnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Scientific Study|Procedure|false|false||studiesnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Iron deficiency anemia|Disorder|false|false||iron deficiency
null|Iron deficiency|Disorder|false|false||iron deficiencynull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Anemia of chronic disease|Disorder|false|false||anemia of chronic diseasenull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Chronic disease|Disorder|false|false||chronic diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Disease|Disorder|false|false||diseasenull|Iron low|Finding|false|false||low ironnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritinnull|Ferritin measurement|Procedure|false|false||ferritinnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Total iron binding capacity measurement|Procedure|false|false||TIBCnull|Total Iron-Binding Capacity result|Lab|false|false||TIBCnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Multifactorial|Finding|false|false||multifactorialnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Insufficiency|Finding|false|false||insufficiencynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Known|Modifier|false|false||knownnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Compression Stockings|Device|false|false||compression stockings
null|Support stockings - garment|Device|false|false||compression stockingsnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Stocking (hosiery)|Device|false|false||stockings
null|Socks|Device|false|false||stockingsnull|Malignant neoplasm of urinary bladder|Disorder|false|false||bladder cancer
null|Carcinoma of bladder|Disorder|false|false||bladder cancer
null|Bladder Neoplasm|Disorder|false|false||bladder cancernull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Transurethral resection of neoplasm of bladder|Procedure|false|false||TURBTnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Membrane Attack Complex|Drug|false|false||TCC
null|triclocarban|Drug|false|false||TCC
null|triclocarban|Drug|false|false||TCC
null|Membrane Attack Complex|Drug|false|false||TCCnull|TARSAL-CARPAL COALITION SYNDROME|Disorder|false|false||TCCnull|membrane attack complex location|Anatomy|false|false||TCCnull|Muscle (organ)|Anatomy|true|false||muscle
null|Muscle Tissue|Anatomy|true|false||musclenull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Magnetic Resonance Imaging (MRI) of Pelvis|Procedure|false|false||pelvic MRInull|Pelvis|Anatomy|false|false||pelvicnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Mass of urinary bladder|Finding|false|false||bladder massnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Tumor Cell Invasion|Disorder|false|false||invasionnull|Cell Invasion|Finding|false|false||invasionnull|Neck+Chest>Soft tissue|Anatomy|false|false||soft tissue
null|soft tissue|Anatomy|false|false||soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false||tissuenull|Body tissue|Anatomy|false|false||tissuenull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Walls of a building|Device|false|false||wallnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Robotics|Subject|false|false||roboticnull|Total abdominal hysterectomy|Procedure|false|false||TAHnull|Tahitian language|Entity|false|false||TAHnull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|pT2b TNM Finding|Finding|false|false||pT2bnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Infantile Neuroaxonal Dystrophy|Disorder|true|false||plannull|Treatment Plan|Finding|true|false||plan
null|Planned|Finding|true|false||plan
null|null|Finding|true|false||plannull|Further|Modifier|false|false||furthernull|Therapy Object (animal model)|Finding|true|false||therapy
null|therapeutic aspects|Finding|true|false||therapynull|Therapeutic procedure|Procedure|true|false||therapynull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Chest CT|Procedure|false|false||chest CTnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|month|Time|false|false||monthsnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Macrobid|Drug|false|false||macrobid
null|Macrobid|Drug|false|false||macrobidnull|Day 7|Finding|false|false||day 7null|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Ambulatory Status - Oxygen therapy|Finding|false|false||oxygen therapynull|Oxygen Therapy Care|Procedure|false|false||oxygen therapy
null|Warburg Therapy|Procedure|false|false||oxygen therapynull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Weaning|Finding|false|false||weannull|Maintain brand of benzocaine|Drug|false|false||maintainnull|Maintenance|Event|false|false||maintainnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Medical Product Stability|Modifier|false|false||stability
null|Stable status|Modifier|false|false||stabilitynull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|nitrofurantoin|Drug|false|false||Nitrofurantoin
null|nitrofurantoin|Drug|false|false||Nitrofurantoinnull|Macrobid|Drug|false|false||MacroBID
null|Macrobid|Drug|false|false||MacroBIDnull|Every twelve hours|Time|false|false||Q12Hnull|Last|Modifier|false|false||Lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|lorazepam|Drug|false|false||lorazepam
null|lorazepam|Drug|false|false||lorazepamnull|Tablet Dosage Form|Drug|false|false||tabnull|Tablet Dosing Unit|LabModifier|false|false||tabnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|has wheelchair at home (history)|Finding|false|false||wheelchair
null|Wheelchair Usually Used|Finding|false|false||wheelchairnull|wheelchair|Device|false|false||wheelchairnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Lung|Anatomy|false|false||lungsnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions