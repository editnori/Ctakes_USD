 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|153,165|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|153,165|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|168,177|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|168,177|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|168,177|false|false|false|C0020517|Hypersensitivity|Allergies
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|180,191|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|180,191|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|180,191|false|false|false|C0030842|penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|180,191|false|false|false|||Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|180,191|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|194,203|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|194,203|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|211,226|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|217,226|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|217,226|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|217,226|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|228,233|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|SIMPLE_SEGMENT|228,233|false|false|false|||Wound
Finding|Body Substance|SIMPLE_SEGMENT|228,233|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|228,233|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|228,233|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Pathologic Function|SIMPLE_SEGMENT|228,243|false|false|false|C0043241|Wound Infection|Wound Infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|234,243|false|false|false|C0009450|Communicable Diseases|Infection
Event|Event|SIMPLE_SEGMENT|234,243|false|false|false|||Infection
Finding|Pathologic Function|SIMPLE_SEGMENT|234,243|false|false|false|C3714514|Infection|Infection
Finding|Classification|SIMPLE_SEGMENT|246,251|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|252,260|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|252,260|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|264,282|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|273,282|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|273,282|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|273,282|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|273,282|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|273,282|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|284,289|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Event|Event|SIMPLE_SEGMENT|290,300|false|false|false|||Craniotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|290,300|false|false|false|C0010280|Craniotomy|Craniotomy
Event|Event|SIMPLE_SEGMENT|305,315|false|false|false|||Evacuation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|305,315|false|false|false|C1282573|Evacuation procedure|Evacuation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|319,326|false|false|false|C0000833|Abscess|Abscess
Event|Event|SIMPLE_SEGMENT|319,326|false|false|false|||Abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|319,326|false|false|false|C1546533||Abscess
Event|Event|SIMPLE_SEGMENT|336,343|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|336,343|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|336,343|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|336,343|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|336,346|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|336,362|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|336,362|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|347,354|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|347,354|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|347,362|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|355,362|false|false|false|C0221423|Illness (finding)|Illness
Finding|Finding|SIMPLE_SEGMENT|398,418|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|past medical history
Finding|Functional Concept|SIMPLE_SEGMENT|403,410|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|403,410|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|403,410|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|403,410|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|403,418|false|false|false|C0262926|Medical History|medical history
Event|Event|SIMPLE_SEGMENT|411,418|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|411,418|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|411,418|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|411,418|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|432,437|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|447,452|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|447,452|false|false|false|C0006111|Brain Diseases|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|447,460|false|false|false|C0006105;C1510428|Brain Abscess;Cerebral abscess|brain abscess
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|453,460|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|453,460|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|453,460|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|471,481|false|false|false|||discovered
Finding|Idea or Concept|SIMPLE_SEGMENT|500,505|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|500,505|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|SIMPLE_SEGMENT|506,509|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|520,529|false|false|false|||presented
Finding|Functional Concept|SIMPLE_SEGMENT|535,539|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|535,543|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|540,543|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|540,543|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|SIMPLE_SEGMENT|540,543|false|false|false|||arm
Finding|Gene or Genome|SIMPLE_SEGMENT|540,543|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|540,543|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|540,543|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|540,543|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Location or Region|SIMPLE_SEGMENT|549,553|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|549,553|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|549,553|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|549,553|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Finding|Sign or Symptom|SIMPLE_SEGMENT|549,562|false|false|false|C0239511|Numbness of face|face numbness
Event|Event|SIMPLE_SEGMENT|554,562|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|554,562|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|554,562|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|568,575|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|568,575|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|568,575|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|580,587|false|false|false|||drained
Event|Event|SIMPLE_SEGMENT|628,635|false|false|false|||started
Finding|Conceptual Entity|SIMPLE_SEGMENT|645,653|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|SIMPLE_SEGMENT|654,665|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|654,665|false|false|false|||antibiotics
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|673,680|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|673,680|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|673,680|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|673,680|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|673,680|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|681,685|false|false|false|||data
Finding|Idea or Concept|SIMPLE_SEGMENT|681,685|false|false|false|C1511726|Data|data
Event|Event|SIMPLE_SEGMENT|686,694|false|false|false|||returned
Finding|Intellectual Product|SIMPLE_SEGMENT|740,744|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|745,757|false|false|false|||transitioned
Drug|Antibiotic|SIMPLE_SEGMENT|761,772|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|761,772|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Event|Event|SIMPLE_SEGMENT|779,783|false|false|false|||q12h
Drug|Organic Chemical|SIMPLE_SEGMENT|789,795|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|789,795|false|false|false|C0699678|Flagyl|flagyl
Event|Event|SIMPLE_SEGMENT|802,805|false|false|false|||TID
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|847,851|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|852,856|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|852,856|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|852,856|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|852,856|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|852,856|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|874,878|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|899,905|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|906,909|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|906,909|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|906,909|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|906,909|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|930,938|false|false|false|||revealed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|949,954|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|949,954|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|949,954|false|false|false|C0013604|Edema|edema
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|971,975|false|false|false|C1882953|Ring Dosage Form|ring
Event|Event|SIMPLE_SEGMENT|976,985|false|false|false|||enhancing
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|986,997|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|986,997|false|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|986,997|false|false|false|C1704258|Abnormality|abnormality
Finding|Functional Concept|SIMPLE_SEGMENT|1005,1010|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Procedure|Health Care Activity|SIMPLE_SEGMENT|1020,1028|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1020,1028|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1029,1033|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|1029,1033|false|false|false|C1546778||site
Event|Event|SIMPLE_SEGMENT|1050,1057|false|false|false|||ongoing
Finding|Idea or Concept|SIMPLE_SEGMENT|1050,1057|false|false|false|C0549178|Continuous|ongoing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1058,1065|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|1058,1065|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|1058,1065|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|1085,1094|false|false|false|||scheduled
Finding|Functional Concept|SIMPLE_SEGMENT|1099,1105|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|1106,1114|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|1106,1114|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|1106,1114|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1106,1114|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|1131,1135|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|1142,1152|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|1142,1152|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|1142,1152|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1160,1170|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1160,1178|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1171,1178|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|1171,1178|false|false|false|||disease
Finding|Idea or Concept|SIMPLE_SEGMENT|1179,1185|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|1209,1220|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|1233,1241|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|1249,1257|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|1262,1265|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1262,1265|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1276,1286|false|false|false|||broadening
Drug|Antibiotic|SIMPLE_SEGMENT|1294,1304|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|1294,1304|false|false|false|||antibiotic
Event|Event|SIMPLE_SEGMENT|1305,1312|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|1305,1312|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1305,1312|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|1322,1330|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|1322,1330|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|1322,1330|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1322,1330|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|1337,1343|false|false|false|||states
Finding|Idea or Concept|SIMPLE_SEGMENT|1363,1368|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|1363,1368|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|SIMPLE_SEGMENT|1374,1382|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1374,1382|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|1374,1382|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1395,1399|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1400,1415|false|false|false|C1140618|Upper Extremity|upper extremity
Finding|Sign or Symptom|SIMPLE_SEGMENT|1400,1424|false|false|false|C0751409|Upper Extremity Paresis|upper extremity weakness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1406,1415|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|SIMPLE_SEGMENT|1406,1424|false|false|false|C0587246|Muscle weakness of limb|extremity weakness
Event|Event|SIMPLE_SEGMENT|1416,1424|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1416,1424|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|1429,1437|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|1429,1437|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1429,1437|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|1453,1457|false|false|false|||gone
Event|Event|SIMPLE_SEGMENT|1472,1478|false|false|false|||thinks
Finding|Intellectual Product|SIMPLE_SEGMENT|1484,1491|false|false|false|C0282416|Overall Publication Type|overall
Event|Event|SIMPLE_SEGMENT|1502,1510|false|false|false|||worsened
Event|Event|SIMPLE_SEGMENT|1526,1532|true|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1537,1543|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1537,1543|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1544,1550|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1544,1550|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1555,1564|true|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|1555,1564|true|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|1569,1576|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1569,1576|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1580,1586|true|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|1580,1586|true|false|false|C0042789|Vision|vision
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1589,1592|true|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|1593,1601|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1593,1601|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|1605,1612|false|false|false|||trouble
Finding|Intellectual Product|SIMPLE_SEGMENT|1605,1630|false|false|false|C3827765|Trouble with Coordination|trouble with coordination
Event|Event|SIMPLE_SEGMENT|1618,1630|false|false|false|||coordination
Finding|Functional Concept|SIMPLE_SEGMENT|1618,1630|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|1618,1630|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|1618,1630|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Drug|Organic Chemical|SIMPLE_SEGMENT|1634,1641|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1634,1641|false|false|false|C4319618|Balance (substance)|balance
Event|Event|SIMPLE_SEGMENT|1634,1641|false|false|false|||balance
Finding|Finding|SIMPLE_SEGMENT|1634,1641|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|SIMPLE_SEGMENT|1634,1641|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1634,1641|false|false|false|C2174421|examination of balance|balance
Event|Event|SIMPLE_SEGMENT|1648,1654|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1655,1664|true|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1655,1674|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|1655,1674|true|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|SIMPLE_SEGMENT|1668,1674|true|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|1668,1674|true|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1676,1681|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1676,1681|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1676,1686|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1676,1686|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1682,1686|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1682,1686|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1682,1686|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1682,1686|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1682,1697|true|false|false|C0000737|Abdominal Pain|pain, abdominal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1688,1697|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1688,1702|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1698,1702|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1698,1702|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1698,1702|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1698,1702|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1707,1727|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1712,1719|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1712,1719|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1712,1719|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1712,1719|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1712,1719|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1712,1727|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1720,1727|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1720,1727|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1720,1727|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1729,1747|false|false|false|C0026769|Multiple Sclerosis|Multiple sclerosis
Event|Event|SIMPLE_SEGMENT|1738,1747|false|false|false|||sclerosis
Finding|Pathologic Function|SIMPLE_SEGMENT|1738,1747|false|false|false|C0036429|Sclerosis|sclerosis
Finding|Functional Concept|SIMPLE_SEGMENT|1750,1756|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1750,1764|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1757,1764|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1757,1764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1757,1764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1757,1764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1770,1776|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1770,1776|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1770,1776|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1770,1776|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1770,1784|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1777,1784|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1777,1784|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1777,1784|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1777,1784|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1786,1792|false|false|false|||Mother
Finding|Idea or Concept|SIMPLE_SEGMENT|1786,1792|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1798,1808|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1798,1808|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|SIMPLE_SEGMENT|1798,1808|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1798,1808|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1798,1815|false|false|false|C0235974;C0346647|Malignant neoplasm of pancreas;Pancreatic carcinoma|pancreatic cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1809,1815|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1809,1815|false|false|false|||cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|1817,1824|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|SIMPLE_SEGMENT|1817,1824|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1825,1829|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1825,1829|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1825,1829|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1825,1829|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1825,1836|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1830,1836|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1830,1836|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1856,1861|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1856,1861|false|false|false|C0006111|Brain Diseases|brain
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1856,1868|false|false|false|C0006118;C0153633|Brain Neoplasms;Malignant neoplasm of brain|brain cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1862,1868|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1862,1868|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1873,1881|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1873,1881|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1873,1881|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1873,1881|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1873,1886|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1873,1886|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1882,1886|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1882,1886|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1882,1886|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|1888,1896|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1888,1896|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1888,1896|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1888,1908|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|1888,1908|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|1897,1908|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|1897,1908|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|1897,1908|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|1912,1921|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Classification|SIMPLE_SEGMENT|1923,1930|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|1923,1930|false|false|false|C3812897|General medical service|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|1923,1944|false|false|false|C0031809|Physical Examination|General Physical Exam
Event|Event|SIMPLE_SEGMENT|1931,1939|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1931,1939|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1931,1939|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1931,1939|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1931,1944|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1931,1944|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1940,1944|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1940,1944|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1940,1944|false|false|false|C0582103|Medical Examination|Exam
Finding|Classification|SIMPLE_SEGMENT|1946,1953|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|1946,1953|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|1964,1975|true|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1964,1975|true|true|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1976,1981|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1984,1987|true|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1984,1987|true|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|1984,1987|true|false|false|||MMM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1992,1999|true|false|false|C0036410|Sclera|scleral
Finding|Finding|SIMPLE_SEGMENT|1992,2007|true|false|false|C0240962|Scleral icterus|scleral icterus
Event|Event|SIMPLE_SEGMENT|2000,2007|true|false|false|||icterus
Finding|Sign or Symptom|SIMPLE_SEGMENT|2000,2007|true|false|false|C0022346|Icterus|icterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2012,2021|true|false|false|C0015300|Exophthalmos|proptosis
Event|Event|SIMPLE_SEGMENT|2012,2021|true|false|false|||proptosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2023,2029|true|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2023,2029|true|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|2023,2029|true|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2023,2029|true|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2034,2045|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2034,2045|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2034,2045|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|SIMPLE_SEGMENT|2034,2045|true|false|false|||conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|2034,2045|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|2034,2045|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|2034,2045|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2054,2059|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2054,2059|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2054,2059|true|false|false|C0013604|Edema|edema
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2060,2069|true|false|false|C1272883|Injection|injection
Event|Event|SIMPLE_SEGMENT|2060,2069|true|false|false|||injection
Finding|Functional Concept|SIMPLE_SEGMENT|2060,2069|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2060,2069|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2071,2075|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2071,2075|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|2071,2075|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|2079,2085|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|2079,2085|false|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|2092,2095|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2100,2107|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2100,2107|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2109,2113|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2109,2113|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2118,2125|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2130,2137|true|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|SIMPLE_SEGMENT|2130,2144|true|false|false|C0007280|Carotid bruit|carotid bruits
Event|Event|SIMPLE_SEGMENT|2138,2144|true|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|2138,2144|true|false|false|C0006318|Bruit|bruits
Event|Event|SIMPLE_SEGMENT|2145,2149|true|false|false|||Pulm
Procedure|Health Care Activity|SIMPLE_SEGMENT|2145,2149|true|false|false|C1315068|Pulmonary ventilator management|Pulm
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2152,2155|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|2152,2155|true|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2152,2155|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2152,2155|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2160,2163|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2160,2163|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2166,2170|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2166,2170|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2191,2196|true|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2191,2203|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|2197,2203|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2197,2203|true|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2204,2215|true|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Event|Event|SIMPLE_SEGMENT|2221,2229|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2221,2229|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2234,2239|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2234,2239|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2234,2239|true|false|false|C0013604|Edema|edema
Anatomy|Body System|SIMPLE_SEGMENT|2240,2244|true|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2240,2244|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2240,2244|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|2240,2244|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2240,2244|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Finding|SIMPLE_SEGMENT|2247,2251|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2247,2251|true|false|false|C0687712|warming process|warm
Event|Event|SIMPLE_SEGMENT|2269,2275|true|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2269,2275|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|2287,2291|true|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2287,2291|true|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2287,2291|true|false|false|C0582103|Medical Examination|Exam
Finding|Mental Process|SIMPLE_SEGMENT|2293,2299|false|false|false|C0229992|Psyche structure|MENTAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2293,2306|false|false|false|C0488568;C0488569||MENTAL STATUS
Finding|Finding|SIMPLE_SEGMENT|2293,2306|false|false|false|C0278060|Mental state|MENTAL STATUS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2300,2306|false|false|false|C5889824||STATUS
Event|Event|SIMPLE_SEGMENT|2300,2306|false|false|false|||STATUS
Finding|Idea or Concept|SIMPLE_SEGMENT|2300,2306|false|false|false|C1546481|What subject filter - Status|STATUS
Event|Event|SIMPLE_SEGMENT|2308,2313|false|false|false|||Awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2318,2323|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2318,2323|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2318,2323|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2318,2323|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2318,2323|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2318,2323|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2318,2323|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|2325,2333|false|false|false|||oriented
Finding|Finding|SIMPLE_SEGMENT|2325,2333|false|false|false|C1961028|Oriented to place|oriented
Event|Event|SIMPLE_SEGMENT|2362,2370|false|false|false|||commands
Event|Event|SIMPLE_SEGMENT|2377,2382|false|false|false|||cross
Anatomy|Cell Component|SIMPLE_SEGMENT|2387,2394|false|false|false|C1660780|midline cell component|midline
Event|Event|SIMPLE_SEGMENT|2396,2401|false|false|false|||Knows
Finding|Pathologic Function|SIMPLE_SEGMENT|2413,2420|false|false|false|C5441917|Distant Metastasis|distant
Event|Event|SIMPLE_SEGMENT|2421,2427|false|false|false|||events
Event|Event|SIMPLE_SEGMENT|2421,2427|false|false|false|C0441471|Event|events
Event|Event|SIMPLE_SEGMENT|2432,2443|true|false|false|||hemisensory
Finding|Functional Concept|SIMPLE_SEGMENT|2447,2453|true|false|false|C0234621|Visual|visual
Finding|Finding|SIMPLE_SEGMENT|2447,2461|true|false|false|C0423000|Visual neglect|visual neglect
Event|Event|SIMPLE_SEGMENT|2454,2461|true|false|false|||neglect
Event|Event|SIMPLE_SEGMENT|2454,2461|true|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|SIMPLE_SEGMENT|2454,2461|true|false|false|C0521874|Victim of neglect (finding)|neglect
Finding|Finding|SIMPLE_SEGMENT|2464,2472|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2464,2472|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2464,2472|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2464,2484|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2464,2484|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|2473,2484|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|2473,2484|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2473,2484|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Finding|Body Substance|SIMPLE_SEGMENT|2488,2497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2488,2497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2488,2497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2488,2497|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2527,2530|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|2527,2530|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2527,2530|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|2527,2530|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2527,2536|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI Brain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2531,2536|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2531,2536|false|false|false|C0006111|Brain Diseases|Brain
Event|Event|SIMPLE_SEGMENT|2531,2536|false|false|false|||Brain
Finding|Functional Concept|SIMPLE_SEGMENT|2551,2559|false|false|false|C0032074;C1301732|Planned|Planning
Finding|Mental Process|SIMPLE_SEGMENT|2551,2559|false|false|false|C0032074;C1301732|Planned|Planning
Finding|Finding|SIMPLE_SEGMENT|2565,2573|false|false|false|C0392756|Reduced|Decrease
Finding|Functional Concept|SIMPLE_SEGMENT|2591,2596|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2605,2611|false|false|false|C0230003|Vertex|vertex
Finding|Conceptual Entity|SIMPLE_SEGMENT|2605,2611|false|false|false|C2697524|Graph Node|vertex
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2612,2615|false|false|false|C1308727|RBBP8 protein, human|rim
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2612,2615|false|false|false|C1308727|RBBP8 protein, human|rim
Event|Event|SIMPLE_SEGMENT|2612,2615|false|false|false|||rim
Finding|Gene or Genome|SIMPLE_SEGMENT|2612,2615|false|false|false|C1419293;C1424873;C2347743;C5575294|RBBP8 gene;RBBP8 wt Allele;RIMS1 gene;RIMS1 wt Allele|rim
Event|Event|SIMPLE_SEGMENT|2616,2625|false|false|false|||enhancing
Event|Event|SIMPLE_SEGMENT|2627,2633|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|2627,2633|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|2627,2633|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Finding|SIMPLE_SEGMENT|2639,2648|false|false|false|C0442739||unchanged
Finding|Finding|SIMPLE_SEGMENT|2649,2664|false|false|false|C2825502|Vasogenic Edema|vasogenic edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2659,2664|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2659,2664|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2659,2664|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|2669,2673|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|2669,2673|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|2669,2673|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|2669,2680|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|2674,2680|false|false|false|||effect
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2696,2700|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2696,2700|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2696,2700|false|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2696,2700|false|false|false|C0876917|Procedure on head|Head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2696,2703|false|false|false|C0202691|CAT scan of head|Head CT
Event|Event|SIMPLE_SEGMENT|2701,2703|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|2717,2721|false|false|false|||SCAN
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2717,2721|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|SCAN
Event|Event|SIMPLE_SEGMENT|2723,2733|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|2723,2733|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|2723,2733|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2737,2743|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|2737,2743|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|2737,2743|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|2754,2759|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2769,2775|true|false|false|C0230003|Vertex|vertex
Finding|Conceptual Entity|SIMPLE_SEGMENT|2769,2775|true|false|false|C2697524|Graph Node|vertex
Event|Event|SIMPLE_SEGMENT|2776,2786|true|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2776,2786|true|false|false|C0010280|Craniotomy|craniotomy
Event|Event|SIMPLE_SEGMENT|2796,2804|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|2796,2804|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|2796,2807|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|2808,2818|true|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|2808,2818|true|false|false|C0019080|Hemorrhage|hemorrhage
Finding|Intellectual Product|SIMPLE_SEGMENT|2821,2827|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Finding|SIMPLE_SEGMENT|2828,2843|false|false|false|C2825502|Vasogenic Edema|vasogenic edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2838,2843|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2838,2843|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2838,2843|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2844,2853|false|false|false|||extending
Finding|Functional Concept|SIMPLE_SEGMENT|2862,2867|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2868,2894|false|false|false|C0546003|Frontal and parietal lobes|frontal and parietal lobes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2880,2894|false|false|false|C0030560|Parietal Lobe|parietal lobes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2889,2894|false|false|false|C0796494|lobe|lobes
Finding|Intellectual Product|SIMPLE_SEGMENT|2900,2905|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|2906,2914|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2906,2921|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|2906,2921|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|2954,2962|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|2970,2982|false|false|false|||neurosurgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2970,2982|false|false|false|C0524850|Neurosurgical Procedures|neurosurgery
Event|Occupational Activity|SIMPLE_SEGMENT|2984,2991|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|2984,2991|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Finding|Idea or Concept|SIMPLE_SEGMENT|2999,3002|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|2999,3002|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|3006,3015|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3006,3015|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3030,3040|false|false|false|C0009450|Communicable Diseases|Infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3042,3049|false|false|false|C0012634|Disease|Disease
Finding|Mental Process|SIMPLE_SEGMENT|3060,3072|false|false|false|C0679106|anticipation|anticipation
Event|Event|SIMPLE_SEGMENT|3077,3087|false|false|false|||evacuation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3077,3087|false|false|false|C1282573|Evacuation procedure|evacuation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3095,3100|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3095,3100|false|false|false|C0006111|Brain Diseases|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3102,3109|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|3102,3109|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|3102,3109|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|3127,3130|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|3127,3130|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3127,3130|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|3127,3130|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Finding|SIMPLE_SEGMENT|3131,3144|false|false|false|C0455610|History of surgery|prior surgery
Event|Event|SIMPLE_SEGMENT|3137,3144|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|3137,3144|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|3137,3144|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|3137,3144|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3137,3144|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|3160,3168|false|false|false|||planning
Finding|Functional Concept|SIMPLE_SEGMENT|3160,3168|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|SIMPLE_SEGMENT|3160,3168|false|false|false|C0032074;C1301732|Planned|planning
Finding|Functional Concept|SIMPLE_SEGMENT|3186,3191|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|3192,3202|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3192,3202|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|SIMPLE_SEGMENT|3207,3217|false|false|false|||evacuation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3207,3217|false|false|false|C1282573|Evacuation procedure|evacuation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3222,3229|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|3222,3229|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|3222,3229|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|3242,3251|false|false|false|||tolerated
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3256,3265|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|3256,3265|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|3256,3265|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|3256,3265|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3256,3265|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|SIMPLE_SEGMENT|3266,3270|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3280,3289|false|false|false|||extubated
Finding|Finding|SIMPLE_SEGMENT|3297,3306|false|false|false|C4738506|Operating|operating
Finding|Intellectual Product|SIMPLE_SEGMENT|3321,3325|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|3326,3337|false|false|false|||transferred
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3346,3349|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Event|Event|SIMPLE_SEGMENT|3346,3349|false|false|false|||ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|3346,3349|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Activity|SIMPLE_SEGMENT|3354,3362|false|false|false|C0237820||recovery
Event|Event|SIMPLE_SEGMENT|3354,3362|false|false|false|||recovery
Finding|Organism Function|SIMPLE_SEGMENT|3354,3362|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|SIMPLE_SEGMENT|3395,3408|false|false|false|||non-contrasat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3410,3414|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3410,3414|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3410,3414|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|3410,3414|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3410,3414|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3410,3417|false|false|false|C0202691|CAT scan of head|head CT
Event|Event|SIMPLE_SEGMENT|3424,3432|true|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|3433,3439|true|false|false|||normal
Finding|Finding|SIMPLE_SEGMENT|3440,3454|true|false|false|C0241311|post operative (finding)|post operative
Event|Event|SIMPLE_SEGMENT|3455,3462|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3455,3462|true|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|3470,3473|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|3470,3473|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|3475,3485|true|false|false|||hemorrahge
Event|Event|SIMPLE_SEGMENT|3505,3512|false|false|false|||sitting
Event|Event|SIMPLE_SEGMENT|3563,3569|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3563,3569|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3575,3585|false|false|false|||transfered
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3593,3598|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|3602,3608|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|3602,3608|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|3610,3620|false|false|false|||conditions
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3649,3659|false|false|false|C0009450|Communicable Diseases|Infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3649,3667|false|false|false|C0009450|Communicable Diseases|Infectious Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3660,3667|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|3660,3667|false|false|false|||Disease
Event|Event|SIMPLE_SEGMENT|3676,3687|false|false|false|||recommended
Finding|Body Substance|SIMPLE_SEGMENT|3697,3704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3697,3704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3697,3704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|3708,3715|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3719,3729|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|3719,3729|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|3719,3729|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3719,3729|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|3735,3744|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|SIMPLE_SEGMENT|3735,3744|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|SIMPLE_SEGMENT|3735,3744|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Event|Event|SIMPLE_SEGMENT|3735,3744|false|false|false|||meropenem
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3751,3758|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|3751,3758|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|3751,3758|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|3751,3758|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3751,3758|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|3759,3763|false|false|false|||data
Finding|Idea or Concept|SIMPLE_SEGMENT|3759,3763|false|false|false|C1511726|Data|data
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3773,3777|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3773,3777|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3773,3777|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3773,3777|false|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3778,3783|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|3778,3783|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|3778,3783|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|3778,3783|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|3778,3783|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|3788,3796|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|3809,3817|true|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|3809,3817|true|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|3818,3826|true|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|3830,3836|true|false|false|||growth
Finding|Finding|SIMPLE_SEGMENT|3830,3836|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3830,3836|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|SIMPLE_SEGMENT|3830,3836|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|SIMPLE_SEGMENT|3830,3836|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3830,3836|true|false|false|C2911660|Growth action|growth
Finding|Body Substance|SIMPLE_SEGMENT|3842,3849|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3842,3849|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3842,3849|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|3854,3863|false|false|false|||continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3868,3878|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|3868,3878|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|3868,3878|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3868,3878|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|3880,3889|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|SIMPLE_SEGMENT|3880,3889|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|SIMPLE_SEGMENT|3880,3889|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Event|Event|SIMPLE_SEGMENT|3880,3889|false|false|false|||meropenem
Event|Event|SIMPLE_SEGMENT|3894,3901|false|false|false|||changed
Event|Event|SIMPLE_SEGMENT|3905,3914|false|false|false|||ertapenum
Finding|Body Substance|SIMPLE_SEGMENT|3921,3928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3921,3928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3921,3928|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|3929,3938|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|3942,3950|false|false|false|||progress
Finding|Finding|SIMPLE_SEGMENT|3951,3955|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3974,3978|false|false|false|||some
Finding|Functional Concept|SIMPLE_SEGMENT|3989,3993|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|4000,4008|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4000,4008|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|4020,4030|false|false|false|||complained
Finding|Functional Concept|SIMPLE_SEGMENT|4040,4044|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|4052,4060|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|4052,4060|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4052,4060|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4065,4069|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4065,4069|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4065,4069|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4065,4069|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|4086,4093|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4086,4093|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4086,4093|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4103,4107|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4103,4107|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4103,4107|true|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|4103,4107|true|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4103,4107|true|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4125,4133|true|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|4125,4133|true|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|4145,4148|true|false|false|||DWI
Finding|Individual Behavior|SIMPLE_SEGMENT|4145,4148|true|false|false|C1171335|Driving While Intoxicated|DWI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4145,4148|true|false|false|C0598801|Diffusion weighted imaging|DWI
Event|Event|SIMPLE_SEGMENT|4156,4162|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|4163,4169|false|false|false|C5202796|Intensity and Distress 1|slight
Event|Event|SIMPLE_SEGMENT|4170,4181|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|4170,4181|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|4192,4202|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|4203,4207|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|4203,4207|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4203,4207|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4203,4207|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|4232,4238|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|4232,4238|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|4232,4238|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|4232,4241|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|4232,4241|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|4239,4241|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|4252,4261|false|false|false|||questions
Event|Event|SIMPLE_SEGMENT|4267,4275|false|false|false|||answered
Event|Event|SIMPLE_SEGMENT|4283,4292|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4283,4292|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4283,4292|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4283,4292|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4283,4292|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4296,4307|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4296,4307|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|4296,4307|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4296,4307|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|4296,4320|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|4311,4320|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4311,4320|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4339,4349|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|4339,4349|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|4339,4354|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|4350,4354|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|4350,4354|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|4358,4366|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|4371,4379|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4371,4379|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|4371,4379|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|4371,4379|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|4371,4379|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|4371,4379|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Antibiotic|SIMPLE_SEGMENT|4384,4395|false|false|false|C0007561|ceftriaxone|CeftriaXONE
Drug|Organic Chemical|SIMPLE_SEGMENT|4384,4395|false|false|false|C0007561|ceftriaxone|CeftriaXONE
Event|Event|SIMPLE_SEGMENT|4404,4408|false|false|false|||Q12H
Drug|Organic Chemical|SIMPLE_SEGMENT|4413,4426|false|false|false|C0025872|metronidazole|MetRONIDAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4413,4426|false|false|false|C0025872|metronidazole|MetRONIDAZOLE
Drug|Organic Chemical|SIMPLE_SEGMENT|4428,4434|false|false|false|C0699678|Flagyl|FLagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4428,4434|false|false|false|C0699678|Flagyl|FLagyl
Event|Event|SIMPLE_SEGMENT|4446,4449|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|4454,4463|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4454,4463|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|SIMPLE_SEGMENT|4454,4463|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4454,4463|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|SIMPLE_SEGMENT|4465,4474|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|4465,4474|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4465,4482|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|SIMPLE_SEGMENT|4475,4482|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|4475,4482|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4475,4482|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4475,4482|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|4497,4500|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4501,4505|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4501,4505|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4501,4505|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4501,4505|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|4510,4523|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4510,4523|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|4510,4523|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4510,4523|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|4542,4545|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4546,4550|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4546,4550|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4546,4550|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4546,4550|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|4555,4568|false|false|false|C0377265|levetiracetam|LeVETiracetam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4555,4568|false|false|false|C0377265|levetiracetam|LeVETiracetam
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4555,4568|false|false|false|C3693636|Measurement of levetiracetam|LeVETiracetam
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4580,4583|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4580,4583|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4580,4583|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|4580,4583|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4580,4583|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|4588,4597|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4588,4597|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4588,4597|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4588,4597|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4588,4597|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4588,4609|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|4588,4609|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4598,4609|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|4598,4609|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|4598,4609|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|4611,4615|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|4611,4615|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|4611,4615|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4611,4615|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|4621,4628|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|4621,4628|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|4631,4639|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|4631,4639|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|4647,4656|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4647,4656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4647,4656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4647,4656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4647,4656|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|4647,4666|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4657,4666|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|4657,4666|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|4657,4666|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4657,4666|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4657,4666|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4668,4673|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4668,4673|false|false|false|C0006111|Brain Diseases|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4668,4681|false|false|false|C0006105;C1510428|Brain Abscess;Cerebral abscess|Brain Abscess
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4674,4681|false|false|false|C0000833|Abscess|Abscess
Event|Event|SIMPLE_SEGMENT|4674,4681|false|false|false|||Abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|4674,4681|false|false|false|C1546533||Abscess
Event|Event|SIMPLE_SEGMENT|4684,4693|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4684,4693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4684,4693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4684,4693|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4684,4693|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4694,4703|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4694,4703|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|4694,4703|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|4694,4703|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|4705,4711|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4705,4718|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|4705,4718|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4712,4718|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4712,4718|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|4720,4725|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4720,4725|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|4730,4738|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|4730,4738|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|4740,4745|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4740,4762|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|4740,4762|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|4749,4762|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|4749,4762|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|4749,4762|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4764,4769|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|4764,4769|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4764,4769|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|4764,4769|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|4764,4769|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|4764,4769|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|4764,4769|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|4774,4785|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|4774,4785|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|4787,4795|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4787,4795|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|4787,4795|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4796,4802|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|4796,4802|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4796,4802|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|4804,4814|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|4804,4814|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|4804,4814|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|4804,4814|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|4804,4814|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|4817,4828|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|4817,4828|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|4817,4828|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|4833,4842|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4833,4842|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4833,4842|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4833,4842|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4833,4842|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4833,4855|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4833,4855|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|4833,4855|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4843,4855|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|4843,4855|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4843,4855|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|4863,4870|false|false|false|||staples
Event|Event|SIMPLE_SEGMENT|4878,4882|false|false|false|||stay
Event|Activity|SIMPLE_SEGMENT|4883,4888|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|SIMPLE_SEGMENT|4883,4888|false|false|false|||clean
Event|Event|SIMPLE_SEGMENT|4912,4919|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|4931,4937|false|false|false|||friend
Finding|Idea or Concept|SIMPLE_SEGMENT|4931,4937|false|false|false|C1546502|Relationship - Friend|friend
Finding|Classification|SIMPLE_SEGMENT|4941,4947|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|4941,4947|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|4941,4947|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|4941,4947|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|4955,4960|false|false|false|||check
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4965,4970|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|4965,4970|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|4965,4970|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|4965,4970|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|4965,4970|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|4975,4980|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|4975,4980|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|4975,4980|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4985,4994|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|4985,4994|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|4985,4994|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5003,5010|false|false|false|C0041834|Erythema|redness
Event|Event|SIMPLE_SEGMENT|5003,5010|false|false|false|||redness
Finding|Finding|SIMPLE_SEGMENT|5003,5010|false|false|false|C0332575|Redness|redness
Event|Event|SIMPLE_SEGMENT|5014,5022|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|5014,5022|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|5014,5022|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5014,5022|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|5032,5036|false|false|false|||Take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5042,5046|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5042,5046|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5042,5046|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5042,5046|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5042,5055|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|SIMPLE_SEGMENT|5042,5055|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5042,5055|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5047,5055|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|SIMPLE_SEGMENT|5047,5055|false|false|false|||medicine
Event|Event|SIMPLE_SEGMENT|5059,5069|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|5073,5079|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|5093,5097|true|false|false|||need
Event|Event|SIMPLE_SEGMENT|5101,5105|true|false|false|||take
Finding|Intellectual Product|SIMPLE_SEGMENT|5123,5132|true|false|false|C2984058|Have Pain|have pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5128,5132|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5128,5132|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5128,5132|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5128,5132|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5135,5143|false|false|false|||Exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5135,5143|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5135,5143|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|SIMPLE_SEGMENT|5154,5161|false|false|false|||limited
Event|Event|SIMPLE_SEGMENT|5165,5172|false|false|false|||walking
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5165,5172|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|SIMPLE_SEGMENT|5165,5172|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|SIMPLE_SEGMENT|5165,5172|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Activity|SIMPLE_SEGMENT|5177,5184|true|false|false|C0206244|Lifting|lifting
Event|Event|SIMPLE_SEGMENT|5177,5184|true|false|false|||lifting
Event|Event|SIMPLE_SEGMENT|5194,5203|true|false|false|||straining
Finding|Physiologic Function|SIMPLE_SEGMENT|5194,5203|true|false|false|C0442694|Straining (finding)|straining
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5218,5225|false|false|false|C0011119|Decompression Sickness|bending
Event|Event|SIMPLE_SEGMENT|5218,5225|false|false|false|||bending
Finding|Finding|SIMPLE_SEGMENT|5218,5225|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|SIMPLE_SEGMENT|5218,5225|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|SIMPLE_SEGMENT|5228,5236|false|false|false|||Increase
Event|Event|SIMPLE_SEGMENT|5242,5248|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|5242,5248|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|5242,5248|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Substance|SIMPLE_SEGMENT|5252,5258|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|5252,5258|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|5252,5258|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5252,5258|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Tissue|SIMPLE_SEGMENT|5263,5268|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|SIMPLE_SEGMENT|5263,5268|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5263,5268|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5273,5281|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5273,5281|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5282,5286|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5282,5286|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5282,5286|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5282,5286|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5288,5296|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|SIMPLE_SEGMENT|5288,5296|false|false|false|||medicine
Event|Event|SIMPLE_SEGMENT|5301,5306|false|false|false|||cause
Event|Event|SIMPLE_SEGMENT|5307,5319|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5307,5319|false|false|false|C0009806|Constipation|constipation
Event|Event|SIMPLE_SEGMENT|5334,5343|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|5344,5350|false|false|false|||taking
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5355,5371|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5364,5371|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|SIMPLE_SEGMENT|5364,5371|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|SIMPLE_SEGMENT|5372,5377|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|5372,5386|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5372,5386|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|SIMPLE_SEGMENT|5378,5386|false|false|false|||softener
Drug|Organic Chemical|SIMPLE_SEGMENT|5396,5404|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5396,5404|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|5406,5412|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5406,5412|false|false|false|C0282139|Colace|Colace
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5428,5436|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5428,5436|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5437,5441|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5437,5441|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5437,5441|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5437,5441|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5442,5452|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|5442,5452|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5442,5452|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|5455,5457|true|false|false|||DO
Event|Event|SIMPLE_SEGMENT|5462,5466|true|false|false|||take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5471,5488|true|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5489,5498|true|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|SIMPLE_SEGMENT|5489,5498|true|false|false|||medicines
Drug|Organic Chemical|SIMPLE_SEGMENT|5507,5513|true|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5507,5513|true|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|SIMPLE_SEGMENT|5516,5523|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5516,5523|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|5525,5530|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5525,5530|false|false|false|C0593507|Advil|Advil
Event|Event|SIMPLE_SEGMENT|5525,5530|false|false|false|||Advil
Finding|Gene or Genome|SIMPLE_SEGMENT|5525,5530|false|false|false|C1422473|AVIL gene|Advil
Drug|Organic Chemical|SIMPLE_SEGMENT|5535,5544|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5535,5544|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Functional Concept|SIMPLE_SEGMENT|5556,5562|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5556,5562|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5556,5565|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5556,5565|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|5563,5565|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|5583,5593|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|5597,5603|false|false|false|C0876060|Keppra|Keppra
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5597,5603|false|false|false|C0876060|Keppra|Keppra
Drug|Organic Chemical|SIMPLE_SEGMENT|5605,5618|false|false|false|C0377265|levetiracetam|Levetiracetam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5605,5618|false|false|false|C0377265|levetiracetam|Levetiracetam
Event|Event|SIMPLE_SEGMENT|5605,5618|false|false|false|||Levetiracetam
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5605,5618|false|false|false|C3693636|Measurement of levetiracetam|Levetiracetam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5638,5646|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|SIMPLE_SEGMENT|5638,5646|false|false|false|||medicine
Event|Event|SIMPLE_SEGMENT|5661,5668|true|false|false|||require
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5669,5674|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5669,5674|true|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5669,5674|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|5675,5679|true|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|5675,5679|true|false|false|C0043227|Work|work
Event|Activity|SIMPLE_SEGMENT|5681,5691|true|false|false|C1283169||monitoring
Event|Event|SIMPLE_SEGMENT|5681,5691|true|false|false|||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|5681,5691|true|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|SIMPLE_SEGMENT|5701,5706|true|false|false|||drive
Event|Event|SIMPLE_SEGMENT|5718,5724|true|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|5718,5724|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5718,5724|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5718,5727|true|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5718,5727|true|false|false|C1522577|follow-up|follow up
Event|Activity|SIMPLE_SEGMENT|5728,5739|true|false|false|C0003629|Appointments|appointment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5744,5752|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5753,5765|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|5753,5765|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5753,5765|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

