 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
.|12,13
Unit|23,27
No|28,30
:|30,31
_|34,35
_|35,36
_|36,37
<EOL>|37,38
<EOL>|39,40
Admission|40,49
Date|50,54
:|54,55
_|57,58
_|58,59
_|59,60
Discharge|74,83
Date|84,88
:|88,89
_|92,93
_|93,94
_|94,95
<EOL>|95,96
<EOL>|97,98
Date|98,102
of|103,105
Birth|106,111
:|111,112
_|114,115
_|115,116
_|116,117
Sex|130,133
:|133,134
F|137,138
<EOL>|138,139
<EOL>|140,141
Service|141,148
:|148,149
MEDICINE|150,158
<EOL>|158,159
<EOL>|160,161
Allergies|161,170
:|170,171
<EOL>|172,173
Patient|173,180
recorded|181,189
as|190,192
having|193,199
No|200,202
Known|203,208
Allergies|209,218
to|219,221
Drugs|222,227
<EOL>|227,228
<EOL>|229,230
Attending|230,239
:|239,240
_|241,242
_|242,243
_|243,244
.|244,245
<EOL>|245,246
<EOL>|247,248
Chief|248,253
Complaint|254,263
:|263,264
<EOL>|264,265
Abdominal|265,274
distention|275,285
/|285,286
pain|286,290
and|291,294
fever|295,300
<EOL>|300,301
<EOL>|302,303
Major|303,308
Surgical|309,317
or|318,320
Invasive|321,329
Procedure|330,339
:|339,340
<EOL>|340,341
Paracentesis|341,353
_|354,355
_|355,356
_|356,357
(|358,359
diagnostic|359,369
)|369,370
and|371,374
_|375,376
_|376,377
_|377,378
(|379,380
therapeutic|380,391
)|391,392
<EOL>|392,393
<EOL>|393,394
<EOL>|395,396
History|396,403
of|404,406
Present|407,414
Illness|415,422
:|422,423
<EOL>|423,424
_|424,425
_|425,426
_|426,427
with|428,432
recently|433,441
diagnosed|442,451
alcoholic|452,461
hepatitis|462,471
,|471,472
persistent|473,483
<EOL>|484,485
ascites|485,492
,|492,493
and|494,497
persistent|498,508
fevers|509,515
and|516,519
leukocytosis|520,532
which|533,538
have|539,543
been|544,548
<EOL>|549,550
atributed|550,559
to|560,562
her|563,566
hepatitis|567,576
who|577,580
presented|581,590
to|591,593
_|594,595
_|595,596
_|596,597
today|598,603
with|604,608
<EOL>|609,610
worsening|610,619
abdominal|620,629
distention|630,640
,|640,641
pain|642,646
,|646,647
and|648,651
persistent|652,662
fever|663,668
.|668,669
She|670,673
<EOL>|674,675
denies|675,681
chills|682,688
but|689,692
did|693,696
have|697,701
sweats|702,708
the|709,712
night|713,718
prior|719,724
to|725,727
admission|728,737
.|737,738
<EOL>|739,740
She|740,743
has|744,747
tried|748,753
to|754,756
be|757,759
strictly|760,768
compliant|769,778
with|779,783
her|784,787
low|788,791
socium|792,798
diet|799,803
<EOL>|804,805
and|805,808
fluid|809,814
restriction|815,826
,|826,827
and|828,831
denies|832,838
any|839,842
increased|843,852
fluid|853,858
or|859,861
sodium|862,868
<EOL>|869,870
intake|870,876
.|876,877
She|878,881
reports|882,889
sobriety|890,898
from|899,903
alcohol|904,911
since|912,917
_|918,919
_|919,920
_|920,921
.|921,922
At|923,925
_|926,927
_|927,928
_|928,929
<EOL>|930,931
she|931,934
was|935,938
febrile|939,946
and|947,950
tender|951,957
to|958,960
palpation|961,970
,|970,971
so|972,974
she|975,978
was|979,982
referred|983,991
to|992,994
<EOL>|995,996
the|996,999
ED|1000,1002
.|1002,1003
<EOL>|1005,1006
.|1006,1007
<EOL>|1009,1010
In|1010,1012
the|1013,1016
ED|1017,1019
initial|1020,1027
vital|1028,1033
signs|1034,1039
were|1040,1044
99.0|1045,1049
113|1050,1053
/|1053,1054
72|1054,1056
132|1057,1060
16|1061,1063
99|1064,1066
%|1066,1067
on|1068,1070
RA|1071,1073
.|1073,1074
<EOL>|1075,1076
Her|1076,1079
temp|1080,1084
increased|1085,1094
to|1095,1097
100.4|1098,1103
and|1104,1107
her|1108,1111
pulse|1112,1117
came|1118,1122
down|1123,1127
to|1128,1130
the|1131,1134
100s|1135,1139
<EOL>|1140,1141
with|1141,1145
Ativan|1146,1152
.|1152,1153
She|1154,1157
received|1158,1166
morphine|1167,1175
4mg|1176,1179
IV|1180,1182
x|1183,1184
4|1185,1186
for|1187,1190
pain|1191,1195
,|1195,1196
tylenol|1197,1204
<EOL>|1205,1206
_|1206,1207
_|1207,1208
_|1208,1209
PO|1210,1212
x1|1213,1215
for|1216,1219
fever|1220,1225
,|1225,1226
ondansetron|1227,1238
4mg|1239,1242
IV|1243,1245
x2|1246,1248
for|1249,1252
nausea|1253,1259
,|1259,1260
and|1261,1264
<EOL>|1265,1266
lorazeman|1266,1275
0.5|1276,1279
mg|1279,1281
IV|1282,1284
x1|1285,1287
for|1288,1291
anxiety|1292,1299
.|1299,1300
She|1301,1304
underwent|1305,1314
a|1315,1316
diagnostic|1317,1327
<EOL>|1328,1329
paracentesis|1329,1341
but|1342,1345
the|1346,1349
samples|1350,1357
were|1358,1362
initially|1363,1372
lost|1373,1377
.|1377,1378
She|1379,1382
was|1383,1386
<EOL>|1387,1388
treated|1388,1395
with|1396,1400
ceftriaxone|1401,1412
2g|1413,1415
IV|1416,1418
x1|1419,1421
for|1422,1425
possible|1426,1434
SBP|1435,1438
.|1438,1439
She|1440,1443
was|1444,1447
<EOL>|1448,1449
admitted|1449,1457
to|1458,1460
Medicine|1461,1469
for|1470,1473
further|1474,1481
management|1482,1492
.|1492,1493
Fortunately|1494,1505
,|1505,1506
her|1507,1510
<EOL>|1511,1512
samples|1512,1519
were|1520,1524
found|1525,1530
after|1531,1536
she|1537,1540
arrived|1541,1548
on|1549,1551
the|1552,1555
floor|1556,1561
.|1561,1562
<EOL>|1564,1565
.|1565,1566
<EOL>|1568,1569
On|1569,1571
the|1572,1575
floor|1576,1581
her|1582,1585
mood|1586,1590
is|1591,1593
labile|1594,1600
.|1600,1601
She|1602,1605
is|1606,1608
at|1609,1611
times|1612,1617
tearful|1618,1625
and|1626,1629
at|1630,1632
<EOL>|1633,1634
times|1634,1639
pleasant|1640,1648
.|1648,1649
She|1650,1653
does|1654,1658
seem|1659,1663
uncomfortable|1664,1677
.|1677,1678
She|1679,1682
is|1683,1685
not|1686,1689
confused|1690,1698
<EOL>|1699,1700
or|1700,1702
obviously|1703,1712
encephalopathic|1713,1728
.|1728,1729
She|1730,1733
denies|1734,1740
cough|1741,1746
,|1746,1747
dysuria|1748,1755
,|1755,1756
<EOL>|1757,1758
diarrhea|1758,1766
,|1766,1767
or|1768,1770
rash|1771,1775
.|1775,1776
She|1777,1780
does|1781,1785
endorse|1786,1793
decreased|1794,1803
UOP|1804,1807
for|1808,1811
the|1812,1815
past|1816,1820
<EOL>|1821,1822
few|1822,1825
days|1826,1830
.|1830,1831
<EOL>|1833,1834
.|1834,1835
<EOL>|1835,1836
Review|1836,1842
of|1843,1845
Systems|1846,1853
:|1853,1854
<EOL>|1856,1857
(|1857,1858
+|1858,1859
)|1859,1860
Per|1861,1864
HPI|1865,1868
<EOL>|1870,1871
(|1871,1872
-|1872,1873
)|1873,1874
Denies|1875,1881
chills|1882,1888
.|1888,1889
Denies|1890,1896
headache|1897,1905
,|1905,1906
sinus|1907,1912
tenderness|1913,1923
,|1923,1924
rhinorrhea|1925,1935
<EOL>|1936,1937
or|1937,1939
congestion|1940,1950
.|1950,1951
Denies|1952,1958
chest|1959,1964
pain|1965,1969
or|1970,1972
tightness|1973,1982
,|1982,1983
palpitations|1984,1996
.|1996,1997
<EOL>|1998,1999
Denies|1999,2005
cough|2006,2011
,|2011,2012
shortness|2013,2022
of|2023,2025
breath|2026,2032
,|2032,2033
or|2034,2036
wheezes|2037,2044
.|2044,2045
Denied|2046,2052
nausea|2053,2059
,|2059,2060
<EOL>|2061,2062
vomiting|2062,2070
,|2070,2071
diarrhea|2072,2080
,|2080,2081
constipation|2082,2094
.|2094,2095
No|2096,2098
recent|2099,2105
change|2106,2112
in|2113,2115
bowel|2116,2121
or|2122,2124
<EOL>|2125,2126
bladder|2126,2133
habits|2134,2140
.|2140,2141
No|2142,2144
dysuria|2145,2152
.|2152,2153
Denies|2154,2160
arthralgias|2161,2172
or|2173,2175
myalgias|2176,2184
.|2184,2185
<EOL>|2186,2187
Denies|2187,2193
rashes|2194,2200
or|2201,2203
skin|2204,2208
breakdown|2209,2218
.|2218,2219
No|2220,2222
numbness|2223,2231
/|2231,2232
tingling|2232,2240
in|2241,2243
<EOL>|2244,2245
extremities|2245,2256
.|2256,2257
No|2258,2260
feelings|2261,2269
of|2270,2272
depression|2273,2283
or|2284,2286
anxiety|2287,2294
.|2294,2295
All|2296,2299
other|2300,2305
<EOL>|2306,2307
review|2307,2313
of|2314,2316
systems|2317,2324
negative|2325,2333
.|2333,2334
<EOL>|2336,2337
<EOL>|2337,2338
<EOL>|2339,2340
Past|2340,2344
Medical|2345,2352
History|2353,2360
:|2360,2361
<EOL>|2361,2362
-|2362,2363
Alcohol|2364,2371
abuse|2372,2377
<EOL>|2379,2380
-|2380,2381
Alcoholic|2382,2391
hepatitis|2392,2401
,|2401,2402
with|2403,2407
persistent|2408,2418
fever|2419,2424
and|2425,2428
leukocytosis|2429,2441
<EOL>|2441,2442
-|2442,2443
Ascites|2444,2451
<EOL>|2452,2453
-|2453,2454
Chronic|2455,2462
back|2463,2467
pain|2468,2472
<EOL>|2473,2474
<EOL>|2475,2476
Social|2476,2482
History|2483,2490
:|2490,2491
<EOL>|2491,2492
_|2492,2493
_|2493,2494
_|2494,2495
<EOL>|2495,2496
Family|2496,2502
History|2503,2510
:|2510,2511
<EOL>|2511,2512
-|2512,2513
Mother|2514,2520
:|2520,2521
_|2522,2523
_|2523,2524
_|2524,2525
cancer|2526,2532
,|2532,2533
age|2534,2537
_|2538,2539
_|2539,2540
_|2540,2541
<EOL>|2543,2544
-|2544,2545
No|2546,2548
family|2549,2555
history|2556,2563
of|2564,2566
liver|2567,2572
disease|2573,2580
<EOL>|2582,2583
-|2583,2584
Multiple|2585,2593
relatives|2594,2603
with|2604,2608
alcoholism|2609,2619
<EOL>|2621,2622
<EOL>|2623,2624
Physical|2624,2632
Exam|2633,2637
:|2637,2638
<EOL>|2638,2639
Physical|2639,2647
Exam|2648,2652
on|2653,2655
Admission|2656,2665
:|2665,2666
<EOL>|2668,2669
GEN|2669,2672
:|2672,2673
NAD|2674,2677
,|2677,2678
labile|2679,2685
affect|2686,2692
between|2693,2700
pleasant|2701,2709
and|2710,2713
tearful|2714,2721
<EOL>|2723,2724
VS|2724,2726
:|2726,2727
101.0|2728,2733
104|2734,2737
/|2737,2738
69|2738,2740
125|2741,2744
18|2745,2747
95|2748,2750
%|2750,2751
on|2752,2754
RA|2755,2757
<EOL>|2759,2760
HEENT|2760,2765
:|2765,2766
Dry|2767,2770
MM|2771,2773
,|2773,2774
no|2775,2777
OP|2778,2780
lesions|2781,2788
,|2788,2789
mild|2790,2794
scleral|2795,2802
icterus|2803,2810
<EOL>|2812,2813
CV|2813,2815
:|2815,2816
RR|2817,2819
,|2819,2820
tachy|2821,2826
,|2826,2827
no|2828,2830
MRG|2831,2834
<EOL>|2836,2837
PULM|2837,2841
:|2841,2842
Bibasilar|2843,2852
crackles|2853,2861
R|2862,2863
>|2864,2865
L|2866,2867
<EOL>|2869,2870
ABD|2870,2873
:|2873,2874
BS|2875,2877
+|2877,2878
,|2878,2879
soft|2880,2884
,|2884,2885
distended|2886,2895
,|2895,2896
diffusely|2897,2906
tender|2907,2913
with|2914,2918
mild|2919,2923
rebound|2924,2931
,|2931,2932
<EOL>|2933,2934
obvious|2934,2941
collateral|2942,2952
veins|2953,2958
,|2958,2959
some|2960,2964
mild|2965,2969
angiomata|2970,2979
<EOL>|2981,2982
LIMBS|2982,2987
:|2987,2988
Trace|2989,2994
_|2995,2996
_|2996,2997
_|2997,2998
edema|2999,3004
,|3004,3005
no|3006,3008
tremors|3009,3016
or|3017,3019
asterixis|3020,3029
<EOL>|3031,3032
SKIN|3032,3036
:|3036,3037
No|3038,3040
rashes|3041,3047
or|3048,3050
skin|3051,3055
breakdown|3056,3065
,|3065,3066
scattered|3067,3076
ecchymoses|3077,3087
at|3088,3090
<EOL>|3091,3092
puncture|3092,3100
sites|3101,3106
<EOL>|3108,3109
NEURO|3109,3114
:|3114,3115
A|3116,3117
and|3118,3121
O|3122,3123
x|3124,3125
3|3126,3127
,|3127,3128
no|3129,3131
pronator|3132,3140
drift|3141,3146
,|3146,3147
reflexes|3148,3156
are|3157,3160
1|3161,3162
+|3162,3163
of|3164,3166
the|3167,3170
<EOL>|3171,3172
upper|3172,3177
and|3178,3181
lower|3182,3187
extremities|3188,3199
<EOL>|3201,3202
<EOL>|3203,3204
Pertinent|3204,3213
Results|3214,3221
:|3221,3222
<EOL>|3222,3223
LABS|3223,3227
:|3227,3228
<EOL>|3228,3229
<EOL>|3229,3230
Blood|3230,3235
_|3236,3237
_|3237,3238
_|3238,3239
:|3239,3240
<EOL>|3240,3241
WBC|3241,3244
-|3244,3245
17|3245,3247
.|3247,3248
9|3248,3249
*|3249,3250
RBC|3251,3254
-|3254,3255
3|3255,3256
.|3256,3257
25|3257,3259
*|3259,3260
HGB|3261,3264
-|3264,3265
11|3265,3267
.|3267,3268
0|3268,3269
*|3269,3270
HCT|3271,3274
-|3274,3275
34|3275,3277
.|3277,3278
1|3278,3279
*|3279,3280
MCV|3281,3284
-|3284,3285
105|3285,3288
*|3288,3289
MCH|3290,3293
-|3293,3294
33|3294,3296
.|3296,3297
9|3297,3298
*|3298,3299
<EOL>|3300,3301
MCHC|3301,3305
-|3305,3306
32.3|3306,3310
RDW|3311,3314
-|3314,3315
14.0|3315,3319
PLT|3320,3323
COUNT|3324,3329
-|3329,3330
198|3330,3333
_|3334,3335
_|3335,3336
_|3336,3337
PTT|3338,3341
-|3341,3342
39|3342,3344
.|3344,3345
3|3345,3346
*|3346,3347
_|3348,3349
_|3349,3350
_|3350,3351
<EOL>|3351,3352
ALBUMIN|3352,3359
-|3359,3360
2|3360,3361
.|3361,3362
7|3362,3363
*|3363,3364
ALT|3365,3368
(|3368,3369
SGPT|3369,3373
)|3373,3374
-|3374,3375
33|3375,3377
AST|3378,3381
(|3381,3382
SGOT|3382,3386
)|3386,3387
-|3387,3388
124|3388,3391
*|3391,3392
ALK|3393,3396
PHOS|3397,3401
-|3401,3402
186|3402,3405
*|3405,3406
TOT|3407,3410
<EOL>|3411,3412
BILI|3412,3416
-|3416,3417
2.4|3417,3420
<EOL>|3420,3421
<EOL>|3421,3422
Ascitic|3422,3429
Fluid|3430,3435
_|3436,3437
_|3437,3438
_|3438,3439
:|3439,3440
<EOL>|3442,3443
WBC|3443,3446
-|3446,3447
52|3447,3449
*|3449,3450
RBC|3451,3454
-|3454,3455
98|3455,3457
*|3457,3458
POLYS|3459,3464
-|3464,3465
13|3465,3467
*|3467,3468
LYMPHS|3469,3475
-|3475,3476
20|3476,3478
*|3478,3479
MONOS|3480,3485
-|3485,3486
0|3486,3487
EOS|3488,3491
-|3491,3492
1|3492,3493
*|3493,3494
<EOL>|3495,3496
MESOTHELI|3496,3505
-|3505,3506
16|3506,3508
*|3508,3509
MACROPHAG|3510,3519
-|3519,3520
50|3520,3522
*|3522,3523
<EOL>|3523,3524
TOT|3524,3527
PROT|3528,3532
-|3532,3533
1.1|3533,3536
LD|3537,3539
(|3539,3540
LDH|3540,3543
)|3543,3544
-|3544,3545
42|3545,3547
ALBUMIN|3548,3555
-|3555,3556
<|3556,3557
1.0|3557,3560
<EOL>|3560,3561
<EOL>|3561,3562
Ascitic|3562,3569
Fluid|3570,3575
_|3576,3577
_|3577,3578
_|3578,3579
:|3579,3580
<EOL>|3580,3581
WBC|3581,3584
-|3584,3585
104|3585,3588
*|3588,3589
RBB|3590,3593
-|3593,3594
290|3594,3597
*|3597,3598
POLYS|3599,3604
-|3604,3605
14|3605,3607
*|3607,3608
LYMPHS|3609,3615
-|3615,3616
17|3616,3618
*|3618,3619
MONOS|3620,3625
-|3625,3626
3|3626,3627
*|3627,3628
EOS|3629,3632
-|3632,3633
21|3633,3635
*|3635,3636
<EOL>|3637,3638
MESOTHELI|3638,3647
-|3647,3648
45|3648,3650
*|3650,3651
<EOL>|3652,3653
<EOL>|3653,3654
Blood|3654,3659
_|3660,3661
_|3661,3662
_|3662,3663
:|3663,3664
<EOL>|3664,3665
WBC|3665,3668
-|3668,3669
11.1|3669,3673
HCT|3674,3677
30.7|3678,3682
<EOL>|3682,3683
<EOL>|3684,3685
RADIOLOGY|3685,3694
:|3694,3695
<EOL>|3695,3696
Lumbo|3696,3701
-|3701,3702
sacral|3702,3708
XR|3709,3711
:|3711,3712
Normal|3713,3719
,|3719,3720
no|3721,3723
evidence|3724,3732
of|3733,3735
osteomyelitis|3736,3749
/|3749,3750
vertebral|3750,3759
<EOL>|3760,3761
compression|3761,3772
fracture|3773,3781
.|3781,3782
<EOL>|3782,3783
<EOL>|3783,3784
<EOL>|3785,3786
Brief|3786,3791
Hospital|3792,3800
Course|3801,3807
:|3807,3808
<EOL>|3808,3809
#|3809,3810
Abdominal|3810,3819
distention|3820,3830
/|3830,3831
pain|3831,3835
:|3835,3836
<EOL>|3836,3837
She|3837,3840
was|3841,3844
treated|3845,3852
empirically|3853,3864
due|3865,3868
to|3869,3871
concern|3872,3879
for|3880,3883
spontaneous|3884,3895
<EOL>|3896,3897
bacterial|3897,3906
peritonitis|3907,3918
with|3919,3923
ceftriaxone|3924,3935
2g|3936,3938
x|3939,3940
1|3941,3942
.|3942,3943
A|3945,3946
diagnostic|3947,3957
<EOL>|3958,3959
paracentesis|3959,3971
was|3972,3975
performed|3976,3985
in|3986,3988
the|3989,3992
ED|3993,3995
.|3995,3996
Ascitic|3998,4005
fluid|4006,4011
analysis|4012,4020
<EOL>|4021,4022
was|4022,4025
performed|4026,4035
.|4035,4036
Spontaneous|4038,4049
bacterial|4050,4059
peritonitis|4060,4071
was|4072,4075
ruled|4076,4081
out|4082,4085
<EOL>|4086,4087
given|4087,4092
that|4093,4097
the|4098,4101
fluid|4102,4107
cell|4108,4112
count|4113,4118
showed|4119,4125
only|4126,4130
52|4131,4133
WBC|4134,4137
;|4137,4138
antibiotics|4139,4150
<EOL>|4151,4152
were|4152,4156
discontinued|4157,4169
in|4170,4172
this|4173,4177
setting|4178,4185
.|4185,4186
Subsequently|4188,4200
,|4200,4201
a|4202,4203
large|4204,4209
volume|4210,4216
<EOL>|4217,4218
paracentesis|4218,4230
was|4231,4234
performed|4235,4244
on|4245,4247
_|4248,4249
_|4249,4250
_|4250,4251
with|4252,4256
4.5|4257,4260
L|4260,4261
of|4262,4264
fluids|4265,4271
<EOL>|4272,4273
removed|4273,4280
.|4280,4281
After|4282,4287
the|4288,4291
procedure|4292,4301
,|4301,4302
her|4303,4306
abdomen|4307,4314
was|4315,4318
less|4319,4323
distended|4324,4333
and|4334,4337
<EOL>|4338,4339
less|4339,4343
painful|4344,4351
.|4351,4352
Fluid|4354,4359
analysis|4360,4368
again|4369,4374
did|4375,4378
not|4379,4382
reveal|4383,4389
SBP|4390,4393
.|4393,4394
<EOL>|4396,4397
.|4397,4398
<EOL>|4398,4399
#|4399,4400
Alcoholic|4400,4409
hepatitis|4410,4419
:|4419,4420
<EOL>|4420,4421
Patient|4421,4428
's|4428,4430
liver|4431,4436
synthetic|4437,4446
function|4447,4455
was|4456,4459
monitored|4460,4469
while|4470,4475
<EOL>|4476,4477
hospitalized|4477,4489
.|4489,4490
She|4491,4494
was|4495,4498
maintained|4499,4509
on|4510,4512
her|4513,4516
home|4517,4521
regimen|4522,4529
of|4530,4532
<EOL>|4533,4534
lactulose|4534,4543
.|4543,4544
She|4545,4548
also|4549,4553
had|4554,4557
24|4558,4560
-|4560,4561
hr|4561,4563
urine|4564,4569
collection|4570,4580
for|4581,4584
copper|4585,4591
to|4592,4594
<EOL>|4595,4596
evaluate|4596,4604
for|4605,4608
_|4609,4610
_|4610,4611
_|4611,4612
disease|4613,4620
.|4620,4621
<EOL>|4622,4623
.|4623,4624
<EOL>|4624,4625
#|4625,4626
Leukocytosis|4626,4638
and|4639,4642
mild|4643,4647
fever|4648,4653
:|4653,4654
<EOL>|4654,4655
She|4655,4658
had|4659,4662
a|4663,4664
temparature|4665,4676
of|4677,4679
101|4680,4683
upon|4684,4688
presentation|4689,4701
in|4702,4704
the|4705,4708
ED|4709,4711
.|4711,4712
She|4714,4717
<EOL>|4718,4719
had|4719,4722
no|4723,4725
signs|4726,4731
or|4732,4734
symptoms|4735,4743
of|4744,4746
any|4747,4750
infection|4751,4760
.|4760,4761
Urine|4763,4768
culture|4769,4776
showed|4777,4783
<EOL>|4784,4785
only|4785,4789
GU|4790,4792
flora|4793,4798
,|4798,4799
consistent|4800,4810
with|4811,4815
contamination|4816,4829
.|4829,4830
After|4831,4836
arrival|4837,4844
to|4845,4847
<EOL>|4848,4849
the|4849,4852
floor|4853,4858
her|4859,4862
temperature|4863,4874
was|4875,4878
stable|4879,4885
,|4885,4886
ranging|4887,4894
from|4895,4899
99|4900,4902
to|4903,4905
101|4906,4909
.|4909,4910
<EOL>|4912,4913
Her|4913,4916
WBC|4917,4920
trended|4921,4928
down|4929,4933
throughout|4934,4944
the|4945,4948
hospitalization|4949,4964
and|4965,4968
was|4969,4972
11|4973,4975
<EOL>|4976,4977
at|4977,4979
the|4980,4983
time|4984,4988
of|4989,4991
discharge|4992,5001
.|5001,5002
<EOL>|5006,5007
.|5007,5008
<EOL>|5008,5009
#|5009,5010
Tachycardia|5010,5021
:|5021,5022
<EOL>|5022,5023
Her|5023,5026
heart|5027,5032
rate|5033,5037
was|5038,5041
elevated|5042,5050
in|5051,5053
the|5054,5057
100|5058,5061
-|5061,5062
120s|5062,5066
throughout|5067,5077
the|5078,5081
<EOL>|5082,5083
hospitalization|5083,5098
.|5098,5099
She|5100,5103
had|5104,5107
good|5108,5112
oxygenation|5113,5124
and|5125,5128
had|5129,5132
no|5133,5135
complaints|5136,5146
<EOL>|5147,5148
of|5148,5150
SOB|5151,5154
,|5154,5155
dyspnea|5156,5163
,|5163,5164
chest|5165,5170
pain|5171,5175
,|5175,5176
palpitations|5177,5189
.|5189,5190
The|5191,5194
most|5195,5199
likely|5200,5206
<EOL>|5207,5208
etiology|5208,5216
of|5217,5219
this|5220,5224
is|5225,5227
pain|5228,5232
,|5232,5233
anxiety|5234,5241
,|5241,5242
and|5243,5246
her|5247,5250
low|5251,5254
intravascular|5255,5268
<EOL>|5269,5270
volume|5270,5276
.|5276,5277
She|5279,5282
was|5283,5286
tachycardic|5287,5298
in|5299,5301
the|5302,5305
100s|5306,5310
upon|5311,5315
discharge|5316,5325
.|5325,5326
<EOL>|5328,5329
.|5329,5330
<EOL>|5330,5331
#|5331,5332
Back|5332,5336
pain|5337,5341
:|5341,5342
<EOL>|5342,5343
Lumbosacral|5343,5354
spine|5355,5360
film|5361,5365
revealed|5366,5374
no|5375,5377
skeletal|5378,5386
abnormalities|5387,5400
<EOL>|5401,5402
(|5402,5403
vertebral|5403,5412
compression|5413,5424
fracture|5425,5433
and|5434,5437
osteomyelitis|5438,5451
)|5451,5452
.|5452,5453
Her|5455,5458
pain|5459,5463
<EOL>|5464,5465
was|5465,5468
present|5469,5476
but|5477,5480
well|5481,5485
-|5485,5486
controlled|5486,5496
throughout|5497,5507
the|5508,5511
hospitalization|5512,5527
<EOL>|5528,5529
with|5529,5533
oxycodone|5534,5543
_|5544,5545
_|5545,5546
_|5546,5547
Q6H|5548,5551
PRN|5552,5555
pain|5556,5560
.|5560,5561
Recommended|5563,5574
follow|5575,5581
up|5582,5584
with|5585,5589
<EOL>|5590,5591
her|5591,5594
primary|5595,5602
care|5603,5607
provider|5608,5616
to|5617,5619
address|5620,5627
management|5628,5638
of|5639,5641
her|5642,5645
chronic|5646,5653
<EOL>|5654,5655
pain|5655,5659
.|5659,5660
<EOL>|5661,5662
.|5662,5663
<EOL>|5663,5664
#|5664,5665
Diet|5665,5669
:|5669,5670
<EOL>|5670,5671
Low|5671,5674
sodium|5675,5681
(|5682,5683
2g|5683,5685
/|5685,5686
day|5686,5689
)|5689,5690
,|5690,5691
fluid|5692,5697
restriction|5698,5709
(|5710,5711
1500mL|5711,5717
/|5717,5718
day|5718,5721
)|5721,5722
<EOL>|5722,5723
.|5723,5724
<EOL>|5724,5725
#|5725,5726
Code|5726,5730
:|5730,5731
Full|5732,5736
<EOL>|5736,5737
<EOL>|5737,5738
<EOL>|5739,5740
Medications|5740,5751
on|5752,5754
Admission|5755,5764
:|5764,5765
<EOL>|5765,5766
-|5766,5767
AMITRIPTYLINE|5768,5781
-|5782,5783
10|5784,5786
mg|5787,5789
PO|5790,5792
HS|5793,5795
<EOL>|5797,5798
-|5798,5799
OXYCODONE|5800,5809
-|5810,5811
5|5812,5813
mg|5814,5816
PO|5817,5819
Q8H|5820,5823
PRN|5824,5827
pain|5828,5832
<EOL>|5834,5835
-|5835,5836
Thiamine|5837,5845
100mg|5846,5851
PO|5852,5854
daily|5855,5860
<EOL>|5862,5863
-|5863,5864
Folic|5865,5870
acid|5871,5875
1mg|5876,5879
PO|5880,5882
daily|5883,5888
<EOL>|5890,5891
-|5891,5892
MVI|5893,5896
PO|5897,5899
daily|5900,5905
<EOL>|5907,5908
<EOL>|5909,5910
Discharge|5910,5919
Medications|5920,5931
:|5931,5932
<EOL>|5932,5933
1.|5933,5935
Thiamine|5936,5944
HCl|5945,5948
100|5949,5952
mg|5953,5955
Tablet|5956,5962
Sig|5963,5966
:|5966,5967
One|5968,5971
(|5972,5973
1|5973,5974
)|5974,5975
Tablet|5976,5982
PO|5983,5985
DAILY|5986,5991
<EOL>|5992,5993
(|5993,5994
Daily|5994,5999
)|5999,6000
.|6000,6001
<EOL>|6001,6002
2.|6002,6004
Folic|6005,6010
Acid|6011,6015
1|6016,6017
mg|6018,6020
Tablet|6021,6027
Sig|6028,6031
:|6031,6032
One|6033,6036
(|6037,6038
1|6038,6039
)|6039,6040
Tablet|6041,6047
PO|6048,6050
DAILY|6051,6056
(|6057,6058
Daily|6058,6063
)|6063,6064
.|6064,6065
<EOL>|6067,6068
<EOL>|6068,6069
3.|6069,6071
Amitriptyline|6072,6085
10|6086,6088
mg|6089,6091
Tablet|6092,6098
Sig|6099,6102
:|6102,6103
One|6104,6107
(|6108,6109
1|6109,6110
)|6110,6111
Tablet|6112,6118
PO|6119,6121
HS|6122,6124
(|6125,6126
at|6126,6128
<EOL>|6129,6130
bedtime|6130,6137
)|6137,6138
.|6138,6139
<EOL>|6141,6142
4.|6142,6144
Multivitamin|6145,6157
Tablet|6162,6168
Sig|6169,6172
:|6172,6173
One|6174,6177
(|6178,6179
1|6179,6180
)|6180,6181
Tablet|6182,6188
PO|6189,6191
DAILY|6192,6197
(|6198,6199
Daily|6199,6204
)|6204,6205
.|6205,6206
<EOL>|6207,6208
<EOL>|6209,6210
5.|6210,6212
Lactulose|6213,6222
10|6223,6225
gram|6226,6230
/|6230,6231
15|6231,6233
mL|6234,6236
Syrup|6237,6242
Sig|6243,6246
:|6246,6247
Thirty|6248,6254
(|6255,6256
30|6256,6258
)|6258,6259
ML|6260,6262
PO|6263,6265
DAILY|6266,6271
<EOL>|6272,6273
(|6273,6274
Daily|6274,6279
)|6279,6280
.|6280,6281
<EOL>|6283,6284
6.|6284,6286
Oxycodone|6287,6296
5|6297,6298
mg|6299,6301
Tablet|6302,6308
Sig|6309,6312
:|6312,6313
One|6314,6317
(|6318,6319
1|6319,6320
)|6320,6321
Tablet|6322,6328
PO|6329,6331
every|6332,6337
eight|6338,6343
(|6344,6345
8|6345,6346
)|6346,6347
<EOL>|6348,6349
hours|6349,6354
as|6355,6357
needed|6358,6364
for|6365,6368
pain|6369,6373
.|6373,6374
<EOL>|6376,6377
<EOL>|6377,6378
<EOL>|6379,6380
Discharge|6380,6389
Disposition|6390,6401
:|6401,6402
<EOL>|6402,6403
Home|6403,6407
<EOL>|6407,6408
<EOL>|6409,6410
Discharge|6410,6419
Diagnosis|6420,6429
:|6429,6430
<EOL>|6430,6431
Primary|6431,6438
:|6438,6439
<EOL>|6439,6440
Ascites|6440,6447
<EOL>|6447,6448
Portal|6448,6454
hypertension|6455,6467
<EOL>|6467,6468
Alcoholic|6468,6477
hepatitis|6478,6487
<EOL>|6487,6488
.|6488,6489
<EOL>|6489,6490
Secondary|6490,6499
:|6499,6500
<EOL>|6500,6501
Chronic|6501,6508
back|6509,6513
pain|6514,6518
<EOL>|6518,6519
<EOL>|6519,6520
<EOL>|6521,6522
Discharge|6522,6531
Condition|6532,6541
:|6541,6542
<EOL>|6542,6543
Alert|6543,6548
and|6549,6552
Oriented|6553,6561
.|6561,6562
Ambulating|6564,6574
without|6575,6582
help|6583,6587
.|6587,6588
Hemodynamically|6590,6605
<EOL>|6606,6607
stable|6607,6613
,|6613,6614
afebrile|6615,6623
,|6623,6624
tachycardic|6625,6636
.|6636,6637
<EOL>|6639,6640
<EOL>|6640,6641
<EOL>|6642,6643
Discharge|6643,6652
Instructions|6653,6665
:|6665,6666
<EOL>|6666,6667
You|6667,6670
were|6671,6675
seen|6676,6680
in|6681,6683
the|6684,6687
_|6688,6689
_|6689,6690
_|6690,6691
Associates|6692,6702
with|6703,6707
<EOL>|6708,6709
complaints|6709,6719
of|6720,6722
increasing|6723,6733
abdominal|6734,6743
distention|6744,6754
and|6755,6758
pain|6759,6763
.|6763,6764
In|6765,6767
the|6768,6771
<EOL>|6772,6773
clinic|6773,6779
,|6779,6780
you|6781,6784
also|6785,6789
had|6790,6793
a|6794,6795
mild|6796,6800
fever|6801,6806
,|6806,6807
fast|6808,6812
heart|6813,6818
rate|6819,6823
,|6823,6824
and|6825,6828
<EOL>|6829,6830
increased|6830,6839
white|6840,6845
blood|6846,6851
count|6852,6857
.|6857,6858
You|6860,6863
were|6864,6868
sent|6869,6873
to|6874,6876
the|6877,6880
emergency|6881,6890
<EOL>|6891,6892
department|6892,6902
and|6903,6906
admitted|6907,6915
to|6916,6918
the|6919,6922
hospital|6923,6931
for|6932,6935
further|6936,6943
workup|6944,6950
.|6950,6951
<EOL>|6953,6954
During|6954,6960
the|6961,6964
hospitalization|6965,6980
your|6981,6985
ascitic|6986,6993
fluid|6994,6999
was|7000,7003
tapped|7004,7010
and|7011,7014
<EOL>|7015,7016
analyzed|7016,7024
.|7024,7025
The|7027,7030
result|7031,7037
showed|7038,7044
that|7045,7049
you|7050,7053
did|7054,7057
not|7058,7061
have|7062,7066
an|7067,7069
infection|7070,7079
<EOL>|7080,7081
of|7081,7083
the|7084,7087
ascitic|7088,7095
fluid|7096,7101
.|7101,7102
Subsequently|7104,7116
,|7116,7117
fluid|7118,7123
was|7124,7127
removed|7128,7135
from|7136,7140
your|7141,7145
<EOL>|7146,7147
abdomen|7147,7154
via|7155,7158
paracentesis|7159,7171
.|7171,7172
We|7173,7175
also|7176,7180
started|7181,7188
a|7189,7190
24|7191,7193
-|7193,7194
hr|7194,7196
urine|7197,7202
<EOL>|7203,7204
collection|7204,7214
for|7215,7218
copper|7219,7225
to|7226,7228
work|7229,7233
up|7234,7236
for|7237,7240
other|7241,7246
potential|7247,7256
causes|7257,7263
of|7264,7266
<EOL>|7267,7268
your|7268,7272
liver|7273,7278
disease|7279,7286
.|7286,7287
The|7289,7292
liver|7293,7298
clinic|7299,7305
will|7306,7310
follow|7311,7317
up|7318,7320
with|7321,7325
you|7326,7329
<EOL>|7330,7331
regarding|7331,7340
the|7341,7344
results|7345,7352
of|7353,7355
these|7356,7361
tests|7362,7367
.|7367,7368
<EOL>|7370,7371
.|7371,7372
<EOL>|7372,7373
Your|7373,7377
back|7378,7382
pain|7383,7387
persisted|7388,7397
during|7398,7404
your|7405,7409
hospitalization|7410,7425
.|7425,7426
You|7428,7431
<EOL>|7432,7433
underwent|7433,7442
x-rays|7443,7449
which|7450,7455
showed|7456,7462
no|7463,7465
evidence|7466,7474
of|7475,7477
fracture|7478,7486
or|7487,7489
bone|7490,7494
<EOL>|7495,7496
infection|7496,7505
.|7505,7506
Please|7508,7514
continue|7515,7523
your|7524,7528
home|7529,7533
pain|7534,7538
regimen|7539,7546
and|7547,7550
readdress|7551,7560
<EOL>|7561,7562
with|7562,7566
your|7567,7571
primary|7572,7579
care|7580,7584
provider|7585,7593
.|7593,7594
<EOL>|7594,7595
.|7595,7596
<EOL>|7596,7597
No|7597,7599
changes|7600,7607
were|7608,7612
made|7613,7617
to|7618,7620
your|7621,7625
home|7626,7630
medications|7631,7642
.|7642,7643
You|7645,7648
should|7649,7655
<EOL>|7656,7657
continue|7657,7665
to|7666,7668
use|7669,7672
lactulose|7673,7682
for|7683,7686
constipation|7687,7699
while|7700,7705
using|7706,7711
pain|7712,7716
<EOL>|7717,7718
medications|7718,7729
.|7729,7730
<EOL>|7732,7733
.|7733,7734
<EOL>|7734,7735
Please|7735,7741
stop|7742,7746
using|7747,7752
all|7753,7756
herbal|7757,7763
or|7764,7766
tonic|7767,7772
remedies|7773,7781
until|7782,7787
your|7788,7792
liver|7793,7798
<EOL>|7799,7800
function|7800,7808
has|7809,7812
recovered|7813,7822
.|7822,7823
Some|7824,7828
of|7829,7831
these|7832,7837
therapies|7838,7847
may|7848,7851
interact|7852,7860
<EOL>|7861,7862
with|7862,7866
your|7867,7871
current|7872,7879
medications|7880,7891
or|7892,7894
make|7895,7899
it|7900,7902
difficult|7903,7912
to|7913,7915
interpret|7916,7925
<EOL>|7926,7927
your|7927,7931
laboratory|7932,7942
results|7943,7950
.|7950,7951
<EOL>|7951,7952
<EOL>|7953,7954
Followup|7954,7962
Instructions|7963,7975
:|7975,7976
<EOL>|7976,7977
_|7977,7978
_|7978,7979
_|7979,7980
<EOL>|7980,7981

