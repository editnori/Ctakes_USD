 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
PLASTIC|156,163
<EOL>|163,164
<EOL>|165,166
Penicillins|178,189
/|190,191
Paxil|192,197
/|198,199
Wellbutrin|200,210
<EOL>|210,211
<EOL>|212,213
Attending|213,222
:|222,223
_|224,225
_|225,226
_|226,227
.|227,228
<EOL>|228,229
<EOL>|230,231
exposed|248,255
craniotomy|256,266
hardware|267,275
<EOL>|276,277
<EOL>|278,279
Major|279,284
Surgical|285,293
or|294,296
Invasive|297,305
Procedure|306,315
:|315,316
<EOL>|316,317
Right|317,322
scalp|323,328
flap|329,333
with|334,338
split|339,344
thickness|345,354
skin|355,359
graft|360,365
and|366,369
wound|370,375
VAC|376,379
<EOL>|380,381
placement|381,390
<EOL>|390,391
<EOL>|391,392
<EOL>|393,394
_|422,423
_|423,424
_|424,425
year|426,430
old|431,434
female|435,441
with|442,446
multiple|447,455
prior|456,461
surgeries|462,471
for|472,475
right|476,481
<EOL>|482,483
parietal|483,491
anaplastic|492,502
astrocytoma|503,514
diagnosed|515,524
in|525,527
_|528,529
_|529,530
_|530,531
.|531,532
She|533,536
has|537,540
also|541,545
<EOL>|546,547
undergone|547,556
chemo|557,562
and|563,566
radiation|567,576
.|576,577
She|578,581
presented|582,591
to|592,594
_|595,596
_|596,597
_|597,598
in|599,601
<EOL>|602,603
_|603,604
_|604,605
_|605,606
with|607,611
_|612,613
_|613,614
_|614,615
month|616,621
history|622,629
of|630,632
pruritus|633,641
on|642,644
the|645,648
top|649,652
of|653,655
her|656,659
head|660,664
.|664,665
<EOL>|666,667
She|667,670
reports|671,678
that|679,683
she|684,687
had|688,691
her|692,695
husband|696,703
look|704,708
at|709,711
the|712,715
top|716,719
of|720,722
her|723,726
head|727,731
<EOL>|732,733
and|733,736
her|737,740
found|741,746
her|747,750
metal|751,756
hardware|757,765
from|766,770
her|771,774
prior|775,780
surgery|781,788
was|789,792
<EOL>|793,794
present|794,801
.|801,802
On|803,805
_|806,807
_|807,808
_|808,809
Dr.|810,813
_|814,815
_|815,816
_|816,817
metal|818,823
hardware|824,832
(|833,834
removal|834,841
of|842,844
<EOL>|845,846
harware|846,853
but|854,857
not|858,861
the|862,865
bone|866,870
flap|871,875
)|875,876
.|876,877
She|878,881
presented|882,891
today|892,897
for|898,901
a|902,903
<EOL>|904,905
rotational|905,915
flap|916,920
and|921,924
skin|925,929
graft|930,935
for|936,939
proper|940,946
coverage|947,955
of|956,958
wound|959,964
.|964,965
<EOL>|966,967
<EOL>|968,969
right|991,996
parietal|997,1005
anaplastic|1006,1016
astrocytoma|1017,1028
,|1028,1029
Craniotomy|1029,1039
_|1040,1041
_|1041,1042
_|1042,1043
by|1044,1046
<EOL>|1048,1049
Dr.|1049,1052
_|1053,1054
_|1054,1055
_|1055,1056
in|1057,1059
_|1060,1061
_|1061,1062
_|1062,1063
irradiation|1064,1075
to|1076,1078
6,120|1079,1084
<EOL>|1085,1086
<EOL>|1087,1088
cGy|1088,1091
_|1092,1093
_|1093,1094
_|1094,1095
in|1096,1098
_|1099,1100
_|1100,1101
_|1101,1102
,|1102,1103
3|1103,1104
cycles|1105,1111
of|1112,1114
Temodar|1115,1122
ended|1123,1128
_|1129,1130
_|1130,1131
_|1131,1132
<EOL>|1134,1135
craniotomy|1135,1145
on|1146,1148
_|1149,1150
_|1150,1151
_|1151,1152
by|1153,1155
Dr.|1156,1159
_|1160,1161
_|1161,1162
_|1162,1163
at|1164,1166
_|1167,1168
_|1168,1169
_|1169,1170
_|1171,1172
_|1172,1173
_|1173,1174
-|1175,1176
<EOL>|1178,1179
_|1179,1180
_|1180,1181
_|1181,1182
wound|1183,1188
revision|1189,1197
and|1198,1201
removal|1202,1209
of|1210,1212
the|1213,1216
exposed|1217,1224
craniotx|1225,1233
<EOL>|1234,1235
hardware|1235,1243
,|1243,1244
Accutane|1245,1253
for|1254,1257
2|1258,1259
weeks|1260,1265
only|1266,1270
_|1271,1272
_|1272,1273
_|1273,1274
disease|1275,1282
since|1283,1288
<EOL>|1289,1290
_|1290,1291
_|1291,1292
_|1292,1293
,|1293,1294
<EOL>|1296,1297
tubal|1297,1302
ligation|1303,1311
,|1311,1312
tonsillectomy|1312,1325
,|1325,1326
bronchitis|1327,1337
,|1337,1338
depression|1339,1349
.|1349,1350
<EOL>|1352,1353
seizures|1353,1361
<EOL>|1363,1364
<EOL>|1364,1365
<EOL>|1366,1367
:|1381,1382
<EOL>|1382,1383
_|1383,1384
_|1384,1385
_|1385,1386
<EOL>|1386,1387
:|1401,1402
<EOL>|1402,1403
NC|1403,1405
<EOL>|1405,1406
<EOL>|1407,1408
Afebrile|1423,1431
.|1431,1432
vital|1433,1438
signs|1439,1444
stable|1445,1451
.|1451,1452
Right|1453,1458
scalp|1459,1464
incision|1465,1473
clean|1474,1479
,|1479,1480
dry|1481,1484
<EOL>|1485,1486
and|1486,1489
intact|1490,1496
with|1497,1501
xeroform|1502,1510
dressing|1511,1519
in|1520,1522
place|1523,1528
.|1528,1529
Right|1530,1535
STSG|1536,1540
site|1541,1545
with|1546,1550
<EOL>|1551,1552
bolstered|1552,1561
xeroform|1562,1570
dressing|1571,1579
in|1580,1582
place|1583,1588
.|1588,1589
No|1590,1592
drainage|1593,1601
or|1602,1604
bleeding|1605,1613
.|1613,1614
<EOL>|1614,1615
<EOL>|1616,1617
Pertinent|1617,1626
Results|1627,1634
:|1634,1635
<EOL>|1635,1636
None|1636,1640
this|1641,1645
admission|1646,1655
.|1655,1656
<EOL>|1656,1657
<EOL>|1658,1659
The|1682,1685
patient|1686,1693
was|1694,1697
admitted|1698,1706
to|1707,1709
the|1710,1713
plastic|1714,1721
surgery|1722,1729
service|1730,1737
on|1738,1740
<EOL>|1741,1742
_|1742,1743
_|1743,1744
_|1744,1745
and|1746,1749
had|1750,1753
a|1754,1755
flap|1756,1760
and|1761,1764
skin|1765,1769
graft|1770,1775
to|1776,1778
your|1779,1783
scalp|1784,1789
defect|1790,1796
.|1796,1797
<EOL>|1799,1800
The|1800,1803
patient|1804,1811
tolerated|1812,1821
the|1822,1825
procedure|1826,1835
well|1836,1840
.|1840,1841
<EOL>|1842,1843
.|1843,1844
<EOL>|1844,1845
Neuro|1845,1850
:|1850,1851
Post-operatively|1852,1868
,|1868,1869
the|1870,1873
patient|1874,1881
received|1882,1890
vicodin|1891,1898
with|1899,1903
good|1904,1908
<EOL>|1909,1910
pain|1910,1914
relief|1915,1921
noted|1922,1927
.|1927,1928
<EOL>|1928,1929
.|1929,1930
<EOL>|1930,1931
CV|1931,1933
:|1933,1934
The|1935,1938
patient|1939,1946
was|1947,1950
stable|1951,1957
from|1958,1962
a|1963,1964
cardiovascular|1965,1979
standpoint|1980,1990
;|1990,1991
<EOL>|1992,1993
vital|1993,1998
signs|1999,2004
were|2005,2009
routinely|2010,2019
monitored|2020,2029
.|2029,2030
<EOL>|2030,2031
.|2031,2032
<EOL>|2032,2033
Pulmonary|2033,2042
:|2042,2043
The|2044,2047
patient|2048,2055
was|2056,2059
stable|2060,2066
from|2067,2071
a|2072,2073
pulmonary|2074,2083
standpoint|2084,2094
;|2094,2095
<EOL>|2096,2097
vital|2097,2102
signs|2103,2108
were|2109,2113
routinely|2114,2123
monitored|2124,2133
.|2133,2134
<EOL>|2134,2135
.|2135,2136
<EOL>|2136,2137
GI|2137,2139
/|2139,2140
GU|2140,2142
:|2142,2143
Post-operatively|2144,2160
,|2160,2161
the|2162,2165
patient|2166,2173
was|2174,2177
given|2178,2183
IV|2184,2186
fluids|2187,2193
until|2194,2199
<EOL>|2200,2201
tolerating|2201,2211
oral|2212,2216
intake|2217,2223
.|2223,2224
Her|2225,2228
diet|2229,2233
was|2234,2237
advanced|2238,2246
when|2247,2251
appropriate|2252,2263
,|2263,2264
<EOL>|2265,2266
which|2266,2271
was|2272,2275
tolerated|2276,2285
well|2286,2290
.|2290,2291
She|2292,2295
was|2296,2299
also|2300,2304
started|2305,2312
on|2313,2315
a|2316,2317
bowel|2318,2323
<EOL>|2324,2325
regimen|2325,2332
to|2333,2335
encourage|2336,2345
bowel|2346,2351
movement|2352,2360
.|2360,2361
Intake|2362,2368
and|2369,2372
output|2373,2379
were|2380,2384
<EOL>|2385,2386
closely|2386,2393
monitored|2394,2403
.|2403,2404
<EOL>|2405,2406
.|2406,2407
<EOL>|2407,2408
ID|2408,2410
:|2410,2411
Post-operatively|2412,2428
,|2428,2429
the|2430,2433
patient|2434,2441
was|2442,2445
started|2446,2453
on|2454,2456
IV|2457,2459
cefazolin|2460,2469
,|2469,2470
<EOL>|2471,2472
then|2472,2476
switched|2477,2485
to|2486,2488
PO|2489,2491
cefadroxil|2492,2502
for|2503,2506
discharge|2507,2516
home|2517,2521
.|2521,2522
The|2523,2526
patient|2527,2534
's|2534,2536
<EOL>|2537,2538
temperature|2538,2549
was|2550,2553
closely|2554,2561
watched|2562,2569
for|2570,2573
signs|2574,2579
of|2580,2582
infection|2583,2592
.|2592,2593
<EOL>|2594,2595
.|2595,2596
<EOL>|2596,2597
Prophylaxis|2597,2608
:|2608,2609
The|2610,2613
patient|2614,2621
received|2622,2630
subcutaneous|2631,2643
heparin|2644,2651
during|2652,2658
<EOL>|2659,2660
this|2660,2664
stay|2665,2669
,|2669,2670
and|2671,2674
was|2675,2678
encouraged|2679,2689
to|2690,2692
get|2693,2696
up|2697,2699
and|2700,2703
ambulate|2704,2712
as|2713,2715
early|2716,2721
as|2722,2724
<EOL>|2725,2726
possible|2726,2734
.|2734,2735
<EOL>|2736,2737
.|2737,2738
<EOL>|2738,2739
At|2739,2741
the|2742,2745
time|2746,2750
of|2751,2753
discharge|2754,2763
on|2764,2766
POD|2767,2770
#|2770,2771
1|2771,2772
,|2772,2773
the|2774,2777
patient|2778,2785
was|2786,2789
doing|2790,2795
well|2796,2800
,|2800,2801
<EOL>|2802,2803
afebrile|2803,2811
with|2812,2816
stable|2817,2823
vital|2824,2829
signs|2830,2835
,|2835,2836
tolerating|2837,2847
a|2848,2849
regular|2850,2857
diet|2858,2862
,|2862,2863
<EOL>|2864,2865
ambulating|2865,2875
,|2875,2876
voiding|2877,2884
without|2885,2892
assistance|2893,2903
,|2903,2904
and|2905,2908
pain|2909,2913
was|2914,2917
well|2918,2922
<EOL>|2923,2924
controlled|2924,2934
.|2934,2935
Her|2936,2939
scalp|2940,2945
graft|2946,2951
site|2952,2956
was|2957,2960
clean|2961,2966
and|2967,2970
pink|2971,2975
and|2976,2979
she|2980,2983
had|2984,2987
<EOL>|2988,2989
xeroform|2989,2997
dressing|2998,3006
intact|3007,3013
.|3013,3014
Her|3016,3019
right|3020,3025
thing|3026,3031
graft|3032,3037
donor|3038,3043
site|3044,3048
had|3049,3052
<EOL>|3053,3054
original|3054,3062
xeroform|3063,3071
dressing|3072,3080
in|3081,3083
place|3084,3089
to|3090,3092
left|3093,3097
open|3098,3102
to|3103,3105
air|3106,3109
to|3110,3112
dry|3113,3116
<EOL>|3117,3118
out|3118,3121
.|3121,3122
<EOL>|3122,3123
<EOL>|3123,3124
<EOL>|3125,3126
Medications|3126,3137
on|3138,3140
Admission|3141,3150
:|3150,3151
<EOL>|3151,3152
_|3152,3153
_|3153,3154
_|3154,3155
:|3155,3156
azathioprine|3157,3169
,|3169,3170
Pentasa|3171,3178
,|3178,3179
topiramate|3180,3190
,|3190,3191
alprazolam|3192,3202
,|3202,3203
omeprazole|3204,3214
,|3214,3215
<EOL>|3216,3217
zolpidem|3217,3225
,|3225,3226
venlafaxine|3227,3238
hcl|3239,3242
er|3243,3245
30|3246,3248
,|3248,3249
popylthiouracil|3250,3265
,|3265,3266
promethazine|3267,3279
,|3279,3280
<EOL>|3281,3282
keflex|3282,3288
<EOL>|3289,3290
<EOL>|3291,3292
Discharge|3292,3301
Medications|3302,3313
:|3313,3314
<EOL>|3314,3315
1.|3315,3317
azathioprine|3318,3330
75|3331,3333
mg|3334,3336
Tablet|3337,3343
Sig|3344,3347
:|3347,3348
One|3349,3352
(|3353,3354
1|3354,3355
)|3355,3356
Tablet|3357,3363
PO|3364,3366
DAILY|3367,3372
<EOL>|3373,3374
(|3374,3375
Daily|3375,3380
)|3380,3381
.|3381,3382
<EOL>|3384,3385
2.|3385,3387
dicyclomine|3388,3399
10|3400,3402
mg|3403,3405
Capsule|3406,3413
Sig|3414,3417
:|3417,3418
One|3419,3422
(|3423,3424
1|3424,3425
)|3425,3426
Capsule|3427,3434
PO|3435,3437
Q8H|3438,3441
(|3442,3443
every|3443,3448
<EOL>|3449,3450
8|3450,3451
hours|3452,3457
)|3457,3458
as|3459,3461
needed|3462,3468
for|3469,3472
abdominal|3473,3482
pain|3483,3487
.|3487,3488
<EOL>|3490,3491
3.|3491,3493
fluticasone|3494,3505
-|3505,3506
salmeterol|3506,3516
500|3517,3520
-|3520,3521
50|3521,3523
mcg|3524,3527
/|3527,3528
dose|3528,3532
Disk|3533,3537
with|3538,3542
Device|3543,3549
Sig|3550,3553
:|3553,3554
<EOL>|3555,3556
One|3556,3559
(|3560,3561
1|3561,3562
)|3562,3563
Disk|3564,3568
with|3569,3573
Device|3574,3580
Inhalation|3581,3591
BID|3592,3595
(|3596,3597
2|3597,3598
times|3599,3604
a|3605,3606
day|3607,3610
)|3610,3611
.|3611,3612
<EOL>|3614,3615
4.|3615,3617
mesalamine|3618,3628
250|3629,3632
mg|3633,3635
Capsule|3636,3643
,|3643,3644
Extended|3645,3653
Release|3654,3661
Sig|3662,3665
:|3665,3666
Two|3667,3670
(|3671,3672
2|3672,3673
)|3673,3674
<EOL>|3675,3676
Capsule|3676,3683
,|3683,3684
Extended|3685,3693
Release|3694,3701
PO|3702,3704
QID|3705,3708
(|3709,3710
4|3710,3711
times|3712,3717
a|3718,3719
day|3720,3723
)|3723,3724
.|3724,3725
<EOL>|3727,3728
5.|3728,3730
omeprazole|3731,3741
20|3742,3744
mg|3745,3747
Capsule|3748,3755
,|3755,3756
Delayed|3757,3764
Release|3765,3772
(|3772,3773
E.C|3773,3776
.|3776,3777
)|3777,3778
Sig|3779,3782
:|3782,3783
One|3784,3787
(|3788,3789
1|3789,3790
)|3790,3791
<EOL>|3792,3793
Capsule|3793,3800
,|3800,3801
Delayed|3802,3809
Release|3810,3817
(|3817,3818
E.C|3818,3821
.|3821,3822
)|3822,3823
PO|3824,3826
DAILY|3827,3832
(|3833,3834
Daily|3834,3839
)|3839,3840
.|3840,3841
<EOL>|3843,3844
6.|3844,3846
topiramate|3847,3857
100|3858,3861
mg|3862,3864
Tablet|3865,3871
Sig|3872,3875
:|3875,3876
Two|3877,3880
(|3881,3882
2|3882,3883
)|3883,3884
Tablet|3885,3891
PO|3892,3894
BID|3895,3898
(|3899,3900
2|3900,3901
times|3902,3907
<EOL>|3908,3909
a|3909,3910
day|3911,3914
)|3914,3915
.|3915,3916
<EOL>|3918,3919
7.|3919,3921
venlafaxine|3922,3933
75|3934,3936
mg|3937,3939
Capsule|3940,3947
,|3947,3948
Ext|3949,3952
Release|3953,3960
24|3961,3963
hr|3964,3966
Sig|3967,3970
:|3970,3971
Three|3972,3977
(|3978,3979
3|3979,3980
)|3980,3981
<EOL>|3982,3983
Capsule|3983,3990
,|3990,3991
Ext|3992,3995
Release|3996,4003
24|4004,4006
hr|4007,4009
PO|4010,4012
DAILY|4013,4018
(|4019,4020
Daily|4020,4025
)|4025,4026
.|4026,4027
<EOL>|4029,4030
8.|4030,4032
propylthiouracil|4033,4049
50|4050,4052
mg|4053,4055
Tablet|4056,4062
Sig|4063,4066
:|4066,4067
Two|4068,4071
(|4072,4073
2|4073,4074
)|4074,4075
Tablet|4076,4082
PO|4083,4085
Q8H|4086,4089
<EOL>|4090,4091
(|4091,4092
every|4092,4097
8|4098,4099
hours|4100,4105
)|4105,4106
.|4106,4107
<EOL>|4109,4110
9.|4110,4112
bacitracin|4113,4123
zinc|4124,4128
500|4129,4132
unit|4133,4137
/|4137,4138
g|4138,4139
Ointment|4140,4148
Sig|4149,4152
:|4152,4153
One|4154,4157
(|4158,4159
1|4159,4160
)|4160,4161
Appl|4162,4166
Topical|4167,4174
<EOL>|4175,4176
BID|4176,4179
(|4180,4181
2|4181,4182
times|4183,4188
a|4189,4190
day|4191,4194
)|4194,4195
.|4195,4196
<EOL>|4196,4197
Disp|4197,4201
:|4201,4202
*|4202,4203
1|4203,4204
tube|4205,4209
*|4209,4210
Refills|4211,4218
:|4218,4219
*|4219,4220
2|4220,4221
*|4221,4222
<EOL>|4222,4223
10.|4223,4226
cefadroxil|4227,4237
500|4238,4241
mg|4242,4244
Capsule|4245,4252
Sig|4253,4256
:|4256,4257
One|4258,4261
(|4262,4263
1|4263,4264
)|4264,4265
Capsule|4266,4273
PO|4274,4276
twice|4277,4282
a|4283,4284
<EOL>|4285,4286
day|4286,4289
for|4290,4293
7|4294,4295
days|4296,4300
.|4300,4301
<EOL>|4301,4302
Disp|4302,4306
:|4306,4307
*|4307,4308
14|4308,4310
Capsule|4311,4318
(|4318,4319
s|4319,4320
)|4320,4321
*|4321,4322
Refills|4323,4330
:|4330,4331
*|4331,4332
0|4332,4333
*|4333,4334
<EOL>|4334,4335
11.|4335,4338
hydrocodone|4339,4350
-|4350,4351
acetaminophen|4351,4364
_|4365,4366
_|4366,4367
_|4367,4368
mg|4369,4371
Tablet|4372,4378
Sig|4379,4382
:|4382,4383
_|4384,4385
_|4385,4386
_|4386,4387
Tablets|4388,4395
<EOL>|4396,4397
PO|4397,4399
every|4400,4405
six|4406,4409
(|4410,4411
6|4411,4412
)|4412,4413
hours|4414,4419
as|4420,4422
needed|4423,4429
for|4430,4433
pain|4434,4438
:|4438,4439
Max|4440,4443
8|4444,4445
/|4445,4446
day|4446,4449
.|4449,4450
.|4451,4452
<EOL>|4452,4453
Disp|4453,4457
:|4457,4458
*|4458,4459
40|4459,4461
Tablet|4462,4468
(|4468,4469
s|4469,4470
)|4470,4471
*|4471,4472
Refills|4473,4480
:|4480,4481
*|4481,4482
0|4482,4483
*|4483,4484
<EOL>|4484,4485
12.|4485,4488
alprazolam|4489,4499
0.25|4500,4504
mg|4505,4507
Tablet|4508,4514
Sig|4515,4518
:|4518,4519
Two|4520,4523
(|4524,4525
2|4525,4526
)|4526,4527
Tablet|4528,4534
PO|4535,4537
TID|4538,4541
(|4542,4543
3|4543,4544
<EOL>|4545,4546
times|4546,4551
a|4552,4553
day|4554,4557
)|4557,4558
as|4559,4561
needed|4562,4568
for|4569,4572
anxiety|4573,4580
.|4580,4581
<EOL>|4583,4584
<EOL>|4584,4585
<EOL>|4586,4587
Discharge|4587,4596
Disposition|4597,4608
:|4608,4609
<EOL>|4609,4610
Home|4610,4614
With|4615,4619
Service|4620,4627
<EOL>|4627,4628
<EOL>|4629,4630
Facility|4630,4638
:|4638,4639
<EOL>|4639,4640
_|4640,4641
_|4641,4642
_|4642,4643
<EOL>|4644,4645
<EOL>|4646,4647
Discharge|4647,4656
Diagnosis|4657,4666
:|4666,4667
<EOL>|4667,4668
exposed|4668,4675
craniotomy|4676,4686
wound|4687,4692
Status|4693,4699
post|4700,4704
hardware|4705,4713
removal|4714,4721
,|4721,4722
split|4723,4728
<EOL>|4729,4730
thickness|4730,4739
skin|4740,4744
graft|4745,4750
application|4751,4762
to|4763,4765
scalp|4766,4771
,|4771,4772
donor|4773,4778
site|4779,4783
from|4784,4788
leg|4789,4792
<EOL>|4792,4793
<EOL>|4793,4794
<EOL>|4795,4796
Mental|4817,4823
Status|4824,4830
:|4830,4831
Clear|4832,4837
and|4838,4841
coherent|4842,4850
.|4850,4851
<EOL>|4851,4852
Level|4852,4857
of|4858,4860
Consciousness|4861,4874
:|4874,4875
Alert|4876,4881
and|4882,4885
interactive|4886,4897
.|4897,4898
<EOL>|4898,4899
Activity|4899,4907
Status|4908,4914
:|4914,4915
Ambulatory|4916,4926
-|4927,4928
Independent|4929,4940
.|4940,4941
<EOL>|4941,4942
<EOL>|4942,4943
<EOL>|4944,4945
-|4969,4970
The|4970,4973
hemovac|4974,4981
drain|4982,4987
should|4988,4994
always|4995,5001
be|5002,5004
collapsed|5005,5014
so|5015,5017
as|5018,5020
to|5021,5023
apply|5024,5029
<EOL>|5030,5031
constant|5031,5039
suction|5040,5047
to|5048,5050
the|5051,5054
wound|5055,5060
.|5060,5061
Does|5062,5066
not|5067,5070
need|5071,5075
to|5076,5078
be|5079,5081
emptied|5082,5089
<EOL>|5090,5091
unless|5091,5097
not|5098,5101
collapsed|5102,5111
and|5112,5115
does|5116,5120
not|5121,5124
have|5125,5129
suction|5130,5137
.|5137,5138
<EOL>|5138,5139
-|5139,5140
Your|5140,5144
skin|5145,5149
graft|5150,5155
site|5156,5160
on|5161,5163
your|5164,5168
scalp|5169,5174
should|5175,5181
be|5182,5184
covered|5185,5192
with|5193,5197
a|5198,5199
<EOL>|5200,5201
Xeroform|5201,5209
dressing|5210,5218
and|5219,5222
you|5223,5226
should|5227,5233
apply|5234,5239
bacitracin|5240,5250
ointment|5251,5259
with|5260,5264
<EOL>|5265,5266
Qtips|5266,5271
UNDER|5272,5277
the|5278,5281
xeroform|5282,5290
dressing|5291,5299
twice|5300,5305
a|5306,5307
day|5308,5311
.|5311,5312
WARNING|5314,5321
:|5321,5322
do|5323,5325
NOT|5326,5329
<EOL>|5330,5331
change|5331,5337
the|5338,5341
xeroform|5342,5350
that|5351,5355
is|5356,5358
sewn|5359,5363
/|5363,5364
sutured|5364,5371
in|5372,5374
place|5375,5380
<EOL>|5381,5382
already|5382,5389
...|5389,5392
leave|5392,5397
that|5398,5402
in|5403,5405
place|5406,5411
.|5411,5412
<EOL>|5412,5413
-|5413,5414
Please|5414,5420
keep|5421,5425
your|5426,5430
skin|5431,5435
graft|5436,5441
site|5442,5446
free|5447,5451
of|5452,5454
any|5455,5458
pressure|5459,5467
or|5468,5470
<EOL>|5471,5472
extreme|5472,5479
temperatures|5480,5492
(|5493,5494
cover|5494,5499
with|5500,5504
loose|5505,5510
hat|5511,5514
that|5515,5519
does|5520,5524
not|5525,5528
sit|5529,5532
on|5533,5535
<EOL>|5536,5537
your|5537,5541
graft|5542,5547
site|5548,5552
)|5552,5553
.|5553,5554
<EOL>|5554,5555
-|5555,5556
You|5556,5559
may|5560,5563
shower|5564,5570
48|5571,5573
hours|5574,5579
after|5580,5585
surgery|5586,5593
but|5594,5597
do|5598,5600
not|5601,5604
let|5605,5608
water|5609,5614
run|5615,5618
<EOL>|5619,5620
on|5620,5622
your|5623,5627
head|5628,5632
/|5632,5633
scalp|5633,5638
area|5639,5643
.|5643,5644
You|5646,5649
may|5650,5653
shower|5654,5660
from|5661,5665
the|5666,5669
neck|5670,5674
down|5675,5679
<EOL>|5680,5681
only|5681,5685
.|5685,5686
<EOL>|5686,5687
-|5687,5688
your|5688,5692
thigh|5693,5698
'|5699,5700
donor|5700,5705
site|5706,5710
'|5710,5711
should|5712,5718
be|5719,5721
left|5722,5726
'|5727,5728
open|5728,5732
to|5733,5735
air|5736,5739
'|5739,5740
and|5741,5744
left|5745,5749
<EOL>|5750,5751
to|5751,5753
dry|5754,5757
out|5758,5761
.|5761,5762
The|5764,5767
old|5768,5771
xeroform|5772,5780
dressing|5781,5789
will|5790,5794
peel|5795,5799
back|5800,5804
/|5804,5805
fall|5805,5809
off|5810,5813
<EOL>|5814,5815
on|5815,5817
its|5818,5821
own|5822,5825
.|5825,5826
When|5828,5832
you|5833,5836
shower|5837,5843
you|5844,5847
must|5848,5852
cover|5853,5858
your|5859,5863
thigh|5864,5869
'|5870,5871
donor|5871,5876
<EOL>|5877,5878
site|5878,5882
'|5882,5883
with|5884,5888
Plastic|5889,5896
wrap|5897,5901
to|5902,5904
keep|5905,5909
it|5910,5912
free|5913,5917
of|5918,5920
water|5921,5926
while|5927,5932
you|5933,5936
<EOL>|5937,5938
shower|5938,5944
.|5944,5945
You|5947,5950
may|5951,5954
remove|5955,5961
plastic|5962,5969
wrap|5970,5974
when|5975,5979
you|5980,5983
are|5984,5987
done|5988,5992
and|5993,5996
leave|5997,6002
<EOL>|6003,6004
the|6004,6007
donor|6008,6013
site|6014,6018
open|6019,6023
to|6024,6026
air|6027,6030
again|6031,6036
to|6037,6039
dry|6040,6043
out|6044,6047
.|6047,6048
<EOL>|6048,6049
.|6049,6050
<EOL>|6050,6051
Diet|6051,6055
/|6055,6056
Activity|6056,6064
:|6064,6065
<EOL>|6066,6067
1|6067,6068
.|6068,6069
You|6070,6073
may|6074,6077
resume|6078,6084
your|6085,6089
regular|6090,6097
diet|6098,6102
.|6102,6103
<EOL>|6104,6105
2.|6105,6107
DO|6108,6110
NOT|6111,6114
bend|6115,6119
over|6120,6124
,|6124,6125
avoid|6126,6131
heavy|6132,6137
lifting|6138,6145
and|6146,6149
do|6150,6152
not|6153,6156
engage|6157,6163
in|6164,6166
<EOL>|6167,6168
strenuous|6168,6177
activity|6178,6186
until|6187,6192
instructed|6193,6203
by|6204,6206
Dr.|6207,6210
_|6211,6212
_|6212,6213
_|6213,6214
.|6214,6215
<EOL>|6216,6217
.|6217,6218
<EOL>|6219,6220
1.|6234,6236
Resume|6237,6243
your|6244,6248
regular|6249,6256
medications|6257,6268
unless|6269,6275
instructed|6276,6286
otherwise|6287,6296
<EOL>|6297,6298
and|6298,6301
take|6302,6306
any|6307,6310
new|6311,6314
meds|6315,6319
as|6320,6322
ordered|6323,6330
.|6330,6331
<EOL>|6332,6333
2|6333,6334
.|6334,6335
You|6336,6339
may|6340,6343
take|6344,6348
your|6349,6353
prescribed|6354,6364
pain|6365,6369
medication|6370,6380
for|6381,6384
moderate|6385,6393
to|6394,6396
<EOL>|6397,6398
severe|6398,6404
pain|6405,6409
.|6409,6410
You|6411,6414
may|6415,6418
switch|6419,6425
to|6426,6428
Tylenol|6429,6436
or|6437,6439
Extra|6440,6445
Strength|6446,6454
Tylenol|6455,6462
<EOL>|6463,6464
<EOL>|6464,6465
for|6465,6468
mild|6469,6473
pain|6474,6478
as|6479,6481
directed|6482,6490
on|6491,6493
the|6494,6497
packaging|6498,6507
.|6507,6508
Please|6509,6515
note|6516,6520
that|6521,6525
<EOL>|6526,6527
Percocet|6527,6535
and|6536,6539
Vicodin|6540,6547
have|6548,6552
Tylenol|6553,6560
as|6561,6563
an|6564,6566
active|6567,6573
ingredient|6574,6584
so|6585,6587
do|6588,6590
<EOL>|6591,6592
not|6592,6595
take|6596,6600
these|6601,6606
meds|6607,6611
with|6612,6616
additional|6617,6627
Tylenol|6628,6635
.|6635,6636
<EOL>|6637,6638
4.|6638,6640
Take|6641,6645
prescription|6646,6658
pain|6659,6663
medications|6664,6675
for|6676,6679
pain|6680,6684
not|6685,6688
relieved|6689,6697
by|6698,6700
<EOL>|6701,6702
tylenol|6702,6709
.|6709,6710
<EOL>|6711,6712
5.|6712,6714
Take|6715,6719
your|6720,6724
antibiotic|6725,6735
as|6736,6738
prescribed|6739,6749
.|6749,6750
<EOL>|6751,6752
6.|6752,6754
Take|6755,6759
Colace|6760,6766
,|6766,6767
100|6768,6771
mg|6772,6774
by|6775,6777
mouth|6778,6783
2|6784,6785
times|6786,6791
per|6792,6795
day|6796,6799
,|6799,6800
while|6801,6806
taking|6807,6813
<EOL>|6814,6815
the|6815,6818
prescription|6819,6831
pain|6832,6836
medication|6837,6847
.|6847,6848
You|6849,6852
may|6853,6856
use|6857,6860
a|6861,6862
different|6863,6872
<EOL>|6873,6874
over-the|6874,6882
-|6882,6883
counter|6883,6890
stool|6891,6896
softener|6897,6905
if|6906,6908
you|6909,6912
wish|6913,6917
.|6917,6918
<EOL>|6919,6920
7.|6920,6922
Do|6923,6925
not|6926,6929
drive|6930,6935
or|6936,6938
operate|6939,6946
heavy|6947,6952
machinery|6953,6962
while|6963,6968
taking|6969,6975
any|6976,6979
<EOL>|6980,6981
narcotic|6981,6989
pain|6990,6994
medication|6995,7005
.|7005,7006
You|7007,7010
may|7011,7014
have|7015,7019
constipation|7020,7032
when|7033,7037
taking|7038,7044
<EOL>|7045,7046
narcotic|7046,7054
pain|7055,7059
medications|7060,7071
(|7072,7073
oxycodone|7073,7082
,|7082,7083
percocet|7084,7092
,|7092,7093
vicodin|7094,7101
,|7101,7102
<EOL>|7103,7104
hydrocodone|7104,7115
,|7115,7116
dilaudid|7117,7125
,|7125,7126
etc|7127,7130
.|7130,7131
)|7131,7132
;|7132,7133
you|7134,7137
should|7138,7144
continue|7145,7153
drinking|7154,7162
<EOL>|7163,7164
fluids|7164,7170
,|7170,7171
you|7172,7175
may|7176,7179
take|7180,7184
stool|7185,7190
softeners|7191,7200
,|7200,7201
and|7202,7205
should|7206,7212
eat|7213,7216
foods|7217,7222
that|7223,7227
<EOL>|7228,7229
are|7229,7232
high|7233,7237
in|7238,7240
fiber|7241,7246
.|7246,7247
<EOL>|7248,7249
8.|7249,7251
do|7252,7254
not|7255,7258
take|7259,7263
any|7264,7267
medicines|7268,7277
such|7278,7282
as|7283,7285
Motrin|7286,7292
,|7292,7293
Aspirin|7294,7301
,|7301,7302
Advil|7303,7308
or|7309,7311
<EOL>|7312,7313
Ibuprofen|7313,7322
etc|7323,7326
<EOL>|7326,7327
.|7327,7328
<EOL>|7329,7330
Call|7330,7334
the|7335,7338
office|7339,7345
IMMEDIATELY|7346,7357
if|7358,7360
you|7361,7364
have|7365,7369
any|7370,7373
of|7374,7376
the|7377,7380
following|7381,7390
:|7390,7391
<EOL>|7392,7393
1.|7393,7395
Signs|7396,7401
of|7402,7404
infection|7405,7414
:|7414,7415
fever|7416,7421
with|7422,7426
chills|7427,7433
,|7433,7434
increased|7435,7444
redness|7445,7452
,|7452,7453
<EOL>|7454,7455
welling|7455,7462
,|7462,7463
warmth|7464,7470
or|7471,7473
tenderness|7474,7484
at|7485,7487
the|7488,7491
surgical|7492,7500
site|7501,7505
,|7505,7506
or|7507,7509
unusual|7510,7517
<EOL>|7518,7519
drainage|7519,7527
from|7528,7532
the|7533,7536
incision|7537,7545
(|7545,7546
s|7546,7547
)|7547,7548
.|7548,7549
<EOL>|7550,7551
2|7551,7552
.|7552,7553
A|7554,7555
large|7556,7561
amount|7562,7568
of|7569,7571
bleeding|7572,7580
from|7581,7585
the|7586,7589
incision|7590,7598
(|7598,7599
s|7599,7600
)|7600,7601
or|7602,7604
drain|7605,7610
(|7610,7611
s|7611,7612
)|7612,7613
.|7613,7614
<EOL>|7615,7616
3.|7616,7618
Fever|7619,7624
greater|7625,7632
than|7633,7637
101.5|7638,7643
oF|7644,7646
<EOL>|7647,7648
4.|7648,7650
Severe|7651,7657
pain|7658,7662
NOT|7663,7666
relieved|7667,7675
by|7676,7678
your|7679,7683
medication|7684,7694
.|7694,7695
<EOL>|7696,7697
.|7697,7698
<EOL>|7699,7700
Return|7700,7706
to|7707,7709
the|7710,7713
ER|7714,7716
if|7717,7719
:|7719,7720
<EOL>|7721,7722
*|7722,7723
If|7724,7726
you|7727,7730
are|7731,7734
vomiting|7735,7743
and|7744,7747
can|7748,7751
not|7751,7754
keep|7755,7759
in|7760,7762
fluids|7763,7769
or|7770,7772
your|7773,7777
<EOL>|7778,7779
medications|7779,7790
.|7790,7791
<EOL>|7792,7793
*|7793,7794
If|7795,7797
you|7798,7801
have|7802,7806
shaking|7807,7814
chills|7815,7821
,|7821,7822
fever|7823,7828
greater|7829,7836
than|7837,7841
101.5|7842,7847
(|7848,7849
F|7849,7850
)|7850,7851
<EOL>|7852,7853
degrees|7853,7860
or|7861,7863
38|7864,7866
(|7867,7868
C|7868,7869
)|7869,7870
degrees|7871,7878
,|7878,7879
increased|7880,7889
redness|7890,7897
,|7897,7898
swelling|7899,7907
or|7908,7910
<EOL>|7911,7912
discharge|7912,7921
from|7922,7926
incision|7927,7935
,|7935,7936
chest|7937,7942
pain|7943,7947
,|7947,7948
shortness|7949,7958
of|7959,7961
breath|7962,7968
,|7968,7969
or|7970,7972
<EOL>|7973,7974
anything|7974,7982
else|7983,7987
that|7988,7992
is|7993,7995
troubling|7996,8005
you|8006,8009
.|8009,8010
<EOL>|8011,8012
*|8012,8013
Any|8014,8017
serious|8018,8025
change|8026,8032
in|8033,8035
your|8036,8040
symptoms|8041,8049
,|8049,8050
or|8051,8053
any|8054,8057
new|8058,8061
symptoms|8062,8070
that|8071,8075
<EOL>|8076,8077
concern|8077,8084
you|8085,8088
.|8088,8089
<EOL>|8090,8091
<EOL>|8091,8092
<EOL>|8093,8094
Followup|8094,8102
Instructions|8103,8115
:|8115,8116
<EOL>|8116,8117
_|8117,8118
_|8118,8119
_|8119,8120
<EOL>|8120,8121

