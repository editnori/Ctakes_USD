 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|52,61|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|52,61|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|52,66|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|86,95|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|86,95|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|86,100|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|142,145|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|153,160|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|153,160|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|162,170|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|173,182|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|173,182|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|173,182|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|188,197|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|188,197|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|188,197|true|false|false|C0020517|Hypersensitivity|Allergies
Event|Event|SIMPLE_SEGMENT|206,210|false|false|false|||File
Finding|Functional Concept|SIMPLE_SEGMENT|206,210|false|false|false|C0016094;C1522646;C1555017|File (record);Filed;URL Scheme - File|File
Finding|Intellectual Product|SIMPLE_SEGMENT|206,210|false|false|false|C0016094;C1522646;C1555017|File (record);Filed;URL Scheme - File|File
Event|Event|SIMPLE_SEGMENT|213,222|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|213,222|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|231,246|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|237,246|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|237,246|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|237,246|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|248,253|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|248,253|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|248,258|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|248,258|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|254,258|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|254,258|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|254,258|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|254,258|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|261,266|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|279,297|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|288,297|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|288,297|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|288,297|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|288,297|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|288,297|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|313,331|false|false|false|||pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|313,331|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Event|Event|SIMPLE_SEGMENT|342,349|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|342,349|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|342,349|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|342,349|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|342,352|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|342,368|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|342,368|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|353,360|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|353,360|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|353,368|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|361,368|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|371,378|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|371,381|false|false|false|C0262926|Medical History|HISTORY OF
Finding|Idea or Concept|SIMPLE_SEGMENT|382,392|true|false|false|C0449450|Presentation|PRESENTING
Event|Event|SIMPLE_SEGMENT|393,400|false|false|false|||ILLNESS
Finding|Sign or Symptom|SIMPLE_SEGMENT|393,400|false|false|false|C0221423|Illness (finding)|ILLNESS
Finding|Finding|SIMPLE_SEGMENT|419,423|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|429,449|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|440,449|false|false|false|C0003864|Arthritis|arthritis
Event|Event|SIMPLE_SEGMENT|440,449|false|false|false|||arthritis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|451,456|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|SIMPLE_SEGMENT|457,464|false|false|false|||holiday
Event|Event|SIMPLE_SEGMENT|457,464|false|false|false|C0019843|Holidays|holiday
Event|Event|SIMPLE_SEGMENT|478,483|false|false|false|||brief
Finding|Intellectual Product|SIMPLE_SEGMENT|478,483|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|SIMPLE_SEGMENT|484,499|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|484,499|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|516,528|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|516,528|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|530,538|false|false|false|||returned
Event|Event|SIMPLE_SEGMENT|551,559|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|551,559|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|SIMPLE_SEGMENT|565,573|false|false|false|C0332148|Probable diagnosis|probable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|574,581|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|574,581|false|true|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|574,591|false|true|false|C0007177|Cardiac Tamponade|cardiac tamponade
Event|Event|SIMPLE_SEGMENT|582,591|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|582,591|false|true|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|582,591|false|true|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|609,627|false|false|false|||pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|609,627|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Drug|Substance|SIMPLE_SEGMENT|633,638|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|633,638|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|633,638|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|633,648|false|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|639,648|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|639,648|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|639,648|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|658,666|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|658,666|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|658,666|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|658,666|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Body Substance|SIMPLE_SEGMENT|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|693,705|false|false|false|||hospitalized
Finding|Intellectual Product|SIMPLE_SEGMENT|725,730|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Sign or Symptom|SIMPLE_SEGMENT|731,751|false|false|false|C0008033|Pleuritic pain|pleuritic chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|741,746|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|741,746|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|741,751|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|741,751|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|747,751|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|747,751|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|759,762|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|759,762|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|763,771|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Event|Event|SIMPLE_SEGMENT|763,771|false|false|false|||duration
Event|Event|SIMPLE_SEGMENT|779,786|false|false|false|||context
Finding|Idea or Concept|SIMPLE_SEGMENT|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|SIMPLE_SEGMENT|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|SIMPLE_SEGMENT|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Event|Event|SIMPLE_SEGMENT|790,803|false|false|false|||constellation
Event|Event|SIMPLE_SEGMENT|807,814|false|false|false|||fatigue
Finding|Sign or Symptom|SIMPLE_SEGMENT|807,814|false|false|false|C0015672|Fatigue|fatigue
Event|Event|SIMPLE_SEGMENT|816,823|false|false|false|||malaise
Finding|Sign or Symptom|SIMPLE_SEGMENT|816,823|false|false|false|C0231218|Malaise|malaise
Attribute|Clinical Attribute|SIMPLE_SEGMENT|831,842|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|SIMPLE_SEGMENT|831,842|false|false|false|||respiratory
Finding|Body Substance|SIMPLE_SEGMENT|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|843,851|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|843,851|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|843,851|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|SIMPLE_SEGMENT|872,877|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|872,877|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|872,877|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|872,877|false|false|false|C0010200|Coughing|cough
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|885,888|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|885,888|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|885,888|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|885,888|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|SIMPLE_SEGMENT|889,899|false|false|false|||exonerated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|900,909|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|900,909|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|900,909|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|900,918|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|910,918|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|910,918|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|910,918|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|SIMPLE_SEGMENT|920,929|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|930,941|false|false|false|C0031050|Pericardial sac structure|pericardium
Event|Event|SIMPLE_SEGMENT|952,960|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|967,972|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|985,997|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|985,997|false|false|false|||pericarditis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|999,1002|false|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|999,1002|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|999,1002|false|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|1003,1011|false|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|1030,1040|false|false|false|||elevations
Event|Event|SIMPLE_SEGMENT|1044,1051|false|false|false|||keeping
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1057,1069|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|1057,1069|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|1071,1085|false|false|false|||Echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1071,1085|false|false|false|C0013516|Echocardiography|Echocardiogram
Event|Event|SIMPLE_SEGMENT|1087,1096|false|false|false|||confirmed
Event|Event|SIMPLE_SEGMENT|1102,1110|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|1122,1130|false|false|false|||features
Event|Event|SIMPLE_SEGMENT|1134,1143|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|1134,1143|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1134,1143|false|false|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|1149,1160|false|false|false|||appreciated
Event|Event|SIMPLE_SEGMENT|1169,1179|false|false|false|||discharged
Finding|Idea or Concept|SIMPLE_SEGMENT|1189,1192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1189,1192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|1198,1207|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1198,1207|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|1198,1207|false|false|false|||ibuprofen
Drug|Organic Chemical|SIMPLE_SEGMENT|1223,1233|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1223,1233|false|false|false|C0009262|colchicine|colchicine
Event|Event|SIMPLE_SEGMENT|1223,1233|false|false|false|||colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1241,1244|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1241,1244|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1241,1244|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|1241,1244|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|1241,1244|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|1253,1264|false|false|false|||persistence
Finding|Mental Process|SIMPLE_SEGMENT|1253,1264|false|false|false|C0546816|Persistence|persistence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1268,1273|false|false|false|C1446899|minor (disease)|minor
Event|Event|SIMPLE_SEGMENT|1268,1273|false|false|false|||minor
Finding|Gene or Genome|SIMPLE_SEGMENT|1268,1273|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1284,1289|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1284,1289|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1290,1294|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1290,1294|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1290,1294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1290,1294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1302,1307|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|1311,1317|false|false|false|||worsen
Event|Event|SIMPLE_SEGMENT|1342,1351|false|false|false|||tolerable
Event|Event|SIMPLE_SEGMENT|1368,1375|false|false|false|||evening
Event|Event|SIMPLE_SEGMENT|1384,1391|false|false|false|||evolved
Event|Event|SIMPLE_SEGMENT|1395,1401|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|1395,1401|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1395,1401|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|1403,1414|false|false|false|||unrelenting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1415,1419|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1415,1419|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1415,1419|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1415,1419|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1431,1441|false|false|false|C0230134|Structure of precordium|precordium
Event|Event|SIMPLE_SEGMENT|1442,1449|false|false|false|||likened
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1462,1470|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1462,1470|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1462,1470|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|SIMPLE_SEGMENT|1471,1475|false|false|false|||pads
Event|Event|SIMPLE_SEGMENT|1501,1506|false|false|false|||notes
Finding|Finding|SIMPLE_SEGMENT|1509,1512|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1509,1512|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1535,1540|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1535,1540|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1541,1545|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1541,1545|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1541,1545|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1541,1545|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1552,1556|false|false|false|||goes
Finding|Social Behavior|SIMPLE_SEGMENT|1557,1565|false|false|false|C0019421|Heterosexuality|straight
Finding|Intellectual Product|SIMPLE_SEGMENT|1583,1587|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1595,1603|false|false|false|||dyspneic
Finding|Finding|SIMPLE_SEGMENT|1595,1603|false|false|false|C0277854|dyspneic|dyspneic
Event|Event|SIMPLE_SEGMENT|1605,1614|false|false|false|||prompting
Event|Event|SIMPLE_SEGMENT|1622,1626|false|false|false|||seek
Event|Activity|SIMPLE_SEGMENT|1627,1631|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|1627,1631|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|1627,1631|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|1627,1631|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|1636,1643|false|false|false|||arrived
Event|Event|SIMPLE_SEGMENT|1651,1662|false|false|false|||hypotensive
Finding|Pathologic Function|SIMPLE_SEGMENT|1651,1662|false|false|false|C0857353|Hypotensive|hypotensive
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1668,1671|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1668,1671|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1668,1671|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|1668,1671|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|1668,1671|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1668,1671|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|SIMPLE_SEGMENT|1682,1687|false|false|false|||range
Finding|Intellectual Product|SIMPLE_SEGMENT|1682,1687|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Event|Event|SIMPLE_SEGMENT|1707,1718|false|false|false|||tachycardic
Finding|Intellectual Product|SIMPLE_SEGMENT|1726,1730|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1731,1742|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|1731,1751|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|1743,1751|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|1743,1751|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|1743,1751|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|1757,1768|false|false|false|||oxygenation
Finding|Cell Function|SIMPLE_SEGMENT|1757,1768|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1757,1768|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Event|Event|SIMPLE_SEGMENT|1773,1783|false|false|false|||acceptable
Drug|Substance|SIMPLE_SEGMENT|1821,1826|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|1821,1826|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|1821,1826|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|1843,1852|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|1843,1852|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1843,1852|false|false|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|1864,1872|false|false|false|||confines
Finding|Intellectual Product|SIMPLE_SEGMENT|1876,1880|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|1881,1888|false|false|false|||windows
Event|Event|SIMPLE_SEGMENT|1900,1914|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1900,1914|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|1916,1934|false|false|false|||Pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1916,1934|false|false|false|C0191234|Pericardiocentesis|Pericardiocentesis
Event|Event|SIMPLE_SEGMENT|1935,1942|false|false|false|||yielded
Finding|Body Substance|SIMPLE_SEGMENT|1961,1973|false|false|false|C0682554|Serous fluid|serous fluid
Drug|Substance|SIMPLE_SEGMENT|1968,1973|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|1968,1973|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1980,1991|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1980,1991|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Drug|Substance|SIMPLE_SEGMENT|1992,1997|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|1992,1997|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|1992,1997|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|2002,2008|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|2010,2022|false|false|false|||Hemodynamics
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2010,2022|false|false|false|C0019010|Hemodynamics|Hemodynamics
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2010,2022|false|false|false|C4281788|hemodynamics (procedure)|Hemodynamics
Event|Event|SIMPLE_SEGMENT|2031,2039|false|false|false|||improved
Event|Activity|SIMPLE_SEGMENT|2044,2051|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|2044,2051|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2044,2051|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Body Substance|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|2082,2104|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|SIMPLE_SEGMENT|2098,2104|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|2098,2104|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|SIMPLE_SEGMENT|2113,2117|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|SIMPLE_SEGMENT|2121,2129|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|2121,2129|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2130,2141|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2130,2150|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|2142,2150|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2142,2150|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2142,2150|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|2152,2161|false|false|false|||requiring
Drug|Organic Chemical|SIMPLE_SEGMENT|2191,2196|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2191,2196|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|2191,2196|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|2215,2229|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2215,2229|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|2234,2241|false|false|false|||limited
Event|Event|SIMPLE_SEGMENT|2261,2271|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|2261,2271|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|2261,2274|false|false|false|C0332299|Suggestive of|suggestive of
Event|Event|SIMPLE_SEGMENT|2291,2299|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|2308,2311|false|false|false|||CCU
Finding|Body Substance|SIMPLE_SEGMENT|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2321,2326|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|2327,2337|false|false|false|||resurgence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2341,2345|false|false|false|C0080151|Simian Acquired Immunodeficiency Syndrome|said
Event|Event|SIMPLE_SEGMENT|2341,2345|false|false|false|||said
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2346,2351|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2346,2351|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2346,2356|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2346,2356|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2352,2356|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2352,2356|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2352,2356|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2352,2356|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2362,2369|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|2362,2369|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2362,2369|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|2373,2382|false|false|false|||improving
Finding|Functional Concept|SIMPLE_SEGMENT|2387,2397|false|false|false|C1524062|Additional|additional
Event|Event|SIMPLE_SEGMENT|2409,2416|false|false|false|||drained
Finding|Finding|SIMPLE_SEGMENT|2421,2441|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2426,2433|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2426,2433|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2426,2433|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2426,2433|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2426,2433|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2426,2441|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2434,2441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2434,2441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2434,2441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2443,2463|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PAST MEDICAL HISTORY
Event|Event|SIMPLE_SEGMENT|2448,2455|false|false|false|||MEDICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2448,2455|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Idea or Concept|SIMPLE_SEGMENT|2448,2455|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Intellectual Product|SIMPLE_SEGMENT|2448,2455|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2448,2455|false|false|false|C0199168|Medical service|MEDICAL
Finding|Finding|SIMPLE_SEGMENT|2448,2463|false|false|false|C0262926|Medical History|MEDICAL HISTORY
Event|Event|SIMPLE_SEGMENT|2456,2463|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|2456,2463|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|2456,2463|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|2456,2463|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2468,2475|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2468,2475|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|SIMPLE_SEGMENT|2476,2483|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2476,2483|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2476,2483|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2476,2483|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2488,2500|false|false|false|C0031046|Pericarditis|Pericarditis
Event|Event|SIMPLE_SEGMENT|2488,2500|false|false|false|||Pericarditis
Finding|Idea or Concept|SIMPLE_SEGMENT|2505,2510|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2513,2525|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|2513,2525|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2528,2540|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|SIMPLE_SEGMENT|2528,2540|false|false|false|||Dyslipidemia
Event|Event|SIMPLE_SEGMENT|2552,2555|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|2552,2555|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2560,2580|false|false|false|C0003873|Rheumatoid Arthritis|Rheumatoid arthritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2571,2580|false|false|false|C0003864|Arthritis|arthritis
Event|Event|SIMPLE_SEGMENT|2571,2580|false|false|false|||arthritis
Finding|Functional Concept|SIMPLE_SEGMENT|2591,2600|false|false|false|C0332663|Traumatic|traumatic
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2601,2604|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2601,2604|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2601,2604|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|2601,2604|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|2607,2622|false|false|false|||Cholecystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2607,2622|false|false|false|C0008320|Cholecystectomy procedure|Cholecystectomy
Event|Event|SIMPLE_SEGMENT|2625,2637|false|false|false|||Appendectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2625,2637|false|false|false|C0003611;C0003612|Appendectomy;Appendectomy; for ruptured appendix with abscess or generalized peritonitis|Appendectomy
Event|Event|SIMPLE_SEGMENT|2640,2653|false|false|false|||Tonsillectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2640,2653|false|false|false|C0040423|Tonsillectomy|Tonsillectomy
Finding|Functional Concept|SIMPLE_SEGMENT|2656,2660|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2656,2666|false|false|false|C0230366|Structure of left wrist|Left wrist
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2661,2666|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2661,2666|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2661,2681|false|false|false|C0845620|Wrist reconstruction|wrist reconstruction
Event|Event|SIMPLE_SEGMENT|2667,2681|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|2667,2681|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2667,2681|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Finding|Functional Concept|SIMPLE_SEGMENT|2684,2689|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2684,2702|false|false|false|C0828608|Right tendinous cuff|Right rotator cuff
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2690,2702|false|false|false|C0085515|Rotator Cuff|rotator cuff
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2698,2702|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|SIMPLE_SEGMENT|2698,2702|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Event|Event|SIMPLE_SEGMENT|2703,2717|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|2703,2717|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2703,2717|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Finding|Functional Concept|SIMPLE_SEGMENT|2722,2728|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2722,2736|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2729,2736|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2729,2736|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2729,2736|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2729,2736|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2742,2748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2742,2748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2742,2748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2742,2748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2742,2756|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2749,2756|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2749,2756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2749,2756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2749,2756|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2758,2774|false|false|false|C0424909|Family history with explicit context pertaining to father|paternal history
Event|Event|SIMPLE_SEGMENT|2767,2774|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2767,2777|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2790,2799|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|SIMPLE_SEGMENT|2790,2799|false|false|false|||carcinoma
Finding|Finding|SIMPLE_SEGMENT|2801,2809|false|false|false|C1858460|Maternal|Maternal
Finding|Finding|SIMPLE_SEGMENT|2801,2817|false|false|false|C0559473|maternal history|Maternal history
Event|Event|SIMPLE_SEGMENT|2810,2817|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2810,2820|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2821,2829|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|2821,2829|false|false|false|||diabetes
Event|Event|SIMPLE_SEGMENT|2835,2843|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2835,2843|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2835,2843|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2835,2843|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2835,2848|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2835,2848|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2844,2848|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2844,2848|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2844,2848|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2850,2859|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|SIMPLE_SEGMENT|2860,2868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2860,2868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2860,2868|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2860,2880|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2860,2880|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|2869,2880|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|2869,2880|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2869,2880|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|2931,2933|false|false|false|||HR
Event|Event|SIMPLE_SEGMENT|2961,2968|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2961,2968|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2961,2968|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2970,2975|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2970,2975|false|false|false|||obese
Finding|Finding|SIMPLE_SEGMENT|2976,2980|false|false|false|C1706180|Male Gender|male
Finding|Intellectual Product|SIMPLE_SEGMENT|2984,2988|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|2992,3000|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|2992,3000|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3001,3012|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|3001,3021|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|3013,3021|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|3013,3021|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3013,3021|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3026,3031|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3033,3042|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3043,3050|false|false|false|||sclerae
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3052,3062|false|false|false|C0521367|Oropharyngeal|Oropharynx
Event|Event|SIMPLE_SEGMENT|3063,3068|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3063,3068|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3073,3077|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3079,3082|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3079,3082|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3086,3096|false|false|false|C0024687|Mandible|mandibular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3106,3113|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3106,3113|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|3128,3135|false|false|false|||regular
Finding|Gene or Genome|SIMPLE_SEGMENT|3141,3145|false|false|false|C1514917|Retinoic Acid Response Element|rare
Event|Event|SIMPLE_SEGMENT|3146,3152|false|false|false|||ectopy
Event|Event|SIMPLE_SEGMENT|3172,3180|false|false|false|||confines
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3184,3188|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3184,3188|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|3184,3188|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3184,3196|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|SIMPLE_SEGMENT|3189,3196|false|false|false|||habitus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3205,3216|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3205,3216|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Finding|Finding|SIMPLE_SEGMENT|3205,3220|false|false|false|C0232267|Pericardial friction rub|pericardial rub
Event|Event|SIMPLE_SEGMENT|3217,3220|false|false|false|||rub
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3222,3233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3222,3233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Drug|Substance|SIMPLE_SEGMENT|3234,3239|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|3234,3239|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|3234,3239|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Body Substance|SIMPLE_SEGMENT|3245,3265|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|SIMPLE_SEGMENT|3260,3265|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|3260,3265|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3260,3265|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3267,3274|false|false|false|C0038293|Sternum|Sternal
Finding|Finding|SIMPLE_SEGMENT|3267,3285|false|false|false|C0241246|tender sternum on palpation|Sternal tenderness
Event|Event|SIMPLE_SEGMENT|3275,3285|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3275,3285|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3275,3285|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3289,3294|false|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|3311,3318|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|3311,3318|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3311,3318|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|3323,3332|false|false|false|||tachypnea
Finding|Finding|SIMPLE_SEGMENT|3323,3332|false|false|false|C0231835|Tachypnea|tachypnea
Event|Event|SIMPLE_SEGMENT|3336,3343|false|false|false|||slowing
Event|Event|SIMPLE_SEGMENT|3353,3361|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|3353,3361|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|3366,3374|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3366,3374|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3388,3392|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3388,3392|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3388,3392|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|3388,3392|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|3393,3399|false|false|false|||fields
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3404,3411|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3404,3411|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3404,3411|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3404,3411|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3413,3418|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3413,3418|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3420,3424|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3420,3424|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3439,3450|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|3452,3456|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|3452,3456|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3452,3456|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3458,3462|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3463,3471|false|false|false|||perfused
Finding|Finding|SIMPLE_SEGMENT|3473,3489|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|3476,3483|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|3476,3489|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3484,3489|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3484,3489|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3484,3489|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3493,3498|false|false|false|C0022742|Knee|knees
Anatomy|Body System|SIMPLE_SEGMENT|3503,3507|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3503,3507|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3503,3507|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3503,3507|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3503,3507|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3503,3507|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3509,3516|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|3509,3516|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3527,3533|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3527,3540|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|3527,3540|false|false|false|C4551518|Venous stasis|venous stasis
Event|Event|SIMPLE_SEGMENT|3534,3540|false|false|false|||stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|3534,3540|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3534,3551|false|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3541,3551|false|false|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|3541,3551|false|false|false|||dermatitis
Drug|Food|SIMPLE_SEGMENT|3556,3562|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|3556,3562|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3556,3562|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3556,3562|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3564,3570|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|SIMPLE_SEGMENT|3571,3577|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3571,3577|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3571,3577|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3571,3577|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|3591,3600|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3591,3600|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3591,3600|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|SIMPLE_SEGMENT|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3624,3633|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|SIMPLE_SEGMENT|3634,3642|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3634,3642|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3634,3642|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3634,3654|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3634,3654|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|3643,3654|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3643,3654|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3643,3654|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3692,3699|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3692,3699|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3692,3699|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3701,3706|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3701,3706|false|false|false|||obese
Finding|Finding|SIMPLE_SEGMENT|3707,3711|false|false|false|C1706180|Male Gender|male
Finding|Intellectual Product|SIMPLE_SEGMENT|3715,3719|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|3723,3731|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|3723,3731|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3732,3743|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|3732,3752|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|3744,3752|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|3744,3752|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3744,3752|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3757,3762|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3764,3773|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3774,3781|false|false|false|||sclerae
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3783,3793|false|false|false|C0521367|Oropharyngeal|Oropharynx
Event|Event|SIMPLE_SEGMENT|3794,3799|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3794,3799|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3804,3808|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3804,3808|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3804,3808|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3810,3813|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3810,3813|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|3818,3829|false|false|false|||appreciated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3833,3840|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3833,3840|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|SIMPLE_SEGMENT|3849,3853|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|3849,3853|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3849,3853|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|3858,3864|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|3858,3864|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3858,3864|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3895,3899|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3895,3899|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|3895,3899|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3895,3907|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|SIMPLE_SEGMENT|3900,3907|false|false|false|||habitus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3912,3923|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3912,3923|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Finding|Finding|SIMPLE_SEGMENT|3912,3927|true|false|false|C0232267|Pericardial friction rub|pericardial rub
Event|Event|SIMPLE_SEGMENT|3924,3927|false|false|false|||rub
Event|Event|SIMPLE_SEGMENT|3928,3939|false|false|false|||appreciated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3943,3948|false|false|false|C0024109|Lung|LUNGS
Finding|Finding|SIMPLE_SEGMENT|3950,3959|false|false|false|C0392756;C0442797|Decreasing;Reduced|Decreased
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3960,3971|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3960,3978|false|false|false|C4050166||respiratory effort
Finding|Finding|SIMPLE_SEGMENT|3960,3978|false|false|false|C0425466|Respiratory effort|respiratory effort
Event|Event|SIMPLE_SEGMENT|3972,3978|false|false|false|||effort
Finding|Organism Function|SIMPLE_SEGMENT|3972,3978|false|false|false|C0015264|Exertion|effort
Event|Event|SIMPLE_SEGMENT|3979,3987|false|false|false|||compared
Finding|Organism Function|SIMPLE_SEGMENT|4002,4012|false|false|false|C0231800|Expiration, Respiratory|Expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|4002,4021|false|false|false|C0231875|Expiratory wheezing|Expiratory wheezing
Event|Event|SIMPLE_SEGMENT|4013,4021|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|4013,4021|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|4036,4044|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|4036,4044|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4047,4054|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4047,4054|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|4047,4054|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4047,4054|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4056,4061|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|4056,4061|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4063,4067|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4063,4067|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4097,4108|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|SIMPLE_SEGMENT|4110,4114|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|4110,4114|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4110,4114|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|4116,4120|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4121,4129|false|false|false|||perfused
Finding|Finding|SIMPLE_SEGMENT|4136,4152|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|4139,4146|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|4139,4152|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4147,4152|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4147,4152|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4147,4152|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4156,4161|false|false|false|C0022742|Knee|knees
Anatomy|Body System|SIMPLE_SEGMENT|4166,4170|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4166,4170|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4166,4170|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|4166,4170|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|4166,4170|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|4166,4170|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|4172,4179|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|4172,4179|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4180,4186|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4180,4193|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4180,4193|false|false|false|C4551518|Venous stasis|venous stasis
Event|Event|SIMPLE_SEGMENT|4187,4193|false|false|false|||stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4187,4193|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4187,4204|false|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4194,4204|false|false|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|4194,4204|false|false|false|||dermatitis
Drug|Food|SIMPLE_SEGMENT|4209,4215|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|4209,4215|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|4209,4215|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|4209,4215|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4217,4223|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|SIMPLE_SEGMENT|4224,4230|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4224,4230|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4224,4230|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4224,4230|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|4244,4253|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|4244,4253|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|4244,4253|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Procedure|Health Care Activity|SIMPLE_SEGMENT|4297,4306|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4307,4311|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4307,4311|false|false|false|C0587081|Laboratory test finding|LABS
Anatomy|Cell|SIMPLE_SEGMENT|4343,4346|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4353,4356|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4353,4356|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4353,4356|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4362,4365|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4362,4365|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|4362,4365|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|4362,4365|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4362,4365|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|4371,4374|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4371,4374|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4371,4374|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|4380,4383|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4380,4383|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4380,4383|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4380,4383|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4380,4383|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4388,4391|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4388,4391|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4388,4391|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4388,4391|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4388,4391|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4388,4391|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4397,4401|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4397,4401|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Finding|Body Substance|SIMPLE_SEGMENT|4453,4459|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4475,4478|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|4475,4478|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|4475,4478|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4590,4593|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4590,4593|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4590,4593|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4617,4624|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4617,4624|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4617,4624|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4630,4634|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|4630,4634|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4630,4634|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|4630,4634|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4630,4634|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|4650,4656|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4650,4656|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4650,4656|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|4662,4671|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4662,4671|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4662,4671|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4676,4684|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|4676,4684|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|4676,4684|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4676,4684|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4695,4698|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4695,4698|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|4695,4698|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|4695,4698|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|4695,4698|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4703,4708|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4703,4712|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4703,4712|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4703,4712|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4709,4712|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4709,4712|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|4709,4712|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|4709,4712|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|4730,4737|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4730,4737|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4730,4737|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4743,4752|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Event|Event|SIMPLE_SEGMENT|4757,4766|false|false|false|||MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4757,4766|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Organic Chemical|SIMPLE_SEGMENT|4813,4820|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4813,4820|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Event|Event|SIMPLE_SEGMENT|4813,4820|false|false|false|||LACTATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4813,4820|false|false|false|C0202115|Lactic acid measurement|LACTATE
Anatomy|Tissue|SIMPLE_SEGMENT|4837,4844|false|false|false|C0032225|Pleura|PLEURAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4837,4844|false|false|false|C0032226|Pleural Diseases|PLEURAL
Finding|Body Substance|SIMPLE_SEGMENT|4837,4850|false|false|false|C0225778|Pleural fluid|PLEURAL FLUID
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4837,4850|false|false|false|C2242629|Pleural fluid analysis|PLEURAL FLUID
Drug|Substance|SIMPLE_SEGMENT|4845,4850|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|4845,4850|false|false|false|C1546638|Fluid Specimen Code|FLUID
Event|Event|SIMPLE_SEGMENT|4851,4858|false|false|false|||STUDIES
Procedure|Research Activity|SIMPLE_SEGMENT|4851,4858|false|false|false|C0947630|Scientific Study|STUDIES
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4864,4869|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|Polys
Finding|Body Substance|SIMPLE_SEGMENT|4874,4880|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Event|Event|SIMPLE_SEGMENT|4894,4901|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4894,4901|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4894,4901|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|4916,4919|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4916,4919|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|SIMPLE_SEGMENT|4924,4928|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4924,4935|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4929,4935|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|4939,4945|false|false|false|||normal
Finding|Social Behavior|SIMPLE_SEGMENT|4959,4967|false|false|false|C0678975|inferiority|inferior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4959,4977|false|false|false|C0042458;C4266635|Abdomen>Vena cava.inferior;Inferior vena cava structure|inferior vena cava
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4968,4972|false|false|false|C0447122|Structure of vein of trunk|vena
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4968,4977|false|false|false|C0042460;C4266402|Chest+Abdomen>Vena cava.superior &or Vena cava.inferior;Vena caval structure|vena cava
Finding|Gene or Genome|SIMPLE_SEGMENT|4973,4977|false|false|false|C1413046|CA5A gene|cava
Event|Event|SIMPLE_SEGMENT|4982,4989|false|false|false|||dilated
Finding|Finding|SIMPLE_SEGMENT|4982,4989|false|false|false|C0700124|Dilated|dilated
Finding|Functional Concept|SIMPLE_SEGMENT|5017,5021|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5022,5033|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|5039,5048|false|false|false|||thickness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5063,5069|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5063,5069|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5063,5069|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5097,5102|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|5097,5102|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|5097,5102|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|SIMPLE_SEGMENT|5114,5120|false|false|false|||assess
Finding|Functional Concept|SIMPLE_SEGMENT|5130,5134|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5135,5146|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|5147,5155|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5157,5164|false|false|false|C0282416|Overall Publication Type|Overall
Finding|Functional Concept|SIMPLE_SEGMENT|5165,5169|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5170,5181|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5182,5190|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5191,5199|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|5203,5209|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|5233,5237|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Physiologic Function|SIMPLE_SEGMENT|5233,5258|false|false|false|C2733342|Left ventricular ejection|left ventricular ejection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5238,5249|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Physiologic Function|SIMPLE_SEGMENT|5238,5258|false|false|false|C2733340|Ventricular ejection|ventricular ejection
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5250,5258|false|false|false|C0812388|Ejection time|ejection
Event|Event|SIMPLE_SEGMENT|5250,5258|false|false|false|||ejection
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5250,5258|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5250,5258|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Event|Event|SIMPLE_SEGMENT|5259,5267|false|false|false|||fraction
Finding|Intellectual Product|SIMPLE_SEGMENT|5259,5267|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Finding|Functional Concept|SIMPLE_SEGMENT|5277,5281|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5277,5307|false|false|false|C4050538||Left ventricular cardiac index
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5282,5293|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5294,5301|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|5294,5301|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Finding|SIMPLE_SEGMENT|5294,5307|false|false|false|C0428776|Cardiac index|cardiac index
Event|Event|SIMPLE_SEGMENT|5302,5307|false|false|false|||index
Finding|Idea or Concept|SIMPLE_SEGMENT|5302,5307|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|SIMPLE_SEGMENT|5302,5307|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Event|Event|SIMPLE_SEGMENT|5311,5317|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5339,5350|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5339,5364|true|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5351,5364|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5351,5364|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5358,5364|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|5358,5364|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|5358,5364|true|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|5368,5372|false|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|5381,5386|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5381,5405|false|false|false|C0503854|Cavity of right ventricle|right ventricular cavity
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5381,5410|false|false|false|C0455865|Right ventricular cavity size|right ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5387,5398|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5387,5405|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5399,5405|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5399,5405|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5399,5405|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5406,5410|false|false|false|||size
Finding|Functional Concept|SIMPLE_SEGMENT|5423,5427|false|false|false|C0332296|Free of (attribute)|free
Event|Event|SIMPLE_SEGMENT|5434,5440|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5434,5440|false|false|false|C0026597|Motion|motion
Finding|Finding|SIMPLE_SEGMENT|5451,5459|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|5451,5459|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|SIMPLE_SEGMENT|5460,5476|false|false|false|||interventricular
Event|Event|SIMPLE_SEGMENT|5484,5490|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5484,5490|false|false|false|C0026597|Motion|motion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5496,5502|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5496,5508|false|false|false|C0037197|Structure of sinus of Valsalva|aortic sinus
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5503,5508|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5503,5508|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|5503,5508|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5503,5508|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|5509,5517|false|false|false|||diameter
Event|Event|SIMPLE_SEGMENT|5521,5527|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|5532,5538|false|false|false|||gender
Finding|Functional Concept|SIMPLE_SEGMENT|5552,5561|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5552,5567|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5562,5567|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|5562,5567|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Finding|SIMPLE_SEGMENT|5562,5576|false|false|false|C0579133|Aortic diameter|aorta diameter
Event|Event|SIMPLE_SEGMENT|5568,5576|false|false|false|||diameter
Event|Event|SIMPLE_SEGMENT|5581,5587|false|false|false|||gender
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5593,5599|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5593,5604|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5593,5604|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|5600,5604|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|5600,5604|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|SIMPLE_SEGMENT|5605,5613|false|false|false|||diameter
Event|Event|SIMPLE_SEGMENT|5617,5623|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|5637,5645|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5637,5645|true|false|false|C3887511|Evidence|evidence
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5654,5660|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5654,5665|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5654,5665|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|5661,5665|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|5661,5665|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5666,5677|false|false|false|C0003492;C0332886|Aortic coarctation;Coarctation|coarctation
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5666,5677|false|false|false|C0003492;C0332886|Aortic coarctation;Coarctation|coarctation
Event|Event|SIMPLE_SEGMENT|5666,5677|false|false|false|||coarctation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5683,5689|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5690,5695|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5696,5704|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5710,5716|false|false|false|||appear
Event|Event|SIMPLE_SEGMENT|5730,5736|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5751,5757|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5751,5763|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5751,5772|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5751,5772|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5751,5772|false|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5758,5763|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5764,5772|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5764,5772|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5786,5792|false|false|false|C0003483|Aorta|aortic
Event|Event|SIMPLE_SEGMENT|5793,5806|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5793,5806|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5793,5806|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5793,5806|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5812,5824|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5819,5824|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|5832,5836|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5837,5847|false|false|false|||visualized
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5854,5869|true|false|false|C0040960|Tricuspid valve structure|tricuspid valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5864,5869|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|5877,5881|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5882,5886|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5892,5901|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5892,5901|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5892,5901|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5902,5908|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5902,5908|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|5909,5917|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5909,5917|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5909,5926|false|false|false|C0871470|Systolic Pressure|systolic pressure
Event|Event|SIMPLE_SEGMENT|5918,5926|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5918,5926|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|5940,5949|false|false|false|||estimated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5964,5975|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5964,5975|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5964,5984|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|5964,5984|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|5976,5984|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5987,5992|false|false|false|||MICRO
Finding|Conceptual Entity|SIMPLE_SEGMENT|5987,5992|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|SIMPLE_SEGMENT|5987,5992|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5987,5992|false|false|false|C0085672|Microbiology procedure|MICRO
Drug|Substance|SIMPLE_SEGMENT|6013,6018|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|6013,6018|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|6013,6018|false|false|false|C1546638|Fluid Specimen Code|FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|6013,6024|false|false|false|C1546636|Fluid, Other|FLUID,OTHER
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6030,6041|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|PERICARDIAL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6030,6041|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|PERICARDIAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6030,6047|false|false|false|C0031039|Pericardial effusion|PERICARDIAL FLUID
Finding|Body Substance|SIMPLE_SEGMENT|6030,6047|false|false|false|C0225973|Pericardial fluid (substance)|PERICARDIAL FLUID
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6030,6047|false|false|false|C3854061|pericardial fluid analysis|PERICARDIAL FLUID
Drug|Substance|SIMPLE_SEGMENT|6042,6047|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|6042,6047|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|6042,6047|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6054,6064|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6054,6064|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6054,6064|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6059,6064|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|6059,6064|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6059,6064|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|6066,6071|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|6104,6109|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|6104,6109|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|6104,6109|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|6114,6131|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|SIMPLE_SEGMENT|6133,6143|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|6133,6143|false|false|false|||LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|6133,6143|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|6133,6143|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|SIMPLE_SEGMENT|6155,6174|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|SIMPLE_SEGMENT|6170,6174|false|false|false|||SEEN
Event|Activity|SIMPLE_SEGMENT|6206,6211|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|SIMPLE_SEGMENT|6206,6211|false|false|false|||smear
Finding|Functional Concept|SIMPLE_SEGMENT|6206,6211|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6206,6211|false|false|false|C0444186|Smear test|smear
Event|Event|SIMPLE_SEGMENT|6229,6235|false|false|false|||method
Finding|Functional Concept|SIMPLE_SEGMENT|6229,6235|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|SIMPLE_SEGMENT|6229,6235|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Event|Event|SIMPLE_SEGMENT|6260,6270|false|false|false|||hematology
Finding|Intellectual Product|SIMPLE_SEGMENT|6260,6270|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6260,6270|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|SIMPLE_SEGMENT|6290,6306|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6290,6312|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6290,6312|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6296,6301|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|6296,6301|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|SIMPLE_SEGMENT|6296,6306|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6296,6312|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|SIMPLE_SEGMENT|6302,6306|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|6302,6306|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6302,6312|false|false|false|C0007584|Cell Count|cell count
Event|Event|SIMPLE_SEGMENT|6307,6312|false|false|false|||count
Drug|Substance|SIMPLE_SEGMENT|6320,6325|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|6320,6325|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6326,6333|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6326,6333|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6326,6333|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6326,6333|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6326,6333|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|6356,6364|false|false|false|||Reported
Event|Event|SIMPLE_SEGMENT|6372,6376|false|false|false|||read
Event|Event|SIMPLE_SEGMENT|6396,6400|false|false|false|||53PM
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6409,6423|false|false|false|C0374989|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|STAPHYLOCOCCUS
Event|Event|SIMPLE_SEGMENT|6409,6423|false|false|false|||STAPHYLOCOCCUS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6425,6434|false|false|false|C0009118|Coagulase|COAGULASE
Drug|Enzyme|SIMPLE_SEGMENT|6425,6434|false|false|false|C0009118|Coagulase|COAGULASE
Anatomy|Cell|SIMPLE_SEGMENT|6450,6456|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Event|Event|SIMPLE_SEGMENT|6463,6468|false|false|false|||PLATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6475,6492|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6485,6492|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6485,6492|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6485,6492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6485,6492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6485,6492|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|6524,6532|false|false|false|||ISOLATED
Finding|Functional Concept|SIMPLE_SEGMENT|6539,6545|false|false|false|C0521033|Fungal|FUNGAL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6539,6553|false|false|false|C0200954|Mycology culture|FUNGAL CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6546,6553|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6546,6553|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6546,6553|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6546,6553|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6546,6553|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|6574,6578|false|false|false|||ACID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6574,6583|false|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|6579,6583|false|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Activity|SIMPLE_SEGMENT|6584,6589|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Event|Event|SIMPLE_SEGMENT|6584,6589|false|false|false|||SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|6584,6589|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6584,6589|false|false|false|C0444186|Smear test|SMEAR
Finding|Idea or Concept|SIMPLE_SEGMENT|6591,6596|false|false|false|C1546485|Diagnosis Type - Final|Final
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6612,6621|true|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|6617,6621|false|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Event|SIMPLE_SEGMENT|6622,6629|false|false|false|||BACILLI
Event|Event|SIMPLE_SEGMENT|6630,6634|false|false|false|||SEEN
Finding|Intellectual Product|SIMPLE_SEGMENT|6638,6644|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Event|Activity|SIMPLE_SEGMENT|6645,6650|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Event|Event|SIMPLE_SEGMENT|6645,6650|false|false|false|||SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|6645,6650|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6645,6650|false|false|false|C0444186|Smear test|SMEAR
Event|Event|SIMPLE_SEGMENT|6657,6661|false|false|false|||ACID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6657,6666|false|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|6662,6666|false|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6667,6674|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6667,6674|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6667,6674|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6667,6674|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6667,6674|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Body Substance|SIMPLE_SEGMENT|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|6692,6701|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|6702,6706|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6702,6706|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6736,6741|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6736,6741|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6736,6741|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|6742,6745|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|6752,6755|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6752,6755|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6752,6755|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6762,6765|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6762,6765|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|6762,6765|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6762,6765|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6772,6775|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6772,6775|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|6783,6786|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|6783,6786|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6783,6786|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6783,6786|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6783,6786|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|6790,6793|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6790,6793|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|6790,6793|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|6790,6793|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|6790,6793|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6790,6793|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|6799,6803|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6799,6803|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6829,6832|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6849,6854|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6849,6854|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6849,6854|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|6849,6862|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6849,6862|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6849,6862|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6855,6862|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|6855,6862|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6855,6862|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|6855,6862|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6855,6862|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6855,6862|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6909,6913|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6909,6913|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6909,6913|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6938,6943|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6938,6943|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6938,6943|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6944,6947|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6944,6947|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|6944,6947|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|6944,6947|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6944,6947|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6952,6955|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6952,6955|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|6952,6955|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|6952,6955|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6959,6966|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|6959,6966|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6994,6999|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6994,6999|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6994,6999|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6994,7007|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|7000,7007|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|7000,7007|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7000,7007|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7041,7046|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7041,7046|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7041,7046|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7047,7053|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|7047,7053|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7070,7075|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7070,7075|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7070,7075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7076,7079|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|7076,7079|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7076,7079|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7097,7102|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7097,7102|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7097,7102|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|7107,7110|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|7107,7110|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|7107,7110|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7107,7110|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7115,7119|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7115,7119|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7144,7148|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|7144,7148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|7144,7148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Intellectual Product|SIMPLE_SEGMENT|7157,7162|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|7163,7171|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7163,7178|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|7163,7178|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|7180,7187|false|false|false|||SUMMARY
Finding|Intellectual Product|SIMPLE_SEGMENT|7180,7187|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Finding|Finding|SIMPLE_SEGMENT|7217,7221|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7227,7247|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7238,7247|false|false|false|C0003864|Arthritis|arthritis
Event|Event|SIMPLE_SEGMENT|7238,7247|false|false|false|||arthritis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7249,7254|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|SIMPLE_SEGMENT|7255,7262|false|false|false|||holiday
Event|Event|SIMPLE_SEGMENT|7255,7262|false|false|false|C0019843|Holidays|holiday
Finding|Intellectual Product|SIMPLE_SEGMENT|7276,7281|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|SIMPLE_SEGMENT|7282,7297|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|7282,7297|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7314,7326|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|7314,7326|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|7328,7336|false|false|false|||returned
Finding|Idea or Concept|SIMPLE_SEGMENT|7348,7356|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7362,7373|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7362,7373|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7362,7382|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|7362,7382|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|7374,7382|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Finding|SIMPLE_SEGMENT|7389,7397|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|7398,7407|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|7398,7407|false|true|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7398,7407|false|true|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|7408,7418|false|false|false|||physiology
Finding|Physiologic Function|SIMPLE_SEGMENT|7408,7418|false|true|false|C0031843|physiological aspects|physiology
Event|Event|SIMPLE_SEGMENT|7437,7455|false|false|false|||pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7437,7455|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Event|Event|SIMPLE_SEGMENT|7465,7473|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|7465,7473|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|7465,7473|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|7465,7473|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7492,7503|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7492,7503|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7492,7512|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|7492,7512|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|7504,7512|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Drug|Substance|SIMPLE_SEGMENT|7521,7526|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|7521,7526|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7521,7536|false|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|7527,7536|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|7527,7536|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7527,7536|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|7542,7548|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|7550,7561|false|false|false|||complicated
Finding|Intellectual Product|SIMPLE_SEGMENT|7565,7570|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7584,7595|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|7584,7604|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|7596,7604|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|7596,7604|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|7596,7604|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|7609,7619|false|false|false|||CORONARIES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|7621,7628|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|7631,7635|false|false|false|||PUMP
Finding|Molecular Function|SIMPLE_SEGMENT|7631,7635|false|false|false|C1150186|matrix metalloproteinase 7 activity|PUMP
Event|Event|SIMPLE_SEGMENT|7658,7667|false|false|false|||structure
Event|Event|SIMPLE_SEGMENT|7672,7680|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|7684,7690|false|false|false|||RHYTHM
Finding|Finding|SIMPLE_SEGMENT|7684,7690|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Finding|Physiologic Function|SIMPLE_SEGMENT|7684,7690|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Event|Event|SIMPLE_SEGMENT|7692,7695|false|false|false|||NSR
Finding|Molecular Function|SIMPLE_SEGMENT|7692,7695|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|SIMPLE_SEGMENT|7692,7695|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7697,7700|false|false|false|C0235480;C0393911|Paroxysmal atrial fibrillation;Pure Autonomic Failure|pAF
Drug|Immunologic Factor|SIMPLE_SEGMENT|7697,7700|false|false|false|C0032172|Platelet Activating Factor|pAF
Drug|Organic Chemical|SIMPLE_SEGMENT|7697,7700|false|false|false|C0032172|Platelet Activating Factor|pAF
Event|Event|SIMPLE_SEGMENT|7697,7700|false|false|false|||pAF
Finding|Gene or Genome|SIMPLE_SEGMENT|7697,7700|false|false|false|C1537443|PCLAF gene|pAF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7697,7700|false|false|false|C0279389|doxorubicin/fluorouracil/melphalan protocol|pAF
Finding|Idea or Concept|SIMPLE_SEGMENT|7706,7718|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|7719,7725|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|7758,7768|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|7772,7781|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7772,7781|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|7772,7781|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|7788,7791|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|7796,7806|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7796,7806|false|false|false|C0009262|colchicine|colchicine
Event|Event|SIMPLE_SEGMENT|7796,7806|false|false|false|||colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7814,7817|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7814,7817|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7814,7817|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7814,7817|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7814,7817|false|false|false|C1332410|BID gene|BID
Finding|Functional Concept|SIMPLE_SEGMENT|7826,7838|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7839,7851|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|7839,7851|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|7863,7871|false|false|false|||continue
Drug|Organic Chemical|SIMPLE_SEGMENT|7873,7883|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7873,7883|false|false|false|C0009262|colchicine|colchicine
Event|Event|SIMPLE_SEGMENT|7873,7883|false|false|false|||colchicine
Drug|Organic Chemical|SIMPLE_SEGMENT|7917,7926|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7917,7926|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|7927,7934|false|false|false|||tapered
Event|Event|SIMPLE_SEGMENT|7953,7963|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|7953,7963|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|7953,7963|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Event|Event|SIMPLE_SEGMENT|7971,7979|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7971,7979|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7971,7979|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|7997,8003|false|false|false|||reduce
Event|Event|SIMPLE_SEGMENT|8008,8012|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|8008,8012|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|SIMPLE_SEGMENT|8008,8015|false|false|false|C0035647|Risk|risk of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8016,8026|false|false|false|C1458156|Recurrent Malignant Neoplasm|recurrence
Event|Event|SIMPLE_SEGMENT|8016,8026|false|false|false|||recurrence
Finding|Pathologic Function|SIMPLE_SEGMENT|8016,8026|false|false|false|C2825055|Recurrence (disease attribute)|recurrence
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8016,8026|false|false|false|C0034897|Recurrence|recurrence
Event|Event|SIMPLE_SEGMENT|8039,8049|false|false|false|||discharged
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8055,8058|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|8055,8058|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|8055,8058|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|SIMPLE_SEGMENT|8070,8078|false|false|false|||continue
Drug|Organic Chemical|SIMPLE_SEGMENT|8094,8103|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8094,8103|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|8094,8103|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|8118,8127|false|false|false|||recommend
Finding|Body Substance|SIMPLE_SEGMENT|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Classification|SIMPLE_SEGMENT|8149,8159|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8149,8159|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8160,8164|false|false|false|||PFTs
Finding|Finding|SIMPLE_SEGMENT|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|8177,8186|false|false|false|||suspicion
Finding|Mental Process|SIMPLE_SEGMENT|8177,8186|false|false|false|C0242114|Suspicion|suspicion
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8191,8199|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|8191,8199|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|8191,8199|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|8200,8211|false|false|false|||obstructive
Finding|Functional Concept|SIMPLE_SEGMENT|8200,8211|false|false|false|C0549186|Obstructed|obstructive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8224,8233|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8224,8233|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|8224,8233|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8235,8242|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8235,8242|false|false|false|||disease
Finding|Body Substance|SIMPLE_SEGMENT|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8255,8264|false|false|false|||developed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8276,8280|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|8276,8280|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8276,8280|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|8286,8289|false|false|false|||RVR
Finding|Finding|SIMPLE_SEGMENT|8286,8289|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|8286,8289|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Event|SIMPLE_SEGMENT|8303,8312|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8303,8312|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|8324,8327|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|8324,8327|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|8324,8337|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8324,8337|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8328,8337|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|8328,8337|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|8328,8337|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8328,8337|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8328,8337|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8355,8367|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|8355,8367|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8373,8381|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|8373,8381|false|false|false|||diabetes
Event|Event|SIMPLE_SEGMENT|8383,8398|false|false|false|||Anticoagulation
Finding|Finding|SIMPLE_SEGMENT|8383,8398|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|8383,8398|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8383,8398|false|false|false|C0003281|Anticoagulation Therapy|Anticoagulation
Event|Event|SIMPLE_SEGMENT|8407,8414|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|8428,8437|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8428,8437|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|8456,8460|false|false|false|||felt
Finding|Finding|SIMPLE_SEGMENT|8480,8483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|8480,8483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|8480,8488|false|false|false|C5201228;C5202762|International Prognostic Index Low Risk Group;Low risk|low risk
Event|Event|SIMPLE_SEGMENT|8484,8488|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|8484,8488|false|false|false|C0035647|Risk|risk
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8494,8497|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8494,8497|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|8494,8497|false|false|false|||CVA
Event|Event|SIMPLE_SEGMENT|8514,8518|false|false|false|||make
Event|Event|SIMPLE_SEGMENT|8521,8525|false|false|false|||note
Finding|Finding|SIMPLE_SEGMENT|8534,8537|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|8534,8537|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|8534,8547|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8534,8547|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8538,8547|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|8538,8547|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|8538,8547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8538,8547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8538,8547|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|SIMPLE_SEGMENT|8562,8566|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|8562,8566|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|8562,8570|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|SIMPLE_SEGMENT|8571,8586|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|8571,8586|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|8571,8586|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8571,8586|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|8600,8611|false|false|false|||appropriate
Finding|Idea or Concept|SIMPLE_SEGMENT|8624,8629|false|false|false|C0750546|newly|newly
Event|Event|SIMPLE_SEGMENT|8630,8639|false|false|false|||diagnosed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8649,8654|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8649,8654|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|SIMPLE_SEGMENT|8649,8654|false|false|false|||HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8649,8654|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Event|Event|SIMPLE_SEGMENT|8679,8689|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|8693,8702|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8693,8702|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|8693,8702|false|false|false|||metformin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8707,8710|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8707,8710|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8707,8710|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8707,8710|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8707,8710|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|8717,8724|false|false|false|||require
Finding|Classification|SIMPLE_SEGMENT|8726,8736|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8726,8736|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8737,8743|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|8737,8743|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8737,8743|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8737,8746|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8737,8746|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|8764,8772|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|8785,8787|false|false|false|||in
Finding|Classification|SIMPLE_SEGMENT|8793,8803|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8793,8803|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8804,8811|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|8804,8811|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|8824,8832|false|false|false|||reassess
Event|Event|SIMPLE_SEGMENT|8833,8837|false|false|false|||need
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8842,8850|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|SIMPLE_SEGMENT|8842,8850|false|false|false|||diuretic
Finding|Classification|SIMPLE_SEGMENT|8858,8868|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|8858,8868|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|8869,8876|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|8869,8876|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|8907,8915|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|8907,8915|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|8907,8918|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8919,8924|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8919,8924|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|8919,8924|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8919,8932|true|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|8925,8932|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|8946,8955|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8946,8955|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|8967,8977|false|false|false|||discharged
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8981,8990|false|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|8981,8990|false|false|false|||diuretics
Finding|Finding|SIMPLE_SEGMENT|8994,8997|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|8994,8997|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8994,9009|false|false|false|C1718097|New medications|New medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8998,9009|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8998,9009|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8998,9009|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8998,9009|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9011,9020|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9011,9020|false|false|false|C0025598|metformin|Metformin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9027,9030|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9027,9030|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9027,9030|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9027,9030|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9027,9030|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9031,9041|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9031,9041|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9054,9064|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9054,9064|false|false|false|C0028978|omeprazole|Omeprazole
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9085,9096|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9085,9096|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9085,9096|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9085,9096|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9098,9110|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9098,9110|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|9116,9119|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9120,9130|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9120,9130|false|false|false|C0009262|colchicine|Colchicine
Event|Event|SIMPLE_SEGMENT|9120,9130|false|false|false|||Colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9137,9140|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9137,9140|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9137,9140|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9137,9140|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9137,9140|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9141,9150|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9141,9150|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|SIMPLE_SEGMENT|9157,9160|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Drug|Vitamin|SIMPLE_SEGMENT|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9161,9171|false|false|false|C0523631|Folic acid measurement|Folic acid
Drug|Organic Chemical|SIMPLE_SEGMENT|9182,9192|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9182,9192|false|false|false|C0074393|sertraline|Sertraline
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9214,9225|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9214,9225|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9214,9225|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9214,9225|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9228,9240|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9228,9240|false|false|false|C0025677|methotrexate|Methotrexate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9228,9240|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Drug|Organic Chemical|SIMPLE_SEGMENT|9249,9259|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9249,9259|false|false|false|C0015620|famotidine|Famotidine
Finding|Intellectual Product|SIMPLE_SEGMENT|9269,9274|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|9275,9281|false|false|false|||ISSUES
Finding|Intellectual Product|SIMPLE_SEGMENT|9301,9306|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9301,9319|false|false|false|C0155679|Acute pericarditis|Acute pericarditis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9307,9319|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|9307,9319|false|false|false|||pericarditis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9323,9330|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|9323,9330|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9323,9340|false|false|false|C0007177|Cardiac Tamponade|Cardiac tamponade
Event|Event|SIMPLE_SEGMENT|9331,9340|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|9331,9340|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9331,9340|false|false|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|9350,9368|false|false|false|||pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9350,9368|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Drug|Substance|SIMPLE_SEGMENT|9373,9378|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|9373,9378|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|9373,9378|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|9379,9388|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|9379,9388|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9379,9388|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|9393,9402|false|false|false|||presented
Finding|Functional Concept|SIMPLE_SEGMENT|9408,9420|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9421,9433|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|9421,9433|false|false|false|||pericarditis
Finding|Finding|SIMPLE_SEGMENT|9437,9445|false|false|false|C0332148|Probable diagnosis|probable
Event|Event|SIMPLE_SEGMENT|9446,9451|false|false|false|||viral
Finding|Functional Concept|SIMPLE_SEGMENT|9446,9451|false|true|false|C0521026|Viral|viral
Event|Event|SIMPLE_SEGMENT|9453,9459|false|false|false|||nature
Finding|Functional Concept|SIMPLE_SEGMENT|9453,9459|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|9453,9459|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|SIMPLE_SEGMENT|9467,9474|false|false|false|||context
Finding|Idea or Concept|SIMPLE_SEGMENT|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|SIMPLE_SEGMENT|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|SIMPLE_SEGMENT|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Functional Concept|SIMPLE_SEGMENT|9478,9483|false|false|false|C0521026|Viral|viral
Event|Event|SIMPLE_SEGMENT|9489,9497|false|false|false|||prodrome
Finding|Sign or Symptom|SIMPLE_SEGMENT|9489,9497|false|false|false|C0240805|Prodrome|prodrome
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9505,9514|false|false|false|C0035435|Rheumatism|rheumatic
Event|Event|SIMPLE_SEGMENT|9505,9514|false|false|false|||rheumatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9516,9528|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|9516,9528|false|false|false|||pericarditis
Event|Event|SIMPLE_SEGMENT|9536,9545|false|false|false|||serologic
Finding|Functional Concept|SIMPLE_SEGMENT|9536,9545|false|false|false|C0205473|Serologic|serologic
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|9546,9554|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|SIMPLE_SEGMENT|9546,9554|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|9546,9554|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9562,9569|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|9562,9569|false|false|false|||disease
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|9578,9585|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|SIMPLE_SEGMENT|9578,9585|false|false|false|||absence
Finding|Functional Concept|SIMPLE_SEGMENT|9578,9585|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|SIMPLE_SEGMENT|9578,9588|false|false|false|C0332197|Absent|absence of
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9589,9594|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|SIMPLE_SEGMENT|9589,9594|false|false|false|||DMARD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9596,9607|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9596,9607|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9596,9613|false|false|false|C0031039|Pericardial effusion|Pericardial fluid
Finding|Body Substance|SIMPLE_SEGMENT|9596,9613|false|false|false|C0225973|Pericardial fluid (substance)|Pericardial fluid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9596,9613|false|false|false|C3854061|pericardial fluid analysis|Pericardial fluid
Drug|Substance|SIMPLE_SEGMENT|9608,9613|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|9608,9613|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9608,9613|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|9614,9622|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|9614,9622|false|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|9633,9641|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|9633,9641|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|9633,9641|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9633,9641|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|9643,9651|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|9643,9651|false|false|false|C0010453|Culture (Anthropological)|cultures
Anatomy|Cell|SIMPLE_SEGMENT|9664,9670|false|false|false|C1947989|Colony (cells or organisms)|colony
Event|Event|SIMPLE_SEGMENT|9685,9689|false|false|false|||coag
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9685,9689|false|false|false|C0005790|Blood coagulation tests|coag
Finding|Classification|SIMPLE_SEGMENT|9691,9699|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|9691,9699|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9691,9699|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9700,9705|false|false|false|C0038160|Staphylococcal Infections|staph
Event|Event|SIMPLE_SEGMENT|9700,9705|false|false|false|||staph
Event|Event|SIMPLE_SEGMENT|9706,9710|false|false|false|||felt
Drug|Substance|SIMPLE_SEGMENT|9717,9728|true|false|false|C2827365|Contaminant|contaminant
Event|Event|SIMPLE_SEGMENT|9717,9728|false|false|false|||contaminant
Finding|Classification|SIMPLE_SEGMENT|9730,9738|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|9730,9738|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9730,9738|false|false|false|C5237010|Expression Negative|negative
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9739,9748|false|false|false|C1318720|Acid fast stain|acid fast
Finding|Finding|SIMPLE_SEGMENT|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|SIMPLE_SEGMENT|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|SIMPLE_SEGMENT|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Event|Activity|SIMPLE_SEGMENT|9749,9754|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|SIMPLE_SEGMENT|9749,9754|false|false|false|||smear
Finding|Functional Concept|SIMPLE_SEGMENT|9749,9754|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9749,9754|false|false|false|C0444186|Smear test|smear
Finding|Functional Concept|SIMPLE_SEGMENT|9760,9771|false|false|false|C0205474|Biochemical|biochemical
Event|Event|SIMPLE_SEGMENT|9772,9780|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|9772,9780|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|9772,9783|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Tissue|SIMPLE_SEGMENT|9784,9794|false|false|false|C0027061|Myocardium|myocardial
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9784,9801|true|false|false|C0746730|Myocardial injury|myocardial injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9795,9801|true|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|9795,9801|false|false|false|||injury
Event|Event|SIMPLE_SEGMENT|9805,9814|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9805,9814|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|9817,9825|false|false|false|||unlikely
Finding|Finding|SIMPLE_SEGMENT|9817,9825|false|false|false|C0750558|Unlikely|unlikely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9845,9856|false|false|false|C0027059|Myocarditis|myocarditis
Event|Event|SIMPLE_SEGMENT|9845,9856|false|false|false|||myocarditis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9860,9867|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|9860,9867|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9860,9873|false|true|false|C0741923|Cardiac Events|cardiac event
Event|Event|SIMPLE_SEGMENT|9868,9873|false|false|false|||event
Event|Event|SIMPLE_SEGMENT|9868,9873|false|false|false|C0441471|Event|event
Event|Event|SIMPLE_SEGMENT|9875,9883|false|false|false|||sequelae
Finding|Pathologic Function|SIMPLE_SEGMENT|9875,9883|false|false|false|C0243088;C0543419|Sequela of disorder;sequelae aspects|sequelae
Event|Event|SIMPLE_SEGMENT|9906,9911|false|false|false|||noted
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9920,9924|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Event|Event|SIMPLE_SEGMENT|9920,9924|false|false|false|||SBPs
Drug|Substance|SIMPLE_SEGMENT|9950,9955|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|9950,9955|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9950,9969|false|false|false|C0150238|Fluid resuscitation|fluid resuscitation
Event|Event|SIMPLE_SEGMENT|9956,9969|false|false|false|||resuscitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9956,9969|false|false|false|C0035273|Resuscitation (procedure)|resuscitation
Event|Event|SIMPLE_SEGMENT|9974,9992|false|false|false|||pericardiocentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9974,9992|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Event|Event|SIMPLE_SEGMENT|10000,10007|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|10000,10007|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|10012,10021|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|10012,10021|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10012,10021|false|false|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|10022,10032|false|false|false|||physiology
Finding|Physiologic Function|SIMPLE_SEGMENT|10022,10032|false|false|false|C0031843|physiological aspects|physiology
Event|Event|SIMPLE_SEGMENT|10034,10046|false|false|false|||Hemodynamics
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10034,10046|false|false|false|C0019010|Hemodynamics|Hemodynamics
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10034,10046|false|false|false|C4281788|hemodynamics (procedure)|Hemodynamics
Event|Event|SIMPLE_SEGMENT|10061,10071|false|false|false|||stabilized
Event|Event|SIMPLE_SEGMENT|10076,10084|false|false|false|||remained
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10103,10111|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Event|Event|SIMPLE_SEGMENT|10120,10129|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|10120,10129|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|10136,10139|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10136,10139|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|10147,10153|false|false|false|||showed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10157,10168|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10157,10168|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Event|Event|SIMPLE_SEGMENT|10170,10178|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10180,10191|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10180,10191|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Drug|Substance|SIMPLE_SEGMENT|10192,10197|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|10192,10197|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|10192,10197|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|10212,10216|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|10212,10216|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|10220,10227|false|false|false|||gravity
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10220,10227|false|false|false|C0282189|Gravity (physical force)|gravity
Event|Event|SIMPLE_SEGMENT|10236,10245|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|10246,10252|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|10246,10252|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|10246,10252|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|10262,10269|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|10282,10289|false|false|false|||treated
Drug|Organic Chemical|SIMPLE_SEGMENT|10296,10306|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10296,10306|false|false|false|C0009262|colchicine|colchicine
Event|Event|SIMPLE_SEGMENT|10296,10306|false|false|false|||colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10313,10316|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10313,10316|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10313,10316|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10313,10316|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10313,10316|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|10331,10339|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|10360,10369|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10360,10369|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|SIMPLE_SEGMENT|10388,10397|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10388,10397|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|10388,10397|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|10407,10410|false|false|false|||TID
Event|Event|SIMPLE_SEGMENT|10424,10434|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|10445,10450|false|false|false|||taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|10445,10450|false|false|false|C0441640||taper
Event|Event|SIMPLE_SEGMENT|10455,10463|false|false|false|||received
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10464,10467|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|10464,10467|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|10464,10467|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|SIMPLE_SEGMENT|10474,10483|false|false|false|||receiving
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10485,10491|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDs
Event|Event|SIMPLE_SEGMENT|10485,10491|false|false|false|||NSAIDs
Finding|Intellectual Product|SIMPLE_SEGMENT|10498,10503|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10498,10535|false|false|false|C4040419|Acute Hypercapnic Respiratory Failure|Acute hypercapnic respiratory failure
Finding|Finding|SIMPLE_SEGMENT|10504,10515|false|false|false|C0020440|Hypercapnia|hypercapnic
Finding|Pathologic Function|SIMPLE_SEGMENT|10504,10535|false|false|false|C0398353|Hypercapnic respiratory failure|hypercapnic respiratory failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10516,10527|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10516,10535|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|10528,10535|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|10538,10547|false|false|false|||resolving
Finding|Finding|SIMPLE_SEGMENT|10548,10556|false|false|false|C0332148|Probable diagnosis|Probable
Event|Event|SIMPLE_SEGMENT|10557,10562|false|false|false|||flash
Finding|Gene or Genome|SIMPLE_SEGMENT|10557,10562|false|true|false|C1413133;C4284306|CASP8AP2 gene;CASP8AP2 wt Allele|flash
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10557,10562|false|true|false|C0262485|Flash|flash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10557,10578|false|true|false|C1168329|Flash pulmonary oedema|flash pulmonary edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10563,10572|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10563,10572|false|true|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10563,10572|false|true|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10563,10578|false|true|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10573,10578|false|true|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10573,10578|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10573,10578|false|true|false|C0013604|Edema|edema
Finding|Gene or Genome|SIMPLE_SEGMENT|10590,10595|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|SIMPLE_SEGMENT|10596,10602|false|false|false|C1705102|Volume (publication)|volume
Drug|Substance|SIMPLE_SEGMENT|10603,10608|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|10603,10608|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|10603,10608|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|10610,10624|false|false|false|||administration
Event|Occupational Activity|SIMPLE_SEGMENT|10610,10624|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10610,10624|false|false|false|C1533734|Administration (procedure)|administration
Event|Event|SIMPLE_SEGMENT|10628,10637|false|false|false|||tamponade
Finding|Functional Concept|SIMPLE_SEGMENT|10628,10637|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10628,10637|false|false|false|C0579016||tamponade
Event|Event|SIMPLE_SEGMENT|10642,10651|false|false|false|||evidenced
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10655,10667|false|false|false|C0444708|Radiographic|radiographic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10669,10678|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10669,10678|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10669,10678|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10669,10684|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10679,10684|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10679,10684|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10679,10684|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|10694,10708|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10694,10708|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|10723,10733|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|10723,10733|true|false|false|C0332299|Suggestive of|suggestive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10738,10749|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|SIMPLE_SEGMENT|10738,10761|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10750,10761|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|10750,10761|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|SIMPLE_SEGMENT|10766,10769|false|false|false|||BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|10766,10769|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10766,10769|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|SIMPLE_SEGMENT|10795,10798|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10795,10798|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|10819,10827|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|10819,10827|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|10819,10830|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10831,10838|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|10831,10838|true|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10831,10847|true|false|false|C0741922|CARDIAC ETIOLOGY|cardiac etiology
Event|Event|SIMPLE_SEGMENT|10839,10847|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|10839,10847|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|10839,10847|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10857,10866|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10857,10866|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10857,10866|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10857,10872|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10867,10872|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10867,10872|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10867,10872|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10873,10884|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10873,10892|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|10885,10892|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Body Substance|SIMPLE_SEGMENT|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|10902,10908|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10902,10908|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10939,10948|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10939,10948|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10939,10948|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|10950,10960|false|false|false|||physiology
Finding|Physiologic Function|SIMPLE_SEGMENT|10950,10960|false|false|false|C0031843|physiological aspects|physiology
Finding|Functional Concept|SIMPLE_SEGMENT|10979,10992|true|false|false|C0333159|Emphysematous|emphysematous
Event|Event|SIMPLE_SEGMENT|10993,11000|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|10993,11000|true|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|11001,11006|false|false|false|||noted
Finding|Intellectual Product|SIMPLE_SEGMENT|11018,11022|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|SIMPLE_SEGMENT|11023,11026|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Conceptual Entity|SIMPLE_SEGMENT|11032,11042|false|false|false|C1706907|Background|background
Finding|Functional Concept|SIMPLE_SEGMENT|11043,11054|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11055,11061|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|11055,11061|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|11055,11061|false|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|11065,11076|false|false|false|||conceivable
Event|Event|SIMPLE_SEGMENT|11084,11094|false|false|false|||compelling
Event|Event|SIMPLE_SEGMENT|11095,11102|false|false|false|||smoking
Event|Event|SIMPLE_SEGMENT|11103,11110|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Classification|SIMPLE_SEGMENT|11121,11129|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|11121,11129|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11121,11129|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11130,11133|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|11130,11133|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|11130,11133|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11130,11133|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|SIMPLE_SEGMENT|11138,11142|false|false|false|||week
Finding|Intellectual Product|SIMPLE_SEGMENT|11138,11142|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|11153,11162|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11153,11162|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11176,11188|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|11176,11188|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|11176,11188|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|11192,11201|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11192,11201|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|11210,11215|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|11210,11215|false|false|false|C1550016|Remote control command - Clear|clear
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11217,11229|false|false|false|C0444708|Radiographic|radiographic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11230,11243|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|11230,11243|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|11244,11254|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|11244,11254|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|11244,11257|false|false|false|C0332299|Suggestive of|suggestive of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11258,11267|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|11258,11267|false|false|false|||pneumonia
Drug|Antibiotic|SIMPLE_SEGMENT|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|SIMPLE_SEGMENT|11291,11303|false|false|false|||azithromycin
Event|Event|SIMPLE_SEGMENT|11314,11323|false|false|false|||overnight
Event|Event|SIMPLE_SEGMENT|11328,11340|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|11365,11373|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|11365,11373|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|SIMPLE_SEGMENT|11379,11390|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|11391,11402|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|11391,11402|false|false|false|C2986411|Improvement|improvement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11411,11422|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11411,11429|false|false|false|C2598168||respiratory status
Finding|Finding|SIMPLE_SEGMENT|11411,11429|false|false|false|C1998827|Respiratory Status|respiratory status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11423,11429|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|11423,11429|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|11423,11429|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|11461,11470|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|11505,11514|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11505,11514|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|11520,11530|false|false|false|||ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|11520,11530|false|false|false|C1561560|ambulatory encounter|ambulatory
Event|Event|SIMPLE_SEGMENT|11532,11543|false|false|false|||saturations
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11532,11543|false|false|false|C0522534|Saturated|saturations
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11566,11570|false|false|false|C0004238|Atrial Fibrillation|AFib
Event|Event|SIMPLE_SEGMENT|11566,11570|false|false|false|||AFib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11566,11570|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Finding|Finding|SIMPLE_SEGMENT|11572,11575|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|11572,11575|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|11572,11585|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11572,11585|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11576,11585|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|11576,11585|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|11576,11585|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|11576,11585|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11576,11585|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Body Substance|SIMPLE_SEGMENT|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|11595,11599|false|false|false|||went
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11605,11609|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11605,11609|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|SIMPLE_SEGMENT|11615,11618|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|SIMPLE_SEGMENT|11615,11618|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Drug|Organic Chemical|SIMPLE_SEGMENT|11654,11664|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11654,11664|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|11654,11664|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|11682,11689|false|false|false|||flipped
Event|Event|SIMPLE_SEGMENT|11700,11703|false|false|false|||NSR
Finding|Molecular Function|SIMPLE_SEGMENT|11700,11703|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|SIMPLE_SEGMENT|11700,11703|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Event|Event|SIMPLE_SEGMENT|11710,11719|false|false|false|||CHADsVASC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11729,11732|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|11729,11732|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|11735,11750|false|false|false|||Anticoagulation
Finding|Finding|SIMPLE_SEGMENT|11735,11750|false|false|true|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|11735,11750|false|false|true|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11735,11750|false|false|true|C0003281|Anticoagulation Therapy|Anticoagulation
Event|Event|SIMPLE_SEGMENT|11755,11764|false|false|false|||discussed
Event|Event|SIMPLE_SEGMENT|11781,11789|false|false|false|||deferred
Finding|Finding|SIMPLE_SEGMENT|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|11805,11814|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11805,11814|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|11815,11820|false|false|false|||given
Finding|Body Substance|SIMPLE_SEGMENT|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11836,11841|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|11836,11841|false|false|false|C2003888|Lower (action)|lower
Finding|Intellectual Product|SIMPLE_SEGMENT|11842,11849|false|false|false|C0282416|Overall Publication Type|overall
Event|Event|SIMPLE_SEGMENT|11850,11854|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|11850,11854|false|false|false|C0035647|Risk|risk
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11859,11862|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11859,11862|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|11859,11862|false|false|false|||CVA
Event|Event|SIMPLE_SEGMENT|11867,11875|false|false|false|||concerns
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11886,11896|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|11886,11896|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11886,11896|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|11898,11907|false|false|false|||adherence
Finding|Functional Concept|SIMPLE_SEGMENT|11898,11907|false|false|false|C1510802|Adherence (attribute)|adherence
Event|Event|SIMPLE_SEGMENT|11908,11912|false|false|false|||cost
Finding|Functional Concept|SIMPLE_SEGMENT|11908,11912|false|false|false|C0220812;C4050363|Comprehensive Score for Financial Toxicity;Cost aspects|cost
Finding|Intellectual Product|SIMPLE_SEGMENT|11908,11912|false|false|false|C0220812;C4050363|Comprehensive Score for Financial Toxicity;Cost aspects|cost
Event|Event|SIMPLE_SEGMENT|11921,11931|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|11935,11945|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11935,11945|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|11935,11945|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|11967,11971|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|11967,11971|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|11967,11975|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|SIMPLE_SEGMENT|11976,11991|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|11976,11991|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|11976,11991|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11976,11991|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|11992,12002|false|false|false|||reassessed
Event|Event|SIMPLE_SEGMENT|12009,12019|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|12009,12019|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|12009,12019|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|12034,12045|false|false|false|||appropriate
Finding|Gene or Genome|SIMPLE_SEGMENT|12052,12056|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|12052,12056|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12052,12068|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12060,12068|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|12060,12068|false|false|false|||diabetes
Finding|Idea or Concept|SIMPLE_SEGMENT|12078,12083|false|false|false|C0750546|newly|newly
Event|Event|SIMPLE_SEGMENT|12084,12093|false|false|false|||diagnosed
Event|Event|SIMPLE_SEGMENT|12109,12112|false|false|false|||A1C
Finding|Classification|SIMPLE_SEGMENT|12109,12112|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12109,12112|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Event|Event|SIMPLE_SEGMENT|12134,12143|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12134,12143|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|12152,12162|false|false|false|||maintained
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|12169,12176|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|12169,12176|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12169,12176|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|12177,12184|false|false|false|||sliding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12185,12190|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|12185,12190|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|12185,12190|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|12185,12190|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|12191,12197|false|false|false|||during
Event|Event|SIMPLE_SEGMENT|12204,12213|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12204,12213|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|12226,12236|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|12240,12249|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12240,12249|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|12250,12255|false|false|false|||500mg
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12256,12259|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12256,12259|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12256,12259|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12256,12259|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12256,12259|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|12263,12270|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|12263,12270|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|12263,12270|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|12271,12277|false|false|false|C1547311|Patient Condition Code - Stable|STABLE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12310,12330|false|false|false|C0003873|Rheumatoid Arthritis|Rheumatoid arthritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12321,12330|false|false|false|C0003864|Arthritis|arthritis
Event|Event|SIMPLE_SEGMENT|12321,12330|false|false|false|||arthritis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12340,12348|false|false|false|C4318437|Anti-Cyclic Citrullinated Protein Antibodies|anti-CCP
Drug|Immunologic Factor|SIMPLE_SEGMENT|12340,12348|false|false|false|C4318437|Anti-Cyclic Citrullinated Protein Antibodies|anti-CCP
Event|Event|SIMPLE_SEGMENT|12340,12348|false|false|false|||anti-CCP
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|12349,12357|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|12349,12357|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|12349,12357|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|12349,12357|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Classification|SIMPLE_SEGMENT|12362,12372|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|12362,12372|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|12373,12385|false|false|false|||rheumatology
Event|Event|SIMPLE_SEGMENT|12414,12424|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|12414,12424|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|12414,12427|false|false|false|C0332299|Suggestive of|suggestive of
Event|Event|SIMPLE_SEGMENT|12431,12436|false|false|false|||flare
Finding|Finding|SIMPLE_SEGMENT|12431,12436|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|SIMPLE_SEGMENT|12431,12436|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|SIMPLE_SEGMENT|12442,12452|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|12442,12452|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12442,12452|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|SIMPLE_SEGMENT|12461,12475|false|false|false|||rheumatologist
Event|Event|SIMPLE_SEGMENT|12477,12485|false|false|false|||deferred
Event|Event|SIMPLE_SEGMENT|12486,12496|false|false|false|||restarting
Drug|Organic Chemical|SIMPLE_SEGMENT|12497,12500|false|false|false|C0025677|methotrexate|MTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12497,12500|false|false|false|C0025677|methotrexate|MTX
Event|Event|SIMPLE_SEGMENT|12497,12500|false|false|false|||MTX
Finding|Gene or Genome|SIMPLE_SEGMENT|12497,12500|false|false|false|C1417487;C5891182|MTX1 gene;Matrix Market File Format|MTX
Finding|Intellectual Product|SIMPLE_SEGMENT|12497,12500|false|false|false|C1417487;C5891182|MTX1 gene;Matrix Market File Format|MTX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12514,12519|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|SIMPLE_SEGMENT|12514,12519|false|false|false|||DMARD
Event|Event|SIMPLE_SEGMENT|12526,12536|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|12526,12536|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|12526,12536|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12542,12545|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|12542,12545|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|12550,12554|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|12550,12554|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12550,12554|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12550,12554|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12558,12562|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|SIMPLE_SEGMENT|12558,12562|false|false|false|||meds
Finding|Intellectual Product|SIMPLE_SEGMENT|12558,12562|false|false|false|C4284232|Medications|meds
Event|Event|SIMPLE_SEGMENT|12568,12572|false|false|false|||held
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12590,12594|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12595,12598|false|false|false|C1849718|POPLITEAL PTERYGIUM SYNDROME, LETHAL TYPE|BPs
Drug|Organic Chemical|SIMPLE_SEGMENT|12595,12598|false|false|false|C2740858|BPS|BPs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12595,12598|false|false|false|C2740858|BPS|BPs
Event|Event|SIMPLE_SEGMENT|12595,12598|false|false|false|||BPs
Event|Event|SIMPLE_SEGMENT|12609,12616|false|false|false|||stopped
Finding|Finding|SIMPLE_SEGMENT|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|12632,12641|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12632,12641|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|12648,12656|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|12657,12669|false|false|false|||normotensive
Anatomy|Cell Component|SIMPLE_SEGMENT|12673,12677|false|false|false|C1167518|viral nucleocapsid location|CORE
Finding|Body Substance|SIMPLE_SEGMENT|12673,12677|false|false|false|C3274653|Core Specimen|CORE
Event|Event|SIMPLE_SEGMENT|12678,12686|false|false|false|||MEASURES
Finding|Functional Concept|SIMPLE_SEGMENT|12678,12686|false|false|false|C1879489|Measures (attribute)|MEASURES
Event|Event|SIMPLE_SEGMENT|12706,12710|false|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|12706,12710|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|12706,12710|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12712,12715|false|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|12712,12715|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|12712,12715|false|false|false|C0011015|daunorubicin|DNR
Event|Event|SIMPLE_SEGMENT|12712,12715|false|false|false|||DNR
Finding|Finding|SIMPLE_SEGMENT|12712,12715|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|12712,12715|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Activity|SIMPLE_SEGMENT|12722,12729|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|12722,12729|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|12722,12729|false|false|false|C0392367|Physical contact|CONTACT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12730,12733|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|12730,12733|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|12730,12733|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12757,12768|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12757,12768|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|12757,12768|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12757,12768|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|12757,12781|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|12772,12781|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12772,12781|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12800,12810|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12800,12810|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12800,12815|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|12811,12815|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|12811,12815|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|12819,12827|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|12832,12840|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|12832,12840|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|12832,12840|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|12845,12857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12845,12857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12875,12885|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12875,12885|false|false|false|C0009262|colchicine|Colchicine
Event|Event|SIMPLE_SEGMENT|12875,12885|false|false|false|||Colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12896,12899|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12896,12899|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12896,12899|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12896,12899|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12896,12899|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12904,12913|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12904,12913|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|SIMPLE_SEGMENT|12924,12927|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|12932,12942|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12932,12942|false|false|false|C0015620|famotidine|Famotidine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12962,12972|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12962,12972|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|12962,12972|false|false|false|||lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12962,12992|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|12973,12992|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12973,12992|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|SIMPLE_SEGMENT|12973,12992|false|false|false|||hydrochlorothiazide
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13000,13004|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13000,13004|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|13000,13004|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|13000,13004|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|13005,13010|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|13015,13027|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13015,13027|false|false|false|C0025677|methotrexate|Methotrexate
Event|Event|SIMPLE_SEGMENT|13015,13027|false|false|false|||Methotrexate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13015,13027|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Finding|Intellectual Product|SIMPLE_SEGMENT|13040,13044|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Organic Chemical|SIMPLE_SEGMENT|13055,13065|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13055,13065|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Vitamin|SIMPLE_SEGMENT|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13086,13096|false|false|false|C0523631|Folic acid measurement|FoLIC Acid
Event|Event|SIMPLE_SEGMENT|13092,13096|false|false|false|||Acid
Event|Event|SIMPLE_SEGMENT|13115,13124|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13115,13124|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|13115,13136|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13125,13136|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13125,13136|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|13125,13136|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13125,13136|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|13142,13151|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13142,13151|false|false|false|C0001927|albuterol|Albuterol
Event|Event|SIMPLE_SEGMENT|13152,13159|false|false|false|||Inhaler
Finding|Functional Concept|SIMPLE_SEGMENT|13152,13159|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|13174,13177|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|13178,13186|false|false|false|||wheezing
Event|Event|SIMPLE_SEGMENT|13188,13197|false|false|false|||shortness
Finding|Body Substance|SIMPLE_SEGMENT|13202,13208|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|13214,13223|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13214,13223|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|13214,13231|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13214,13231|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|13224,13231|false|false|false|||sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|13233,13239|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13233,13239|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|SIMPLE_SEGMENT|13233,13243|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13233,13243|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13240,13243|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|SIMPLE_SEGMENT|13240,13243|false|false|false|||HFA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13240,13243|false|false|false|C0430649|High frequency audiometry|HFA
Event|Event|SIMPLE_SEGMENT|13281,13287|false|false|false|||needed
Finding|Functional Concept|SIMPLE_SEGMENT|13297,13304|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Event|Event|SIMPLE_SEGMENT|13305,13312|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13305,13312|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13321,13330|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13321,13330|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|SIMPLE_SEGMENT|13332,13342|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13332,13342|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13354,13357|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13354,13357|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13354,13357|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13354,13357|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13354,13357|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13363,13372|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13363,13372|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|13363,13372|false|false|false|||metformin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13382,13388|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|13392,13400|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13395,13400|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13395,13400|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|13409,13412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|13409,13412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13424,13430|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13431,13438|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13431,13438|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13447,13457|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13447,13457|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|13447,13467|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13447,13467|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|13458,13467|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|13491,13501|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13491,13501|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|13491,13511|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13491,13511|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|13502,13511|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|SIMPLE_SEGMENT|13502,13511|false|false|false|||succinate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13520,13526|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|13530,13538|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13533,13538|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13533,13538|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|13545,13549|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|13545,13549|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13556,13562|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13563,13570|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13563,13570|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13579,13589|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13579,13589|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|13610,13620|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13610,13620|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|SIMPLE_SEGMENT|13610,13620|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13629,13636|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|13629,13636|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13629,13636|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|13640,13648|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13643,13648|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13643,13648|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13666,13673|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|13666,13673|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13666,13673|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|13674,13681|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13674,13681|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13690,13702|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13690,13702|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|13722,13732|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13722,13732|false|false|false|C0009262|colchicine|Colchicine
Event|Event|SIMPLE_SEGMENT|13722,13732|false|false|false|||Colchicine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13743,13746|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13743,13746|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13743,13746|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13743,13746|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13743,13746|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13752,13762|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13752,13762|false|false|false|C0009262|colchicine|colchicine
Event|Event|SIMPLE_SEGMENT|13752,13762|false|false|false|||colchicine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13772,13779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|13772,13779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13772,13779|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|13783,13791|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13786,13791|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13786,13791|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|13800,13803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|13800,13803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|13804,13808|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|13804,13808|false|false|false|C2828567|PRSS30P gene|Disp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13815,13822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|13815,13822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13815,13822|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|13823,13830|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|13823,13830|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Vitamin|SIMPLE_SEGMENT|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13839,13849|false|false|false|C0523631|Folic acid measurement|FoLIC Acid
Event|Event|SIMPLE_SEGMENT|13845,13849|false|false|false|||Acid
Drug|Organic Chemical|SIMPLE_SEGMENT|13870,13879|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13870,13879|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|SIMPLE_SEGMENT|13890,13893|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|13900,13910|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13900,13910|false|false|false|C0074393|sertraline|Sertraline
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13933,13937|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13933,13937|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|13933,13937|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|13933,13937|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|13933,13937|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13939,13949|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13939,13949|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|13939,13949|false|false|false|||lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13939,13969|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|13950,13969|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13950,13969|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|SIMPLE_SEGMENT|13950,13969|false|false|false|||hydrochlorothiazide
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13977,13981|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13977,13981|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|13977,13981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|13977,13981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|13982,13987|false|false|false|||DAILY
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13995,14005|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|13995,14005|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13995,14005|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|14010,14014|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|14023,14030|false|false|false|||restart
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14032,14042|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14032,14042|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|14032,14042|false|false|false|||lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14032,14062|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|14043,14062|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14043,14062|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|SIMPLE_SEGMENT|14043,14062|false|false|false|||hydrochlorothiazide
Event|Event|SIMPLE_SEGMENT|14069,14079|false|false|false|||instructed
Event|Activity|SIMPLE_SEGMENT|14097,14101|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|14097,14101|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14097,14101|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|14102,14108|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|14102,14108|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|14112,14124|false|false|false|||cardiologist
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14129,14133|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14129,14133|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|14129,14133|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|14129,14133|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|14129,14133|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|SIMPLE_SEGMENT|14135,14147|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14135,14147|false|false|false|C0025677|methotrexate|Methotrexate
Event|Event|SIMPLE_SEGMENT|14135,14147|false|false|false|||Methotrexate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14135,14147|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Finding|Intellectual Product|SIMPLE_SEGMENT|14160,14164|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14177,14187|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|14177,14187|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|14177,14187|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|14193,14197|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|14206,14213|false|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|14214,14226|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14214,14226|false|false|false|C0025677|methotrexate|Methotrexate
Event|Event|SIMPLE_SEGMENT|14214,14226|false|false|false|||Methotrexate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14214,14226|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Event|Event|SIMPLE_SEGMENT|14235,14241|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|14235,14241|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|14259,14268|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14259,14268|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14259,14280|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|14259,14280|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14269,14280|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|14269,14280|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|14269,14280|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|14282,14286|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|14282,14286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|14282,14286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|14282,14286|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|14289,14298|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14289,14298|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14289,14308|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14299,14308|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14299,14308|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14299,14308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14299,14308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14299,14308|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14310,14327|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14318,14327|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14318,14327|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14318,14327|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14318,14327|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14318,14327|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14329,14341|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14342,14354|false|false|false|C0031046|Pericarditis|pericarditis
Event|Event|SIMPLE_SEGMENT|14342,14354|false|false|false|||pericarditis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14355,14364|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|14355,14364|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|14355,14364|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14355,14374|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|SIMPLE_SEGMENT|14355,14374|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14365,14374|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|14365,14374|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|14365,14374|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|14365,14374|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14365,14374|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14376,14396|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14387,14396|false|false|false|C0003864|Arthritis|arthritis
Event|Event|SIMPLE_SEGMENT|14387,14396|false|false|false|||arthritis
Event|Event|SIMPLE_SEGMENT|14401,14410|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14401,14410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14401,14410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14401,14410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14401,14410|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14411,14420|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14411,14420|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|14411,14420|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|14411,14420|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|14422,14428|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14422,14435|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|14422,14435|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14429,14435|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14429,14435|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|14437,14442|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|14437,14442|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|14447,14455|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|14447,14455|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|14457,14462|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14457,14479|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|14457,14479|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|14466,14479|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|14466,14479|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|14466,14479|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14481,14486|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|14481,14486|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14481,14486|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|14481,14486|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|14491,14502|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|14491,14502|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|14504,14512|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|14504,14512|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|14504,14512|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14513,14519|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|14513,14519|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|14513,14519|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|14521,14531|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|14521,14531|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|14534,14545|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|14534,14545|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|14534,14545|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|14550,14559|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14550,14559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14550,14559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14550,14559|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14550,14559|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14550,14572|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14550,14572|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|14550,14572|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14560,14572|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14560,14572|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14560,14572|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|14574,14578|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|14592,14595|false|false|false|||WHY
Event|Event|SIMPLE_SEGMENT|14596,14600|false|false|false|||WERE
Event|Event|SIMPLE_SEGMENT|14605,14613|false|false|false|||ADMITTED
Event|Event|SIMPLE_SEGMENT|14621,14629|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|14621,14629|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|14644,14652|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|14660,14668|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14674,14679|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|14674,14679|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14674,14684|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|14674,14684|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14680,14684|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|14680,14684|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|14680,14684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|14680,14684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|14694,14697|false|false|false|||WAS
Event|Event|SIMPLE_SEGMENT|14709,14712|false|false|false|||YOU
Event|Event|SIMPLE_SEGMENT|14713,14717|false|false|false|||WERE
Finding|Idea or Concept|SIMPLE_SEGMENT|14725,14733|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|14749,14754|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|14763,14775|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|14763,14775|false|false|false|C0021368|Inflammation|inflammation
Finding|Conceptual Entity|SIMPLE_SEGMENT|14782,14787|false|false|false|C1707059|Pre-Release Version|build
Event|Event|SIMPLE_SEGMENT|14788,14790|false|false|false|||up
Drug|Substance|SIMPLE_SEGMENT|14794,14799|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|14794,14799|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|14794,14799|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14822,14827|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14822,14827|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|14822,14827|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14841,14850|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|14841,14850|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|14841,14850|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|14841,14850|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14841,14850|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|SIMPLE_SEGMENT|14854,14860|false|false|false|||remove
Drug|Substance|SIMPLE_SEGMENT|14865,14870|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|14865,14870|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|14865,14870|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14895,14900|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14895,14900|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|14895,14900|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|14895,14900|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Idea or Concept|SIMPLE_SEGMENT|14907,14916|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Finding|Intellectual Product|SIMPLE_SEGMENT|14907,14916|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Drug|Substance|SIMPLE_SEGMENT|14917,14922|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|SIMPLE_SEGMENT|14917,14922|false|false|false|||drain
Finding|Intellectual Product|SIMPLE_SEGMENT|14917,14922|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|SIMPLE_SEGMENT|14923,14929|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|14940,14947|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|14960,14964|false|false|false|||left
Event|Event|SIMPLE_SEGMENT|14969,14977|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|14969,14977|false|false|false|C1547192|Organization unit type - Hospital|hospital
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14995,15005|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|14995,15005|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|14995,15005|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|15009,15013|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|15018,15021|false|false|false|||pee
Finding|Pathologic Function|SIMPLE_SEGMENT|15030,15042|false|false|false|C0013604;C0546817|Edema;Hypervolemia (finding)|excess fluid
Drug|Substance|SIMPLE_SEGMENT|15037,15042|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|15037,15042|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|15037,15042|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|15052,15056|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15052,15056|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|15052,15056|false|false|false|C1551342|Document Body|body
Event|Event|SIMPLE_SEGMENT|15065,15074|false|false|false|||developed
Finding|Finding|SIMPLE_SEGMENT|15078,15086|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|15078,15086|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15087,15092|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|15087,15092|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|15087,15092|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|15087,15099|false|false|false|C0232187|Cardiac rhythm type|heart rhythm
Event|Event|SIMPLE_SEGMENT|15093,15099|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|15093,15099|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|15093,15099|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15101,15105|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|15101,15105|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|15101,15105|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|SIMPLE_SEGMENT|15121,15129|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|15121,15129|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|15140,15147|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|15153,15156|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|15153,15156|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15157,15167|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|15157,15167|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|15157,15167|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|SIMPLE_SEGMENT|15179,15189|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15179,15189|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|15203,15212|false|false|false|||diagnosed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15218,15226|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|15218,15226|false|false|false|||diabetes
Event|Event|SIMPLE_SEGMENT|15239,15248|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|15239,15248|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|15260,15267|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|15273,15276|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|15273,15276|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15277,15287|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|15277,15287|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|15277,15287|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|SIMPLE_SEGMENT|15298,15307|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15298,15307|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|15298,15307|false|false|false|||metformin
Event|Event|SIMPLE_SEGMENT|15321,15324|false|false|false|||YOU
Event|Event|SIMPLE_SEGMENT|15325,15329|false|false|false|||NEED
Finding|Functional Concept|SIMPLE_SEGMENT|15325,15329|false|false|false|C0686904|Patient need for (contextual qualifier)|NEED
Event|Event|SIMPLE_SEGMENT|15333,15335|false|false|false|||DO
Event|Event|SIMPLE_SEGMENT|15345,15350|false|false|false|||LEAVE
Event|Event|SIMPLE_SEGMENT|15355,15363|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|15355,15363|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|15369,15373|false|false|false|||Take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15386,15397|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15386,15397|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|15386,15397|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|15386,15397|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|15401,15411|false|false|false|||prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|15431,15437|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|SIMPLE_SEGMENT|15431,15437|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|SIMPLE_SEGMENT|15431,15440|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|15431,15440|false|false|false|C1522577|follow-up|Follow up
Event|Event|SIMPLE_SEGMENT|15438,15440|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|15509,15513|false|false|false|||seek
Finding|Functional Concept|SIMPLE_SEGMENT|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|15514,15521|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|15522,15531|false|false|false|||attention
Finding|Intellectual Product|SIMPLE_SEGMENT|15522,15531|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|15522,15531|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15541,15547|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|15541,15547|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|15541,15547|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|15541,15547|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|15541,15547|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|15548,15552|false|false|false|||goes
Event|Event|SIMPLE_SEGMENT|15568,15571|false|false|false|||lbs
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15568,15571|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Intellectual Product|SIMPLE_SEGMENT|15577,15581|false|false|false|C5239649|PANEL.SURVEY.SEEK|Seek
Finding|Functional Concept|SIMPLE_SEGMENT|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|15582,15589|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|15590,15599|false|false|false|||attention
Finding|Intellectual Product|SIMPLE_SEGMENT|15590,15599|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|15590,15599|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Finding|SIMPLE_SEGMENT|15612,15615|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|15612,15615|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|15630,15638|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|15630,15638|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|15630,15638|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|15655,15663|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|15655,15663|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|15655,15663|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15672,15676|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15672,15676|false|false|false|C5781420||legs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|15678,15687|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|15678,15698|false|false|false|C0000731|Abdomen distended|abdominal distention
Event|Event|SIMPLE_SEGMENT|15688,15698|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|15688,15698|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|15688,15698|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Event|Event|SIMPLE_SEGMENT|15704,15713|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15704,15723|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|15704,15723|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|SIMPLE_SEGMENT|15717,15723|false|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|15717,15723|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|15744,15747|false|false|false|||see
Finding|Idea or Concept|SIMPLE_SEGMENT|15763,15774|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Finding|Intellectual Product|SIMPLE_SEGMENT|15763,15774|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Event|Event|SIMPLE_SEGMENT|15783,15798|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|15783,15798|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|15810,15818|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|15810,15818|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|15810,15818|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|SIMPLE_SEGMENT|15826,15830|false|false|false|||part
Finding|Idea or Concept|SIMPLE_SEGMENT|15826,15830|false|false|false|C1552020|Role Class - part|part
Event|Activity|SIMPLE_SEGMENT|15839,15843|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|15839,15843|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|15839,15843|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|15839,15843|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15880,15884|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|15880,15884|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|15880,15884|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|SIMPLE_SEGMENT|15900,15904|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|15900,15904|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|15900,15904|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15900,15909|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|15900,15909|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|15914,15922|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15923,15935|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|15923,15935|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|15923,15935|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

