 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Chief|276,281
Complaint|282,291
:|291,292
<EOL>|292,293
Shortness|293,302
of|303,305
breath|306,312
<EOL>|312,313
<EOL>|314,315
Major|315,320
Surgical|321,329
or|330,332
Invasive|333,341
Procedure|342,351
:|351,352
<EOL>|352,353
None|353,357
<EOL>|357,358
<EOL>|358,359
<EOL>|360,361
History|361,368
of|369,371
Present|372,379
Illness|380,387
:|387,388
<EOL>|388,389
Ms.|389,392
_|393,394
_|394,395
_|395,396
is|397,399
a|400,401
_|402,403
_|403,404
_|404,405
with|406,410
hx|411,413
COPD|414,418
on|419,421
home|422,426
O2|427,429
,|429,430
atrial|431,437
<EOL>|438,439
fibrillation|439,451
on|452,454
apixaban|455,463
,|463,464
hypertension|465,477
,|477,478
CAD|479,482
,|482,483
and|484,487
hyperlipidemia|488,502
,|502,503
<EOL>|504,505
with|505,509
recurrent|510,519
hospitalizations|520,536
for|537,540
COPD|541,545
exacerbations|546,559
,|559,560
who|561,564
<EOL>|565,566
presented|566,575
with|576,580
dyspnea|581,588
.|588,589
<EOL>|589,590
<EOL>|592,593
She|593,596
has|597,600
had|601,604
multiple|605,613
prior|614,619
admissions|620,630
for|631,634
dyspnea|635,642
.|642,643
She|644,647
was|648,651
<EOL>|652,653
recently|653,661
discharged|662,672
on|673,675
_|676,677
_|677,678
_|678,679
after|680,685
3|686,687
day|688,691
inpatient|692,701
admission|702,711
for|712,715
<EOL>|716,717
COPD|717,721
exacerbation|722,734
.|734,735
She|736,739
was|740,743
discharged|744,754
on|755,757
extended|758,766
prednisone|767,777
<EOL>|778,779
taper|779,784
with|785,789
plan|790,794
for|795,798
5d|799,801
40mg|802,806
Prednisone|807,817
(|818,819
to|819,821
finish|822,828
_|829,830
_|830,831
_|831,832
followed|833,841
<EOL>|842,843
by|843,845
10mg|846,850
taper|851,856
every|857,862
5|863,864
days|865,869
(|870,871
35mg|871,875
from|876,880
_|881,882
_|882,883
_|883,884
,|884,885
30mg|886,890
_|891,892
_|892,893
_|893,894
,|894,895
<EOL>|896,897
etc|897,900
...|900,903
)|903,904
.|904,905
<EOL>|906,907
<EOL>|907,908
On|908,910
the|911,914
evening|915,922
prior|923,928
to|929,931
presentation|932,944
,|944,945
patient|946,953
experienced|954,965
<EOL>|966,967
worsening|967,976
shortness|977,986
of|987,989
breath|990,996
,|996,997
nonproductive|998,1011
cough|1012,1017
and|1018,1021
wheezing|1022,1030
<EOL>|1031,1032
c|1032,1033
/|1033,1034
w|1034,1035
prior|1036,1041
COPD|1042,1046
exacerbations|1047,1060
.|1060,1061
She|1062,1065
reported|1066,1074
taking|1075,1081
inhalers|1082,1090
as|1091,1093
<EOL>|1094,1095
directed|1095,1103
,|1103,1104
without|1105,1112
relief|1113,1119
.|1119,1120
The|1121,1124
patient|1125,1132
reported|1133,1141
that|1142,1146
this|1147,1151
is|1152,1154
<EOL>|1155,1156
almost|1156,1162
identical|1163,1172
to|1173,1175
her|1176,1179
last|1180,1184
presentation|1185,1197
.|1197,1198
She|1199,1202
also|1203,1207
felt|1208,1212
that|1213,1217
<EOL>|1218,1219
she|1219,1222
was|1223,1226
taking|1227,1233
too|1234,1237
many|1238,1242
medications|1243,1254
and|1255,1258
does|1259,1263
not|1264,1267
wish|1268,1272
to|1273,1275
<EOL>|1276,1277
continue|1277,1285
to|1286,1288
take|1289,1293
prednisone|1294,1304
.|1304,1305
The|1306,1309
patient|1310,1317
was|1318,1321
also|1322,1326
noted|1327,1332
to|1333,1335
have|1336,1340
<EOL>|1341,1342
increased|1342,1351
O2|1352,1354
requirement|1355,1366
and|1367,1370
she|1371,1374
was|1375,1378
referred|1379,1387
to|1388,1390
the|1391,1394
_|1395,1396
_|1396,1397
_|1397,1398
ED|1399,1401
<EOL>|1402,1403
for|1403,1406
further|1407,1414
management|1415,1425
.|1425,1426
Of|1427,1429
note|1430,1434
,|1434,1435
please|1436,1442
see|1443,1446
prior|1447,1452
admission|1453,1462
note|1463,1467
<EOL>|1468,1469
for|1469,1472
details|1473,1480
regarding|1481,1490
prior|1491,1496
admission|1497,1506
.|1506,1507
<EOL>|1509,1510
<EOL>|1511,1512
In|1512,1514
the|1515,1518
ED|1519,1521
,|1521,1522
initial|1523,1530
vital|1531,1536
signs|1537,1542
were|1543,1547
:|1547,1548
88|1549,1551
143|1552,1555
/|1555,1556
105|1556,1559
26|1560,1562
94|1563,1565
%|1565,1566
RA|1567,1569
.|1569,1570
Labs|1571,1575
<EOL>|1576,1577
were|1577,1581
notable|1582,1589
for|1590,1593
normal|1594,1600
BNP|1601,1604
and|1605,1608
a|1609,1610
creatinine|1611,1621
of|1622,1624
1.2|1625,1628
.|1628,1629
Patient|1630,1637
was|1638,1641
<EOL>|1642,1643
given|1643,1648
azithromycin|1649,1661
and|1662,1665
duoneb|1666,1672
.|1672,1673
Patient|1674,1681
was|1682,1685
scheduled|1686,1695
to|1696,1698
have|1699,1703
<EOL>|1704,1705
methylpred|1705,1715
but|1716,1719
did|1720,1723
not|1724,1727
have|1728,1732
it|1733,1735
administered|1736,1748
until|1749,1754
arrival|1755,1762
to|1763,1765
the|1766,1769
<EOL>|1770,1771
floor|1771,1776
.|1776,1777
<EOL>|1779,1780
Upon|1781,1785
arrival|1786,1793
to|1794,1796
the|1797,1800
floor|1801,1806
,|1806,1807
she|1808,1811
complained|1812,1822
of|1823,1825
wheezing|1826,1834
and|1835,1838
SOB|1839,1842
.|1842,1843
<EOL>|1844,1845
She|1845,1848
otherwise|1849,1858
felt|1859,1863
well|1864,1868
.|1868,1869
She|1870,1873
agreed|1874,1880
to|1881,1883
take|1884,1888
the|1889,1892
methyprednisone|1893,1908
<EOL>|1909,1910
but|1910,1913
does|1914,1918
not|1919,1922
wish|1923,1927
to|1928,1930
take|1931,1935
prednisone|1936,1946
any|1947,1950
more|1951,1955
.|1955,1956
<EOL>|1958,1959
<EOL>|1960,1961
REVIEW|1961,1967
OF|1968,1970
SYSTEMS|1971,1978
:|1978,1979
Per|1980,1983
HPI|1984,1987
.|1987,1988
Denies|1989,1995
headache|1996,2004
,|2004,2005
visual|2006,2012
changes|2013,2020
,|2020,2021
<EOL>|2022,2023
pharyngitis|2023,2034
,|2034,2035
fevers|2036,2042
,|2042,2043
chills|2044,2050
,|2050,2051
sweats|2052,2058
,|2058,2059
weight|2060,2066
loss|2067,2071
,|2071,2072
chest|2073,2078
pain|2079,2083
,|2083,2084
<EOL>|2085,2086
abdominal|2086,2095
pain|2096,2100
,|2100,2101
nausea|2102,2108
,|2108,2109
vomiting|2110,2118
,|2118,2119
diarrhea|2120,2128
,|2128,2129
constipation|2130,2142
,|2142,2143
<EOL>|2144,2145
hematochezia|2145,2157
,|2157,2158
dysuria|2159,2166
,|2166,2167
rash|2168,2172
,|2172,2173
paresthesias|2174,2186
,|2186,2187
and|2188,2191
weakness|2192,2200
.|2200,2201
<EOL>|2201,2202
<EOL>|2203,2204
Past|2204,2208
Medical|2209,2216
History|2217,2224
:|2224,2225
<EOL>|2225,2226
-|2226,2227
COPD|2228,2232
/|2232,2233
Asthma|2233,2239
on|2240,2242
home|2243,2247
2L|2248,2250
O2|2251,2253
<EOL>|2253,2254
-|2254,2255
Atypical|2256,2264
Chest|2265,2270
Pain|2271,2275
<EOL>|2275,2276
-|2276,2277
Hypertension|2278,2290
<EOL>|2290,2291
-|2291,2292
Hyperlipidemia|2293,2307
<EOL>|2307,2308
-|2308,2309
Osteroarthritis|2310,2325
<EOL>|2325,2326
-|2326,2327
Atrial|2328,2334
Fibrillation|2335,2347
on|2348,2350
Apixaban|2351,2359
<EOL>|2359,2360
-|2360,2361
Anxiety|2362,2369
<EOL>|2369,2370
-|2370,2371
Cervical|2372,2380
Radiculitis|2381,2392
<EOL>|2392,2393
-|2393,2394
Cervical|2395,2403
Spondylosis|2404,2415
<EOL>|2415,2416
-|2416,2417
Coronary|2418,2426
Artery|2427,2433
Disease|2434,2441
<EOL>|2441,2442
-|2442,2443
Headache|2444,2452
<EOL>|2452,2453
-|2453,2454
Herpes|2455,2461
Zoster|2462,2468
<EOL>|2468,2469
-|2469,2470
GI|2471,2473
Bleeding|2474,2482
<EOL>|2482,2483
-|2483,2484
Peripheral|2485,2495
Vascular|2496,2504
Disease|2505,2512
s|2513,2514
/|2514,2515
p|2515,2516
bilateral|2517,2526
iliac|2527,2532
stents|2533,2539
<EOL>|2539,2540
-|2540,2541
s|2542,2543
/|2543,2544
p|2544,2545
hip|2546,2549
replacement|2550,2561
<EOL>|2561,2562
<EOL>|2563,2564
Social|2564,2570
History|2571,2578
:|2578,2579
<EOL>|2579,2580
_|2580,2581
_|2581,2582
_|2582,2583
<EOL>|2583,2584
Family|2584,2590
History|2591,2598
:|2598,2599
<EOL>|2599,2600
Mother|2600,2606
with|2607,2611
asthma|2612,2618
and|2619,2622
hypertension|2623,2635
.|2635,2636
Father|2637,2643
with|2644,2648
colon|2649,2654
cancer|2655,2661
.|2661,2662
<EOL>|2663,2664
Brother|2664,2671
with|2672,2676
leukemia|2677,2685
.|2685,2686
<EOL>|2686,2687
<EOL>|2687,2688
<EOL>|2689,2690
Physical|2690,2698
Exam|2699,2703
:|2703,2704
<EOL>|2704,2705
PHYSICAL|2705,2713
EXAMINATION|2714,2725
ON|2726,2728
ADMISSION|2729,2738
:|2738,2739
<EOL>|2739,2740
=|2740,2741
=|2741,2742
=|2742,2743
=|2743,2744
=|2744,2745
=|2745,2746
=|2746,2747
=|2747,2748
=|2748,2749
=|2749,2750
=|2750,2751
=|2751,2752
=|2752,2753
=|2753,2754
=|2754,2755
=|2755,2756
=|2756,2757
=|2757,2758
=|2758,2759
=|2759,2760
=|2760,2761
=|2761,2762
=|2762,2763
=|2763,2764
=|2764,2765
=|2765,2766
=|2766,2767
=|2767,2768
=|2768,2769
=|2769,2770
=|2770,2771
=|2771,2772
=|2772,2773
=|2773,2774
<EOL>|2774,2775
VITALS|2776,2782
:|2782,2783
97.3|2784,2788
159|2789,2792
/|2792,2793
91|2793,2795
75|2796,2798
16|2800,2802
94|2804,2806
%|2806,2807
on|2808,2810
2L|2811,2813
<EOL>|2815,2816
GENERAL|2817,2824
:|2824,2825
Pleasant|2826,2834
,|2834,2835
well|2836,2840
-|2840,2841
appearing|2841,2850
,|2850,2851
in|2852,2854
no|2855,2857
apparent|2858,2866
distress|2867,2875
.|2875,2876
<EOL>|2878,2879
HEENT|2880,2885
:|2885,2886
Normocephalic|2887,2900
,|2900,2901
atraumatic|2902,2912
,|2912,2913
no|2914,2916
conjunctival|2917,2929
pallor|2930,2936
or|2937,2939
<EOL>|2940,2941
scleral|2941,2948
icterus|2949,2956
,|2956,2957
PERRLA|2958,2964
,|2964,2965
EOMI|2966,2970
,|2970,2971
OP|2972,2974
clear|2975,2980
.|2980,2981
<EOL>|2983,2984
NECK|2985,2989
:|2989,2990
Supple|2991,2997
,|2997,2998
no|2999,3001
LAD|3002,3005
,|3005,3006
no|3007,3009
thyromegaly|3010,3021
,|3021,3022
JVP|3023,3026
flat|3027,3031
.|3031,3032
<EOL>|3034,3035
CARDIAC|3036,3043
:|3043,3044
Normal|3045,3051
S1|3052,3054
/|3054,3055
S2|3055,3057
,|3057,3058
no|3059,3061
murmurs|3062,3069
rubs|3070,3074
or|3075,3077
gallops|3078,3085
.|3085,3086
<EOL>|3088,3089
PULMONARY|3090,3099
:|3099,3100
Mild|3101,3105
expiratory|3106,3116
wheezes|3117,3124
in|3125,3127
all|3128,3131
lung|3132,3136
fields|3137,3143
<EOL>|3145,3146
ABDOMEN|3147,3154
:|3154,3155
Normal|3156,3162
bowel|3163,3168
sounds|3169,3175
,|3175,3176
soft|3177,3181
,|3181,3182
non-tender|3183,3193
,|3193,3194
non-distended|3195,3208
,|3208,3209
<EOL>|3210,3211
no|3211,3213
organomegaly|3214,3226
.|3226,3227
<EOL>|3229,3230
EXTREMITIES|3231,3242
:|3242,3243
Warm|3244,3248
,|3248,3249
well|3250,3254
-|3254,3255
perfused|3255,3263
,|3263,3264
no|3265,3267
cyanosis|3268,3276
,|3276,3277
clubbing|3278,3286
or|3287,3289
<EOL>|3290,3291
edema|3291,3296
.|3296,3297
<EOL>|3299,3300
SKIN|3301,3305
:|3305,3306
Without|3307,3314
rash|3315,3319
.|3319,3320
<EOL>|3322,3323
NEUROLOGIC|3324,3334
:|3334,3335
A|3336,3337
&|3337,3338
Ox3|3338,3341
,|3341,3342
CN|3343,3345
II|3346,3348
-|3348,3349
XII|3349,3352
grossly|3353,3360
normal|3361,3367
,|3367,3368
normal|3369,3375
sensation|3376,3385
,|3385,3386
<EOL>|3387,3388
with|3388,3392
strength|3393,3401
_|3402,3403
_|3403,3404
_|3404,3405
throughout|3406,3416
.|3416,3417
<EOL>|3420,3421
<EOL>|3421,3422
PHYSICAL|3422,3430
EXAMINATION|3431,3442
ON|3443,3445
DISCHARGE|3446,3455
:|3455,3456
<EOL>|3456,3457
=|3457,3458
=|3458,3459
=|3459,3460
=|3460,3461
=|3461,3462
=|3462,3463
=|3463,3464
=|3464,3465
=|3465,3466
=|3466,3467
=|3467,3468
=|3468,3469
=|3469,3470
=|3470,3471
=|3471,3472
=|3472,3473
=|3473,3474
=|3474,3475
=|3475,3476
=|3476,3477
=|3477,3478
=|3478,3479
=|3479,3480
=|3480,3481
=|3481,3482
=|3482,3483
=|3483,3484
=|3484,3485
=|3485,3486
=|3486,3487
=|3487,3488
=|3488,3489
=|3489,3490
=|3490,3491
<EOL>|3491,3492
VITALS|3493,3499
:|3499,3500
98.6|3501,3505
127|3506,3509
-|3509,3510
150|3510,3513
/|3513,3514
50|3514,3516
-|3516,3517
60|3517,3519
70|3521,3523
-|3523,3524
90'S|3524,3528
16|3529,3531
98|3533,3535
%|3535,3536
on|3537,3539
3L|3540,3542
<EOL>|3544,3545
GENERAL|3546,3553
:|3553,3554
Pleasant|3555,3563
,|3563,3564
well|3565,3569
-|3569,3570
appearing|3570,3579
,|3579,3580
in|3581,3583
no|3584,3586
apparent|3587,3595
distress|3596,3604
.|3604,3605
<EOL>|3607,3608
HEENT|3609,3614
:|3614,3615
Normocephalic|3616,3629
,|3629,3630
atraumatic|3631,3641
,|3641,3642
no|3643,3645
conjunctival|3646,3658
pallor|3659,3665
or|3666,3668
<EOL>|3669,3670
scleral|3670,3677
icterus|3678,3685
,|3685,3686
PERRLA|3687,3693
,|3693,3694
EOMI|3695,3699
,|3699,3700
OP|3701,3703
clear|3704,3709
.|3709,3710
<EOL>|3712,3713
NECK|3714,3718
:|3718,3719
Supple|3720,3726
,|3726,3727
no|3728,3730
LAD|3731,3734
,|3734,3735
no|3736,3738
thyromegaly|3739,3750
,|3750,3751
JVP|3752,3755
flat|3756,3760
.|3760,3761
<EOL>|3763,3764
CARDIAC|3765,3772
:|3772,3773
Normal|3774,3780
S1|3781,3783
/|3783,3784
S2|3784,3786
,|3786,3787
no|3788,3790
murmurs|3791,3798
rubs|3799,3803
or|3804,3806
gallops|3807,3814
.|3814,3815
<EOL>|3817,3818
PULMONARY|3819,3828
:|3828,3829
Minimally|3830,3839
decreased|3840,3849
bilateral|3850,3859
air|3860,3863
entry|3864,3869
,|3869,3870
no|3871,3873
wheezes|3874,3881
<EOL>|3882,3883
in|3883,3885
all|3886,3889
lung|3890,3894
fields|3895,3901
<EOL>|3903,3904
ABDOMEN|3905,3912
:|3912,3913
Normal|3914,3920
bowel|3921,3926
sounds|3927,3933
,|3933,3934
soft|3935,3939
,|3939,3940
non-tender|3941,3951
,|3951,3952
non-distended|3953,3966
,|3966,3967
<EOL>|3968,3969
no|3969,3971
organomegaly|3972,3984
.|3984,3985
<EOL>|3987,3988
EXTREMITIES|3989,4000
:|4000,4001
Warm|4002,4006
,|4006,4007
well|4008,4012
-|4012,4013
perfused|4013,4021
,|4021,4022
no|4023,4025
cyanosis|4026,4034
,|4034,4035
clubbing|4036,4044
or|4045,4047
<EOL>|4048,4049
edema|4049,4054
.|4054,4055
<EOL>|4057,4058
SKIN|4059,4063
:|4063,4064
Without|4065,4072
rash|4073,4077
.|4077,4078
<EOL>|4080,4081
NEUROLOGIC|4082,4092
:|4092,4093
A|4094,4095
&|4095,4096
Ox3|4096,4099
,|4099,4100
CN|4101,4103
II|4104,4106
-|4106,4107
XII|4107,4110
grossly|4111,4118
normal|4119,4125
,|4125,4126
normal|4127,4133
sensation|4134,4143
,|4143,4144
<EOL>|4145,4146
with|4146,4150
strength|4151,4159
_|4160,4161
_|4161,4162
_|4162,4163
throughout|4164,4174
.|4174,4175
<EOL>|4177,4178
<EOL>|4179,4180
Pertinent|4180,4189
Results|4190,4197
:|4197,4198
<EOL>|4198,4199
LABS|4199,4203
ON|4204,4206
ADMISSION|4207,4216
:|4216,4217
<EOL>|4217,4218
=|4218,4219
=|4219,4220
=|4220,4221
=|4221,4222
=|4222,4223
=|4223,4224
=|4224,4225
=|4225,4226
=|4226,4227
=|4227,4228
=|4228,4229
=|4229,4230
=|4230,4231
=|4231,4232
=|4232,4233
=|4233,4234
=|4234,4235
=|4235,4236
<EOL>|4236,4237
_|4237,4238
_|4238,4239
_|4239,4240
06|4241,4243
:|4243,4244
15PM|4244,4248
BLOOD|4249,4254
WBC|4255,4258
-|4258,4259
7.7|4259,4262
RBC|4263,4266
-|4266,4267
4|4267,4268
.|4268,4269
92|4269,4271
Hgb|4272,4275
-|4275,4276
13.5|4276,4280
Hct|4281,4284
-|4284,4285
42.4|4285,4289
MCV|4290,4293
-|4293,4294
86|4294,4296
<EOL>|4297,4298
MCH|4298,4301
-|4301,4302
27.4|4302,4306
MCHC|4307,4311
-|4311,4312
31|4312,4314
.|4314,4315
8|4315,4316
*|4316,4317
RDW|4318,4321
-|4321,4322
19|4322,4324
.|4324,4325
6|4325,4326
*|4326,4327
RDWSD|4328,4333
-|4333,4334
61|4334,4336
.|4336,4337
2|4337,4338
*|4338,4339
Plt|4340,4343
_|4344,4345
_|4345,4346
_|4346,4347
<EOL>|4347,4348
_|4348,4349
_|4349,4350
_|4350,4351
06|4352,4354
:|4354,4355
15PM|4355,4359
BLOOD|4360,4365
Neuts|4366,4371
-|4371,4372
87|4372,4374
.|4374,4375
4|4375,4376
*|4376,4377
Lymphs|4378,4384
-|4384,4385
5|4385,4386
.|4386,4387
7|4387,4388
*|4388,4389
Monos|4390,4395
-|4395,4396
6.1|4396,4399
<EOL>|4400,4401
Eos|4401,4404
-|4404,4405
0|4405,4406
.|4406,4407
0|4407,4408
*|4408,4409
Baso|4410,4414
-|4414,4415
0.1|4415,4418
Im|4419,4421
_|4422,4423
_|4423,4424
_|4424,4425
AbsNeut|4426,4433
-|4433,4434
6|4434,4435
.|4435,4436
72|4436,4438
*|4438,4439
AbsLymp|4440,4447
-|4447,4448
0|4448,4449
.|4449,4450
44|4450,4452
*|4452,4453
<EOL>|4454,4455
AbsMono|4455,4462
-|4462,4463
0|4463,4464
.|4464,4465
47|4465,4467
AbsEos|4468,4474
-|4474,4475
0|4475,4476
.|4476,4477
00|4477,4479
*|4479,4480
AbsBaso|4481,4488
-|4488,4489
0.01|4489,4493
<EOL>|4493,4494
_|4494,4495
_|4495,4496
_|4496,4497
06|4498,4500
:|4500,4501
15PM|4501,4505
BLOOD|4506,4511
_|4512,4513
_|4513,4514
_|4514,4515
PTT|4516,4519
-|4519,4520
29.6|4520,4524
_|4525,4526
_|4526,4527
_|4527,4528
<EOL>|4528,4529
_|4529,4530
_|4530,4531
_|4531,4532
06|4533,4535
:|4535,4536
15PM|4536,4540
BLOOD|4541,4546
Plt|4547,4550
_|4551,4552
_|4552,4553
_|4553,4554
<EOL>|4554,4555
_|4555,4556
_|4556,4557
_|4557,4558
06|4559,4561
:|4561,4562
15PM|4562,4566
BLOOD|4567,4572
Glucose|4573,4580
-|4580,4581
122|4581,4584
*|4584,4585
UreaN|4586,4591
-|4591,4592
21|4592,4594
*|4594,4595
Creat|4596,4601
-|4601,4602
1|4602,4603
.|4603,4604
2|4604,4605
*|4605,4606
Na|4607,4609
-|4609,4610
136|4610,4613
<EOL>|4614,4615
K|4615,4616
-|4616,4617
3.4|4617,4620
Cl|4621,4623
-|4623,4624
92|4624,4626
*|4626,4627
HCO3|4628,4632
-|4632,4633
31|4633,4635
AnGap|4636,4641
-|4641,4642
16|4642,4644
<EOL>|4644,4645
_|4645,4646
_|4646,4647
_|4647,4648
06|4649,4651
:|4651,4652
15PM|4652,4656
BLOOD|4657,4662
ALT|4663,4666
-|4666,4667
52|4667,4669
*|4669,4670
AST|4671,4674
-|4674,4675
34|4675,4677
AlkPhos|4678,4685
-|4685,4686
69|4686,4688
TotBili|4689,4696
-|4696,4697
0.3|4697,4700
<EOL>|4700,4701
_|4701,4702
_|4702,4703
_|4703,4704
06|4705,4707
:|4707,4708
15PM|4708,4712
BLOOD|4713,4718
Lipase|4719,4725
-|4725,4726
28|4726,4728
<EOL>|4728,4729
_|4729,4730
_|4730,4731
_|4731,4732
06|4733,4735
:|4735,4736
15PM|4736,4740
BLOOD|4741,4746
cTropnT|4747,4754
-|4754,4755
<|4755,4756
0|4756,4757
.|4757,4758
01|4758,4760
proBNP|4761,4767
-|4767,4768
325|4768,4771
<EOL>|4771,4772
_|4772,4773
_|4773,4774
_|4774,4775
06|4776,4778
:|4778,4779
15PM|4779,4783
BLOOD|4784,4789
Albumin|4790,4797
-|4797,4798
4.2|4798,4801
<EOL>|4801,4802
<EOL>|4802,4803
LABS|4803,4807
ON|4808,4810
DISHCHARGE|4811,4821
:|4821,4822
<EOL>|4822,4823
=|4823,4824
=|4824,4825
=|4825,4826
=|4826,4827
=|4827,4828
=|4828,4829
=|4829,4830
=|4830,4831
=|4831,4832
=|4832,4833
=|4833,4834
=|4834,4835
=|4835,4836
=|4836,4837
=|4837,4838
=|4838,4839
=|4839,4840
=|4840,4841
=|4841,4842
<EOL>|4842,4843
_|4843,4844
_|4844,4845
_|4845,4846
06|4847,4849
:|4849,4850
40AM|4850,4854
BLOOD|4855,4860
WBC|4861,4864
-|4864,4865
10|4865,4867
.|4867,4868
3|4868,4869
*|4869,4870
RBC|4871,4874
-|4874,4875
4.20|4875,4879
Hgb|4880,4883
-|4883,4884
11.8|4884,4888
Hct|4889,4892
-|4892,4893
37.0|4893,4897
<EOL>|4898,4899
MCV|4899,4902
-|4902,4903
88|4903,4905
MCH|4906,4909
-|4909,4910
28.1|4910,4914
MCHC|4915,4919
-|4919,4920
31|4920,4922
.|4922,4923
9|4923,4924
*|4924,4925
RDW|4926,4929
-|4929,4930
19|4930,4932
.|4932,4933
9|4933,4934
*|4934,4935
RDWSD|4936,4941
-|4941,4942
65|4942,4944
.|4944,4945
1|4945,4946
*|4946,4947
Plt|4948,4951
_|4952,4953
_|4953,4954
_|4954,4955
<EOL>|4955,4956
_|4956,4957
_|4957,4958
_|4958,4959
06|4960,4962
:|4962,4963
40AM|4963,4967
BLOOD|4968,4973
Plt|4974,4977
_|4978,4979
_|4979,4980
_|4980,4981
<EOL>|4981,4982
_|4982,4983
_|4983,4984
_|4984,4985
06|4986,4988
:|4988,4989
40AM|4989,4993
BLOOD|4994,4999
Glucose|5000,5007
-|5007,5008
112|5008,5011
*|5011,5012
UreaN|5013,5018
-|5018,5019
18|5019,5021
Creat|5022,5027
-|5027,5028
0.9|5028,5031
Na|5032,5034
-|5034,5035
137|5035,5038
<EOL>|5039,5040
K|5040,5041
-|5041,5042
3.6|5042,5045
Cl|5046,5048
-|5048,5049
96|5049,5051
HCO3|5052,5056
-|5056,5057
28|5057,5059
AnGap|5060,5065
-|5065,5066
17|5066,5068
<EOL>|5068,5069
_|5069,5070
_|5070,5071
_|5071,5072
06|5073,5075
:|5075,5076
40AM|5076,5080
BLOOD|5081,5086
Calcium|5087,5094
-|5094,5095
9.5|5095,5098
Phos|5099,5103
-|5103,5104
2|5104,5105
.|5105,5106
6|5106,5107
*|5107,5108
Mg|5109,5111
-|5111,5112
2.1|5112,5115
<EOL>|5115,5116
<EOL>|5116,5117
IMAGING|5117,5124
:|5124,5125
<EOL>|5125,5126
=|5126,5127
=|5127,5128
=|5128,5129
=|5129,5130
=|5130,5131
=|5131,5132
=|5132,5133
=|5133,5134
<EOL>|5134,5135
_|5135,5136
_|5136,5137
_|5137,5138
CXR|5139,5142
:|5142,5143
<EOL>|5143,5144
No|5144,5146
acute|5147,5152
cardiopulmonary|5153,5168
process|5169,5176
.|5176,5177
<EOL>|5177,5178
<EOL>|5178,5179
<EOL>|5180,5181
Brief|5181,5186
Hospital|5187,5195
Course|5196,5202
:|5202,5203
<EOL>|5203,5204
_|5204,5205
_|5205,5206
_|5206,5207
yo|5208,5210
F|5211,5212
with|5213,5217
history|5218,5225
of|5226,5228
COPD|5229,5233
on|5234,5236
home|5237,5241
O2|5242,5244
,|5244,5245
atrial|5246,5252
fibrillation|5253,5265
on|5266,5268
<EOL>|5269,5270
apixaban|5270,5278
,|5278,5279
hypertension|5280,5292
,|5292,5293
CAD|5294,5297
,|5297,5298
hyperlipidemia|5299,5313
,|5313,5314
and|5315,5318
recurrent|5319,5328
<EOL>|5329,5330
hospitalization|5330,5345
for|5346,5349
COPD|5350,5354
exacerbation|5355,5367
over|5368,5372
the|5373,5376
last|5377,5381
4|5382,5383
months|5384,5390
,|5390,5391
<EOL>|5392,5393
who|5393,5396
presented|5397,5406
with|5407,5411
dyspnea|5412,5419
and|5420,5423
increased|5424,5433
wheezing|5434,5442
secondary|5443,5452
to|5453,5455
<EOL>|5456,5457
severe|5457,5463
COPD|5464,5468
.|5468,5469
<EOL>|5469,5470
<EOL>|5471,5472
#|5472,5473
Recurrent|5473,5482
COPD|5483,5487
exacerbation|5488,5500
:|5500,5501
Patient|5502,5509
presented|5510,5519
with|5520,5524
increased|5525,5534
<EOL>|5535,5536
dyspnea|5536,5543
and|5544,5547
diffuse|5548,5555
wheezing|5556,5564
,|5564,5565
likely|5566,5572
secondary|5573,5582
to|5583,5585
COPD|5586,5590
<EOL>|5591,5592
exacerbation|5592,5604
.|5604,5605
She|5606,5609
has|5610,5613
a|5614,5615
history|5616,5623
of|5624,5626
multiple|5627,5635
recurrent|5636,5645
COPD|5646,5650
<EOL>|5651,5652
hospitalizations|5652,5668
.|5668,5669
According|5670,5679
to|5680,5682
Pulmonary|5683,5692
,|5692,5693
patient|5694,5701
has|5702,5705
severe|5706,5712
<EOL>|5713,5714
COPD|5714,5718
based|5719,5724
on|5725,5727
her|5728,5731
obstructive|5732,5743
deficits|5744,5752
on|5753,5755
PFTs|5756,5760
as|5761,5763
well|5764,5768
as|5769,5771
her|5772,5775
<EOL>|5776,5777
severe|5777,5783
symptoms|5784,5792
even|5793,5797
at|5798,5800
rest|5801,5805
,|5805,5806
as|5807,5809
well|5810,5814
as|5815,5817
her|5818,5821
more|5822,5826
frequent|5827,5835
<EOL>|5836,5837
exacerbations|5837,5850
and|5851,5854
is|5855,5857
likely|5858,5864
approaching|5865,5876
end|5877,5880
-|5880,5881
stage|5881,5886
disease|5887,5894
.|5894,5895
We|5896,5898
<EOL>|5899,5900
continued|5900,5909
Advair|5910,5916
500|5917,5920
/|5920,5921
50|5921,5923
BID|5924,5927
,|5927,5928
Spiriva|5929,5936
,|5936,5937
standing|5938,5946
nebulizers|5947,5957
,|5957,5958
and|5959,5962
<EOL>|5963,5964
theophylline|5964,5976
.|5976,5977
Pulmonary|5978,5987
recommended|5988,5999
additional|6000,6010
budesonide|6011,6021
<EOL>|6022,6023
inhalers|6023,6031
to|6032,6034
allow|6035,6040
reduction|6041,6050
of|6051,6053
PO|6054,6056
prednisone|6057,6067
dose|6068,6072
.|6072,6073
Prednisone|6074,6084
<EOL>|6085,6086
dose|6086,6090
was|6091,6094
increased|6095,6104
back|6105,6109
to|6110,6112
40mg|6113,6117
(|6118,6119
where|6119,6124
patient|6125,6132
was|6133,6136
better|6137,6143
)|6143,6144
with|6145,6149
<EOL>|6150,6151
a|6151,6152
plan|6153,6157
for|6158,6161
slow|6162,6166
wean|6167,6171
by|6172,6174
5mg|6175,6178
every|6179,6184
2|6185,6186
weeks|6187,6192
.|6192,6193
Also|6194,6198
,|6198,6199
patient|6200,6207
was|6208,6211
<EOL>|6212,6213
started|6213,6220
on|6221,6223
chronic|6224,6231
azithromycin|6232,6244
for|6245,6248
chronic|6249,6256
anti-inflammation|6257,6274
;|6274,6275
<EOL>|6276,6277
after|6277,6282
discussion|6283,6293
with|6294,6298
Dr.|6299,6302
_|6303,6304
_|6304,6305
_|6305,6306
was|6307,6310
agreed|6311,6317
to|6318,6320
stop|6321,6325
<EOL>|6326,6327
azithromycin|6327,6339
on|6340,6342
discharge|6343,6352
due|6353,6356
to|6357,6359
inability|6360,6369
to|6370,6372
monitor|6373,6380
QT|6381,6383
the|6384,6387
<EOL>|6388,6389
week|6389,6393
after|6394,6399
discharge|6400,6409
,|6409,6410
with|6411,6415
plan|6416,6420
to|6421,6423
restart|6424,6431
azithromycin|6432,6444
once|6445,6449
Dr|6450,6452
.|6452,6453
<EOL>|6454,6455
_|6455,6456
_|6456,6457
_|6457,6458
is|6459,6461
able|6462,6466
to|6467,6469
see|6470,6473
the|6474,6477
patient|6478,6485
.|6485,6486
Patient|6487,6494
did|6495,6498
not|6499,6502
want|6503,6507
to|6508,6510
go|6511,6513
to|6514,6516
<EOL>|6517,6518
pulmonary|6518,6527
rehab|6528,6533
.|6533,6534
She|6535,6538
was|6539,6542
seen|6543,6547
by|6548,6550
Palliative|6551,6561
Care|6562,6566
who|6567,6570
recommended|6571,6582
<EOL>|6583,6584
initiation|6584,6594
of|6595,6597
morphine|6598,6606
liquid|6607,6613
suspension|6614,6624
as|6625,6627
needed|6628,6634
for|6635,6638
shortness|6639,6648
<EOL>|6649,6650
of|6650,6652
breath|6653,6659
.|6659,6660
<EOL>|6660,6661
<EOL>|6661,6662
#|6662,6663
Acute|6664,6669
kidney|6670,6676
injury|6677,6683
:|6683,6684
Creatinine|6685,6695
was|6696,6699
slightly|6700,6708
elevated|6709,6717
to|6718,6720
1.2|6721,6724
<EOL>|6725,6726
from|6726,6730
a|6731,6732
baseline|6733,6741
of|6742,6744
1.0|6745,6748
.|6748,6749
She|6750,6753
likely|6754,6760
had|6761,6764
poor|6765,6769
PO|6770,6772
intake|6773,6779
.|6779,6780
<EOL>|6781,6782
Creatinine|6782,6792
on|6793,6795
discharge|6796,6805
was|6806,6809
0.9|6810,6813
.|6813,6814
<EOL>|6814,6815
<EOL>|6816,6817
CHRONIC|6817,6824
ISSUES|6825,6831
:|6831,6832
<EOL>|6834,6835
=|6835,6836
=|6836,6837
=|6837,6838
=|6838,6839
=|6839,6840
=|6840,6841
=|6841,6842
=|6842,6843
=|6843,6844
=|6844,6845
=|6845,6846
=|6846,6847
=|6847,6848
=|6848,6849
=|6849,6850
=|6850,6851
=|6851,6852
=|6852,6853
<EOL>|6855,6856
#|6856,6857
Anxiety|6858,6865
/|6865,6866
Insomnia|6866,6874
:|6874,6875
We|6876,6878
continued|6879,6888
home|6889,6893
lorazepam|6894,6903
.|6903,6904
<EOL>|6904,6905
<EOL>|6906,6907
#|6907,6908
Atrial|6909,6915
fibrillation|6916,6928
:|6928,6929
We|6930,6932
continued|6933,6942
diltiazem|6943,6952
for|6953,6956
rate|6957,6961
control|6962,6969
<EOL>|6970,6971
and|6971,6974
apixaban|6975,6983
for|6984,6987
anticoagulation|6988,7003
.|7003,7004
<EOL>|7006,7007
<EOL>|7008,7009
#|7009,7010
Hypertension|7011,7023
:|7023,7024
We|7025,7027
continued|7028,7037
home|7038,7042
imdur|7043,7048
,|7048,7049
hydrochlorothiazide|7050,7069
,|7069,7070
<EOL>|7071,7072
and|7072,7075
diltiazem|7076,7085
.|7085,7086
<EOL>|7088,7089
<EOL>|7090,7091
#|7091,7092
CAD|7093,7096
:|7096,7097
Cardiac|7098,7105
catheterization|7106,7121
in|7122,7124
_|7125,7126
_|7126,7127
_|7127,7128
showed|7129,7135
no|7136,7138
evidence|7139,7147
of|7148,7150
<EOL>|7151,7152
significant|7152,7163
stenosis|7164,7172
of|7173,7175
coronaries|7176,7186
.|7186,7187
ECHO|7188,7192
on|7193,7195
_|7196,7197
_|7197,7198
_|7198,7199
showed|7200,7206
EF|7207,7209
>|7210,7211
<EOL>|7212,7213
55|7213,7215
%|7215,7216
and|7217,7220
no|7221,7223
regional|7224,7232
or|7233,7235
global|7236,7242
wall|7243,7247
motion|7248,7254
abnormalities|7255,7268
.|7268,7269
We|7270,7272
<EOL>|7273,7274
continued|7274,7283
home|7284,7288
aspirin|7289,7296
and|7297,7300
atorvastatin|7301,7313
.|7313,7314
<EOL>|7314,7315
<EOL>|7316,7317
#|7317,7318
Anemia|7319,7325
:|7325,7326
We|7327,7329
continued|7330,7339
home|7340,7344
iron|7345,7349
supplements|7350,7361
.|7361,7362
<EOL>|7363,7364
<EOL>|7364,7365
*|7365,7366
*|7366,7367
*|7367,7368
TRANSITIONAL|7368,7380
ISSUES|7381,7387
:|7387,7388
*|7388,7389
*|7389,7390
*|7390,7391
<EOL>|7392,7393
-|7393,7394
Continue|7395,7403
Advair|7404,7410
500|7411,7414
/|7414,7415
50|7415,7417
BID|7418,7421
,|7421,7422
Spiriva|7423,7430
,|7430,7431
and|7432,7435
theophylline|7436,7448
<EOL>|7449,7450
-|7450,7451
Make|7452,7456
sure|7457,7461
patient|7462,7469
receives|7470,7478
standing|7479,7487
nebulizers|7488,7498
<EOL>|7499,7500
-|7500,7501
Added|7502,7507
additional|7508,7518
budesonide|7519,7529
inhalers|7530,7538
to|7539,7541
allow|7542,7547
reduction|7548,7557
of|7558,7560
PO|7561,7563
<EOL>|7564,7565
prednisone|7565,7575
dose|7576,7580
<EOL>|7581,7582
-|7582,7583
Start|7584,7589
chronic|7590,7597
azithromycin|7598,7610
for|7611,7614
chronic|7615,7622
anti-inflammation|7623,7640
.|7640,7641
<EOL>|7642,7643
(|7643,7644
Patient|7644,7651
was|7652,7655
started|7656,7663
on|7664,7666
azithromycin|7667,7679
in|7680,7682
the|7683,7686
hospital|7687,7695
and|7696,7699
QTc|7700,7703
on|7704,7706
<EOL>|7707,7708
_|7708,7709
_|7709,7710
_|7710,7711
was|7712,7715
472|7716,7719
ms|7720,7722
.|7722,7723
_|7724,7725
_|7725,7726
_|7726,7727
discussion|7728,7738
with|7739,7743
Dr.|7744,7747
_|7748,7749
_|7749,7750
_|7750,7751
was|7752,7755
agreed|7756,7762
<EOL>|7763,7764
to|7764,7766
stop|7767,7771
azithromycin|7772,7784
on|7785,7787
discharge|7788,7797
due|7798,7801
to|7802,7804
inability|7805,7814
to|7815,7817
monitor|7818,7825
QT|7826,7828
<EOL>|7829,7830
the|7830,7833
week|7834,7838
after|7839,7844
discharge|7845,7854
,|7854,7855
with|7856,7860
the|7861,7864
plan|7865,7869
to|7870,7872
restart|7873,7880
azithromycin|7881,7893
<EOL>|7894,7895
once|7895,7899
Dr.|7900,7903
_|7904,7905
_|7905,7906
_|7906,7907
is|7908,7910
able|7911,7915
to|7916,7918
see|7919,7922
the|7923,7926
patient|7927,7934
.|7934,7935
)|7935,7936
<EOL>|7936,7937
-|7937,7938
Would|7939,7944
recommend|7945,7954
audiology|7955,7964
testing|7965,7972
at|7973,7975
some|7976,7980
point|7981,7986
while|7987,7992
patient|7993,8000
<EOL>|8001,8002
is|8002,8004
on|8005,8007
chronic|8008,8015
azithromycin|8016,8028
<EOL>|8028,8029
-|8029,8030
Continue|8031,8039
supplemental|8040,8052
oxygen|8053,8059
for|8060,8063
comfort|8064,8071
<EOL>|8071,8072
-|8072,8073
Follow|8074,8080
up|8081,8083
with|8084,8088
Dr.|8089,8092
_|8093,8094
_|8094,8095
_|8095,8096
discharge|8097,8106
<EOL>|8107,8108
-|8108,8109
Continue|8110,8118
Bactrim|8119,8126
PPX|8127,8130
(|8131,8132
1|8132,8133
tab|8134,8137
SS|8138,8140
daily|8141,8146
)|8146,8147
given|8148,8153
extended|8154,8162
courses|8163,8170
<EOL>|8171,8172
of|8172,8174
steroids|8175,8183
<EOL>|8184,8185
-|8185,8186
Patient|8187,8194
was|8195,8198
discharged|8199,8209
on|8210,8212
prednisone|8213,8223
40|8224,8226
mg|8227,8229
with|8230,8234
plan|8235,8239
for|8240,8243
taper|8244,8249
<EOL>|8250,8251
by|8251,8253
5mg|8254,8257
every|8258,8263
2|8264,8265
weeks|8266,8271
:|8271,8272
<EOL>|8272,8273
Prednisone|8274,8284
40|8285,8287
mg|8288,8290
for|8291,8294
two|8295,8298
weeks|8299,8304
(|8305,8306
Day|8306,8309
1|8310,8311
=|8311,8312
_|8313,8314
_|8314,8315
_|8315,8316
end|8317,8320
<EOL>|8321,8322
_|8322,8323
_|8323,8324
_|8324,8325
<EOL>|8325,8326
Prednisone|8327,8337
35|8338,8340
mg|8341,8343
for|8344,8347
two|8348,8351
weeks|8352,8357
(|8358,8359
Day|8359,8362
1|8363,8364
=|8364,8365
_|8366,8367
_|8367,8368
_|8368,8369
end|8370,8373
<EOL>|8374,8375
_|8375,8376
_|8376,8377
_|8377,8378
<EOL>|8378,8379
Prednisone|8380,8390
30|8391,8393
mg|8394,8396
for|8397,8400
two|8401,8404
weeks|8405,8410
(|8411,8412
Day|8412,8415
1|8416,8417
=|8417,8418
_|8419,8420
_|8420,8421
_|8421,8422
end|8423,8426
<EOL>|8427,8428
_|8428,8429
_|8429,8430
_|8430,8431
<EOL>|8431,8432
etc|8433,8436
...|8436,8439
<EOL>|8439,8440
#|8440,8441
CONTACT|8442,8449
:|8449,8450
_|8451,8452
_|8452,8453
_|8453,8454
(|8455,8456
husband|8456,8463
/|8463,8464
HCP|8464,8467
)|8467,8468
_|8469,8470
_|8470,8471
_|8471,8472
<EOL>|8473,8474
#|8474,8475
CODE|8476,8480
STATUS|8481,8487
:|8487,8488
Full|8489,8493
confirmed|8494,8503
<EOL>|8504,8505
<EOL>|8506,8507
Medications|8507,8518
on|8519,8521
Admission|8522,8531
:|8531,8532
<EOL>|8532,8533
The|8533,8536
Preadmission|8537,8549
Medication|8550,8560
list|8561,8565
is|8566,8568
accurate|8569,8577
and|8578,8581
complete|8582,8590
.|8590,8591
<EOL>|8591,8592
1.|8592,8594
Acetaminophen|8595,8608
325|8609,8612
mg|8613,8615
PO|8616,8618
Q4H|8619,8622
:|8622,8623
PRN|8623,8626
Pain|8627,8631
<EOL>|8632,8633
2.|8633,8635
albuterol|8636,8645
sulfate|8646,8653
90|8654,8656
mcg|8657,8660
/|8660,8661
actuation|8661,8670
inhalation|8671,8681
Q4H|8682,8685
<EOL>|8686,8687
3.|8687,8689
Apixaban|8690,8698
5|8699,8700
mg|8701,8703
PO|8704,8706
BID|8707,8710
<EOL>|8711,8712
4.|8712,8714
Aspirin|8715,8722
81|8723,8725
mg|8726,8728
PO|8729,8731
DAILY|8732,8737
<EOL>|8738,8739
5.|8739,8741
Atorvastatin|8742,8754
10|8755,8757
mg|8758,8760
PO|8761,8763
QPM|8764,8767
<EOL>|8768,8769
6.|8769,8771
Diltiazem|8772,8781
Extended|8782,8790
-|8790,8791
Release|8791,8798
240|8799,8802
mg|8803,8805
PO|8806,8808
BID|8809,8812
<EOL>|8813,8814
7.|8814,8816
Docusate|8817,8825
Sodium|8826,8832
100|8833,8836
mg|8837,8839
PO|8840,8842
BID|8843,8846
<EOL>|8847,8848
8.|8848,8850
Dorzolamide|8851,8862
2|8863,8864
%|8864,8865
Ophth|8866,8871
.|8871,8872
Soln.|8873,8878
1|8879,8880
DROP|8881,8885
BOTH|8886,8890
EYES|8891,8895
BID|8896,8899
<EOL>|8900,8901
9.|8901,8903
Ferrous|8904,8911
Sulfate|8912,8919
325|8920,8923
mg|8924,8926
PO|8927,8929
DAILY|8930,8935
<EOL>|8936,8937
10.|8937,8940
Fluticasone|8941,8952
Propionate|8953,8963
NASAL|8964,8969
2|8970,8971
SPRY|8972,8976
NU|8977,8979
DAILY|8980,8985
:|8985,8986
PRN|8986,8989
allergies|8990,8999
<EOL>|9000,9001
11|9001,9003
.|9003,9004
Fluticasone|9005,9016
-|9016,9017
Salmeterol|9017,9027
Diskus|9028,9034
(|9035,9036
500|9036,9039
/|9039,9040
50|9040,9042
)|9042,9043
1|9045,9046
INH|9047,9050
IH|9051,9053
BID|9054,9057
<EOL>|9058,9059
12.|9059,9062
Guaifenesin|9063,9074
_|9075,9076
_|9076,9077
_|9077,9078
mL|9079,9081
PO|9082,9084
Q4H|9085,9088
:|9088,9089
PRN|9089,9092
cough|9093,9098
<EOL>|9099,9100
13.|9100,9103
Hydrochlorothiazide|9104,9123
50|9124,9126
mg|9127,9129
PO|9130,9132
DAILY|9133,9138
<EOL>|9139,9140
14.|9140,9143
Isosorbide|9144,9154
Mononitrate|9155,9166
(|9167,9168
Extended|9168,9176
Release|9177,9184
)|9184,9185
240|9186,9189
mg|9190,9192
PO|9193,9195
DAILY|9196,9201
<EOL>|9202,9203
15.|9203,9206
Latanoprost|9207,9218
0.005|9219,9224
%|9224,9225
Ophth|9226,9231
.|9231,9232
Soln.|9233,9238
1|9239,9240
DROP|9241,9245
BOTH|9246,9250
EYES|9251,9255
QHS|9256,9259
<EOL>|9260,9261
16|9261,9263
.|9263,9264
Lorazepam|9265,9274
0.5|9275,9278
mg|9279,9281
PO|9282,9284
Q8H|9285,9288
:|9288,9289
PRN|9289,9292
Insomnia|9293,9301
,|9301,9302
anxiety|9303,9310
,|9310,9311
vertigo|9312,9319
<EOL>|9320,9321
17.|9321,9324
Multivitamins|9325,9338
1|9339,9340
TAB|9341,9344
PO|9345,9347
DAILY|9348,9353
<EOL>|9354,9355
18.|9355,9358
PredniSONE|9359,9369
30|9370,9372
mg|9373,9375
PO|9376,9378
DAILY|9379,9384
<EOL>|9385,9386
Tapered|9386,9393
dose|9394,9398
-|9399,9400
DOWN|9401,9405
<EOL>|9406,9407
19|9407,9409
.|9409,9410
Ranitidine|9411,9421
300|9422,9425
mg|9426,9428
PO|9429,9431
DAILY|9432,9437
<EOL>|9438,9439
20|9439,9441
.|9441,9442
Theophylline|9443,9455
SR|9456,9458
300|9459,9462
mg|9463,9465
PO|9466,9468
BID|9469,9472
<EOL>|9473,9474
21|9474,9476
.|9476,9477
Tiotropium|9478,9488
Bromide|9489,9496
1|9497,9498
CAP|9499,9502
IH|9503,9505
DAILY|9506,9511
<EOL>|9512,9513
22.|9513,9516
Levofloxacin|9517,9529
750|9530,9533
mg|9534,9536
PO|9537,9539
DAILY|9540,9545
<EOL>|9546,9547
23|9547,9549
.|9549,9550
Sulfameth|9551,9560
/|9560,9561
Trimethoprim|9561,9573
SS|9574,9576
1|9577,9578
TAB|9579,9582
PO|9583,9585
DAILY|9586,9591
prophylaxis|9592,9603
for|9604,9607
<EOL>|9608,9609
long|9609,9613
term|9614,9618
steroid|9619,9626
use|9627,9630
<EOL>|9631,9632
24|9632,9634
.|9634,9635
Calcitrate|9636,9646
-|9646,9647
Vitamin|9647,9654
D|9655,9656
(|9657,9658
calcium|9658,9665
citrate|9666,9673
-|9673,9674
vitamin|9674,9681
D3|9682,9684
)|9684,9685
315|9686,9689
mg|9690,9692
-|9693,9694
<EOL>|9695,9696
200|9696,9699
units|9700,9705
oral|9707,9711
DAILY|9712,9717
<EOL>|9718,9719
25.|9719,9722
cod|9723,9726
liver|9727,9732
oil|9733,9736
1|9737,9738
capsule|9739,9746
oral|9748,9752
BID|9753,9756
<EOL>|9757,9758
26|9758,9760
.|9760,9761
Ipratropium|9762,9773
Bromide|9774,9781
Neb|9782,9785
1|9786,9787
NEB|9788,9791
IH|9792,9794
Q6H|9795,9798
:|9798,9799
PRN|9799,9802
Wheezing|9803,9811
<EOL>|9812,9813
<EOL>|9813,9814
<EOL>|9815,9816
Discharge|9816,9825
Medications|9826,9837
:|9837,9838
<EOL>|9838,9839
1.|9839,9841
Acetaminophen|9842,9855
325|9856,9859
mg|9860,9862
PO|9863,9865
Q4H|9866,9869
:|9869,9870
PRN|9870,9873
Pain|9874,9878
<EOL>|9879,9880
2.|9880,9882
Calcitrate|9883,9893
-|9893,9894
Vitamin|9894,9901
D|9902,9903
(|9904,9905
calcium|9905,9912
citrate|9913,9920
-|9920,9921
vitamin|9921,9928
D3|9929,9931
)|9931,9932
315|9933,9936
mg|9937,9939
-|9940,9941
<EOL>|9942,9943
200|9943,9946
units|9947,9952
oral|9954,9958
DAILY|9959,9964
<EOL>|9965,9966
3.|9966,9968
Tiotropium|9969,9979
Bromide|9980,9987
1|9988,9989
CAP|9990,9993
IH|9994,9996
DAILY|9997,10002
<EOL>|10003,10004
4.|10004,10006
Theophylline|10007,10019
SR|10020,10022
300|10023,10026
mg|10027,10029
PO|10030,10032
BID|10033,10036
<EOL>|10037,10038
5.|10038,10040
Sulfameth|10041,10050
/|10050,10051
Trimethoprim|10051,10063
SS|10064,10066
1|10067,10068
TAB|10069,10072
PO|10073,10075
DAILY|10076,10081
prophylaxis|10082,10093
for|10094,10097
long|10098,10102
<EOL>|10103,10104
term|10104,10108
steroid|10109,10116
use|10117,10120
<EOL>|10121,10122
6.|10122,10124
Ranitidine|10125,10135
300|10136,10139
mg|10140,10142
PO|10143,10145
DAILY|10146,10151
<EOL>|10152,10153
7.|10153,10155
PredniSONE|10156,10166
40|10167,10169
mg|10170,10172
PO|10173,10175
DAILY|10176,10181
<EOL>|10182,10183
8.|10183,10185
Lorazepam|10186,10195
0.5|10196,10199
mg|10200,10202
PO|10203,10205
Q8H|10206,10209
:|10209,10210
PRN|10210,10213
Insomnia|10214,10222
,|10222,10223
anxiety|10224,10231
,|10231,10232
vertigo|10233,10240
<EOL>|10241,10242
9.|10242,10244
Latanoprost|10245,10256
0.005|10257,10262
%|10262,10263
Ophth|10264,10269
.|10269,10270
Soln.|10271,10276
1|10277,10278
DROP|10279,10283
BOTH|10284,10288
EYES|10289,10293
QHS|10294,10297
<EOL>|10298,10299
10.|10299,10302
Isosorbide|10303,10313
Mononitrate|10314,10325
(|10326,10327
Extended|10327,10335
Release|10336,10343
)|10343,10344
240|10345,10348
mg|10349,10351
PO|10352,10354
DAILY|10355,10360
<EOL>|10361,10362
11.|10362,10365
Ipratropium|10366,10377
Bromide|10378,10385
Neb|10386,10389
1|10390,10391
NEB|10392,10395
IH|10396,10398
Q6H|10399,10402
Wheezing|10403,10411
<EOL>|10412,10413
12.|10413,10416
Hydrochlorothiazide|10417,10436
50|10437,10439
mg|10440,10442
PO|10443,10445
DAILY|10446,10451
<EOL>|10452,10453
13.|10453,10456
Guaifenesin|10457,10468
_|10469,10470
_|10470,10471
_|10471,10472
mL|10473,10475
PO|10476,10478
Q4H|10479,10482
:|10482,10483
PRN|10483,10486
cough|10487,10492
<EOL>|10493,10494
14.|10494,10497
Fluticasone|10498,10509
-|10509,10510
Salmeterol|10510,10520
Diskus|10521,10527
(|10528,10529
500|10529,10532
/|10532,10533
50|10533,10535
)|10535,10536
1|10538,10539
INH|10540,10543
IH|10544,10546
BID|10547,10550
<EOL>|10551,10552
15.|10552,10555
Fluticasone|10556,10567
Propionate|10568,10578
NASAL|10579,10584
2|10585,10586
SPRY|10587,10591
NU|10592,10594
DAILY|10595,10600
:|10600,10601
PRN|10601,10604
allergies|10605,10614
<EOL>|10615,10616
16|10616,10618
.|10618,10619
Ferrous|10620,10627
Sulfate|10628,10635
325|10636,10639
mg|10640,10642
PO|10643,10645
DAILY|10646,10651
<EOL>|10652,10653
17.|10653,10656
Dorzolamide|10657,10668
2|10669,10670
%|10670,10671
Ophth|10672,10677
.|10677,10678
Soln.|10679,10684
1|10685,10686
DROP|10687,10691
BOTH|10692,10696
EYES|10697,10701
BID|10702,10705
<EOL>|10706,10707
18.|10707,10710
albuterol|10711,10720
sulfate|10721,10728
90|10729,10731
mcg|10732,10735
/|10735,10736
actuation|10736,10745
inhalation|10746,10756
Q4H|10757,10760
<EOL>|10761,10762
19|10762,10764
.|10764,10765
Apixaban|10766,10774
5|10775,10776
mg|10777,10779
PO|10780,10782
BID|10783,10786
<EOL>|10787,10788
20|10788,10790
.|10790,10791
Aspirin|10792,10799
81|10800,10802
mg|10803,10805
PO|10806,10808
DAILY|10809,10814
<EOL>|10815,10816
21|10816,10818
.|10818,10819
Atorvastatin|10820,10832
10|10833,10835
mg|10836,10838
PO|10839,10841
QPM|10842,10845
<EOL>|10846,10847
22.|10847,10850
Diltiazem|10851,10860
Extended|10861,10869
-|10869,10870
Release|10870,10877
240|10878,10881
mg|10882,10884
PO|10885,10887
BID|10888,10891
<EOL>|10892,10893
23|10893,10895
.|10895,10896
Docusate|10897,10905
Sodium|10906,10912
100|10913,10916
mg|10917,10919
PO|10920,10922
BID|10923,10926
<EOL>|10927,10928
24|10928,10930
.|10930,10931
Sodium|10932,10938
Chloride|10939,10947
Nasal|10948,10953
_|10954,10955
_|10955,10956
_|10956,10957
SPRY|10958,10962
NU|10963,10965
QID|10966,10969
:|10969,10970
PRN|10970,10973
nasal|10974,10979
discomfort|10980,10990
<EOL>|10991,10992
RX|10992,10994
*|10995,10996
sodium|10996,11002
chloride|11003,11011
0.65|11012,11016
%|11017,11018
_|11019,11020
_|11020,11021
_|11021,11022
spray|11023,11028
QID|11029,11032
nasal|11033,11038
congestion|11039,11049
Disp|11050,11054
<EOL>|11055,11056
#|11056,11057
*|11057,11058
1|11058,11059
Spray|11060,11065
Refills|11066,11073
:|11073,11074
*|11074,11075
0|11075,11076
<EOL>|11076,11077
25|11077,11079
.|11079,11080
Morphine|11081,11089
Sulfate|11090,11097
(|11098,11099
Oral|11099,11103
Solution|11104,11112
)|11112,11113
2|11114,11115
mg|11116,11118
/|11118,11119
mL|11119,11121
5|11122,11123
mg|11124,11126
PO|11127,11129
Q4H|11130,11133
:|11133,11134
PRN|11134,11137
<EOL>|11138,11139
shortness|11139,11148
of|11149,11151
breath|11152,11158
<EOL>|11159,11160
RX|11160,11162
*|11163,11164
morphine|11164,11172
10|11173,11175
mg|11176,11178
/|11178,11179
5|11179,11180
mL|11181,11183
2.5|11184,11187
mL|11188,11190
by|11191,11193
mouth|11194,11199
every|11200,11205
four|11206,11210
(|11211,11212
4|11212,11213
)|11213,11214
hours|11215,11220
<EOL>|11221,11222
Disp|11222,11226
_|11227,11228
_|11228,11229
_|11229,11230
Milliliter|11231,11241
Milliliter|11242,11252
Refills|11253,11260
:|11260,11261
*|11261,11262
0|11262,11263
<EOL>|11263,11264
26|11264,11266
.|11266,11267
Budesonide|11268,11278
Nasal|11279,11284
Inhaler|11285,11292
180|11293,11296
mcg|11297,11300
Other|11301,11306
DAILY|11307,11312
<EOL>|11313,11314
RX|11314,11316
*|11317,11318
budesonide|11318,11328
[|11329,11330
Pulmicort|11330,11339
Flexhaler|11340,11349
]|11349,11350
180|11351,11354
mcg|11355,11358
/|11358,11359
actuation|11359,11368
(|11369,11370
160|11370,11373
mcg|11374,11377
<EOL>|11378,11379
delivered|11379,11388
)|11388,11389
1|11390,11391
puff|11392,11396
INH|11397,11400
DAILY|11401,11406
Disp|11407,11411
#|11412,11413
*|11413,11414
1|11414,11415
Inhaler|11416,11423
Refills|11424,11431
:|11431,11432
*|11432,11433
0|11433,11434
<EOL>|11434,11435
<EOL>|11435,11436
<EOL>|11437,11438
Discharge|11438,11447
Disposition|11448,11459
:|11459,11460
<EOL>|11460,11461
Home|11461,11465
With|11466,11470
Service|11471,11478
<EOL>|11478,11479
<EOL>|11480,11481
Facility|11481,11489
:|11489,11490
<EOL>|11490,11491
_|11491,11492
_|11492,11493
_|11493,11494
<EOL>|11494,11495
<EOL>|11496,11497
Discharge|11497,11506
Diagnosis|11507,11516
:|11516,11517
<EOL>|11517,11518
PRIMARY|11518,11525
DIAGNOSIS|11526,11535
:|11535,11536
<EOL>|11536,11537
Severe|11537,11543
COPD|11544,11548
<EOL>|11548,11549
<EOL>|11549,11550
SECONDARY|11550,11559
DIAGNOSES|11560,11569
:|11569,11570
<EOL>|11570,11571
CAD|11571,11574
<EOL>|11574,11575
Hypertension|11575,11587
<EOL>|11587,11588
Atrial|11588,11594
fibrillation|11595,11607
<EOL>|11607,11608
<EOL>|11608,11609
<EOL>|11610,11611
Discharge|11611,11620
Condition|11621,11630
:|11630,11631
<EOL>|11631,11632
Mental|11632,11638
Status|11639,11645
:|11645,11646
Clear|11647,11652
and|11653,11656
coherent|11657,11665
.|11665,11666
<EOL>|11666,11667
Level|11667,11672
of|11673,11675
Consciousness|11676,11689
:|11689,11690
Alert|11691,11696
and|11697,11700
interactive|11701,11712
.|11712,11713
<EOL>|11713,11714
Activity|11714,11722
Status|11723,11729
:|11729,11730
Ambulatory|11731,11741
-|11742,11743
Independent|11744,11755
.|11755,11756
<EOL>|11756,11757
<EOL>|11757,11758
<EOL>|11759,11760
Discharge|11760,11769
Instructions|11770,11782
:|11782,11783
<EOL>|11783,11784
Dear|11784,11788
_|11789,11790
_|11790,11791
_|11791,11792
,|11792,11793
<EOL>|11793,11794
<EOL>|11794,11795
_|11795,11796
_|11796,11797
_|11797,11798
was|11799,11802
a|11803,11804
great|11805,11810
pleasure|11811,11819
taking|11820,11826
care|11827,11831
of|11832,11834
you|11835,11838
at|11839,11841
_|11842,11843
_|11843,11844
_|11844,11845
<EOL>|11846,11847
_|11847,11848
_|11848,11849
_|11849,11850
.|11850,11851
You|11852,11855
came|11856,11860
to|11861,11863
the|11864,11867
hospital|11868,11876
because|11877,11884
you|11885,11888
<EOL>|11889,11890
were|11890,11894
experiencing|11895,11907
worsening|11908,11917
shortness|11918,11927
of|11928,11930
breath|11931,11937
.|11937,11938
Pulmonary|11939,11948
team|11949,11953
<EOL>|11954,11955
saw|11955,11958
you|11959,11962
and|11963,11966
reviewed|11967,11975
your|11976,11980
condition|11981,11990
,|11990,11991
and|11992,11995
your|11996,12000
symptoms|12001,12009
are|12010,12013
<EOL>|12014,12015
thought|12015,12022
to|12023,12025
be|12026,12028
related|12029,12036
to|12037,12039
severe|12040,12046
COPD|12047,12051
.|12051,12052
We|12053,12055
did|12056,12059
some|12060,12064
changes|12065,12072
in|12073,12075
<EOL>|12076,12077
your|12077,12081
medications|12082,12093
and|12094,12097
increased|12098,12107
the|12108,12111
dose|12112,12116
of|12117,12119
prednisone|12120,12130
.|12130,12131
The|12132,12135
<EOL>|12136,12137
Palliative|12137,12147
Care|12148,12152
team|12153,12157
was|12158,12161
consulted|12162,12171
and|12172,12175
started|12176,12183
you|12184,12187
on|12188,12190
morphine|12191,12199
<EOL>|12200,12201
liquid|12201,12207
suspension|12208,12218
to|12219,12221
help|12222,12226
with|12227,12231
your|12232,12236
breathing|12237,12246
symptoms|12247,12255
.|12255,12256
<EOL>|12256,12257
<EOL>|12257,12258
Please|12258,12264
take|12265,12269
all|12270,12273
your|12274,12278
medications|12279,12290
on|12291,12293
time|12294,12298
and|12299,12302
follow|12303,12309
up|12310,12312
with|12313,12317
your|12318,12322
<EOL>|12323,12324
doctors|12324,12331
as|12332,12334
_|12335,12336
_|12336,12337
_|12337,12338
.|12338,12339
<EOL>|12339,12340
<EOL>|12340,12341
Best|12341,12345
regards|12346,12353
,|12353,12354
<EOL>|12354,12355
Your|12355,12359
_|12360,12361
_|12361,12362
_|12362,12363
team|12364,12368
<EOL>|12368,12369
<EOL>|12370,12371
Followup|12371,12379
Instructions|12380,12392
:|12392,12393
<EOL>|12393,12394
_|12394,12395
_|12395,12396
_|12396,12397
<EOL>|12397,12398

