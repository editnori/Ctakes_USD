 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
<EOL>|272,273
<EOL>|274,275
Chief|275,280
Complaint|281,290
:|290,291
<EOL>|291,292
Dyspnea|292,299
,|299,300
Atrial|301,307
Fibrillation|308,320
<EOL>|320,321
<EOL>|322,323
Major|323,328
Surgical|329,337
or|338,340
Invasive|341,349
Procedure|350,359
:|359,360
<EOL>|360,361
None|361,365
<EOL>|365,366
<EOL>|366,367
<EOL>|368,369
History|369,376
of|377,379
Present|380,387
Illness|388,395
:|395,396
<EOL>|396,397
_|397,398
_|398,399
_|399,400
F|401,402
with|403,407
pmhx|408,412
of|413,415
COPD|416,420
(|421,422
nighttime|422,431
O2|432,434
)|434,435
,|435,436
htn|437,440
,|440,441
afib|442,446
who|447,450
presents|451,459
<EOL>|460,461
with|461,465
dyspnea|466,473
,|473,474
currently|475,484
being|485,490
treated|491,498
for|499,502
COPD|503,507
and|508,511
admitted|512,520
for|521,524
<EOL>|525,526
Afib|526,530
with|531,535
RVR|536,539
.|539,540
<EOL>|542,543
The|544,547
patient|548,555
went|556,560
to|561,563
the|564,567
ED|568,570
on|571,573
_|574,575
_|575,576
_|576,577
and|578,581
was|582,585
diagnosed|586,595
with|596,600
a|601,602
<EOL>|603,604
COPD|604,608
flare|609,614
.|614,615
She|616,619
was|620,623
discharged|624,634
with|635,639
a|640,641
prednisone|642,652
taper|653,658
<EOL>|659,660
(|660,661
currently|661,670
on|671,673
60mg|674,678
)|678,679
and|680,683
azithromycin|684,696
.|696,697
This|698,702
AM|703,705
she|706,709
initially|710,719
felt|720,724
<EOL>|725,726
well|726,730
,|730,731
then|732,736
developed|737,746
dyspnea|747,754
at|755,757
rest|758,762
,|762,763
worsening|764,773
with|774,778
exertion|779,787
.|787,788
<EOL>|789,790
Her|790,793
inhalers|794,802
improved|803,811
her|812,815
SOB|816,819
.|819,820
She|821,824
felt|825,829
that|830,834
these|835,840
symptoms|841,849
were|850,854
<EOL>|855,856
consistent|856,866
with|867,871
her|872,875
COPD|876,880
.|880,881
She|882,885
saw|886,889
her|890,893
PCP|894,897
_|898,899
_|899,900
_|900,901
today|902,907
in|908,910
<EOL>|911,912
clinic|912,918
where|919,924
she|925,928
was|929,932
found|933,938
to|939,941
be|942,944
in|945,947
Afib|948,952
w|953,954
/|954,955
RVR|956,959
,|959,960
rate|961,965
around|966,972
<EOL>|973,974
110|974,977
-|977,978
120|978,981
.|981,982
She|983,986
has|987,990
a|991,992
history|993,1000
of|1001,1003
afib|1004,1008
.|1008,1009
He|1010,1012
referred|1013,1021
her|1022,1025
to|1026,1028
the|1029,1032
ED|1033,1035
<EOL>|1036,1037
for|1037,1040
persistent|1041,1051
SOB|1052,1055
and|1056,1059
afib|1060,1064
with|1065,1069
RVR|1070,1073
.|1073,1074
She|1075,1078
states|1079,1085
she|1086,1089
been|1090,1094
<EOL>|1095,1096
compliant|1096,1105
with|1106,1110
nebs|1111,1115
and|1116,1119
steroid|1120,1127
/|1127,1128
azithro|1128,1135
regimen|1136,1143
.|1143,1144
She|1145,1148
denies|1149,1155
any|1156,1159
<EOL>|1160,1161
_|1161,1162
_|1162,1163
_|1163,1164
edema|1165,1170
,|1170,1171
orthopnea|1172,1181
.|1181,1182
She|1183,1186
denies|1187,1193
recent|1194,1200
travel|1201,1207
,|1207,1208
surgeries|1209,1218
.|1218,1219
She|1220,1223
<EOL>|1224,1225
had|1225,1228
an|1229,1231
episode|1232,1239
of|1240,1242
chest|1243,1248
tightness|1249,1258
this|1259,1263
AM|1264,1266
that|1267,1271
felt|1272,1276
like|1277,1281
her|1282,1285
<EOL>|1286,1287
COPD|1287,1291
flares|1292,1298
.|1298,1299
Denies|1300,1306
fevers|1307,1313
or|1314,1316
coughing|1317,1325
or|1326,1328
production|1329,1339
of|1340,1342
sputum|1343,1349
,|1349,1350
<EOL>|1351,1352
hemomptysis|1352,1363
.|1363,1364
<EOL>|1366,1367
<EOL>|1368,1369
Past|1369,1373
Medical|1374,1381
History|1382,1389
:|1389,1390
<EOL>|1390,1391
ASTHMA|1391,1397
/|1397,1398
COPD|1398,1402
<EOL>|1404,1405
ATYPICAL|1406,1414
CHEST|1415,1420
PAIN|1421,1425
<EOL>|1427,1428
CERVICAL|1429,1437
RADICULITIS|1438,1449
<EOL>|1451,1452
CERVICAL|1453,1461
SPONDYLOSIS|1462,1473
<EOL>|1475,1476
CORONARY|1477,1485
ARTERY|1486,1492
DISEASE|1493,1500
<EOL>|1502,1503
HEADACHE|1504,1512
<EOL>|1514,1515
HIP|1516,1519
REPLACEMENT|1520,1531
<EOL>|1533,1534
HYPERLIPIDEMIA|1535,1549
<EOL>|1551,1552
HYPERTENSION|1553,1565
<EOL>|1567,1568
OSTEOARTHRITIS|1569,1583
<EOL>|1585,1586
HERPES|1587,1593
ZOSTER|1594,1600
<EOL>|1602,1603
ATRIAL|1604,1610
FIBRILLATION|1611,1623
<EOL>|1625,1626
ANXIETY|1627,1634
<EOL>|1636,1637
GASTROINTESTINAL|1638,1654
BLEEDING|1655,1663
<EOL>|1665,1666
OSTEOARTHRITIS|1667,1681
<EOL>|1683,1684
ATHEROSCLEROTIC|1685,1700
CARDIOVASCULAR|1701,1715
DISEASE|1716,1723
<EOL>|1725,1726
PERIPHERAL|1727,1737
VASCULAR|1738,1746
DISEASE|1747,1754
<EOL>|1754,1755
<EOL>|1756,1757
Social|1757,1763
History|1764,1771
:|1771,1772
<EOL>|1772,1773
_|1773,1774
_|1774,1775
_|1775,1776
<EOL>|1776,1777
Family|1777,1783
History|1784,1791
:|1791,1792
<EOL>|1792,1793
Mother|1793,1799
:|1799,1800
_|1801,1802
_|1802,1803
_|1803,1804
,|1804,1805
HTN|1806,1809
<EOL>|1811,1812
Father|1812,1818
:|1818,1819
_|1820,1821
_|1821,1822
_|1822,1823
CA|1824,1826
<EOL>|1828,1829
Brother|1829,1836
:|1836,1837
CA|1838,1840
?|1840,1841
<EOL>|1843,1844
Brother|1844,1851
:|1851,1852
_|1853,1854
_|1854,1855
_|1855,1856
<EOL>|1857,1858
<EOL>|1859,1860
Physical|1860,1868
_|1869,1870
_|1870,1871
_|1871,1872
:|1872,1873
<EOL>|1873,1874
ADMISSION|1874,1883
PHYSICAL|1884,1892
EXAM|1893,1897
:|1897,1898
<EOL>|1898,1899
VS|1899,1901
:|1901,1902
98.14|1903,1908
154|1909,1912
/|1912,1913
74|1913,1915
71|1916,1918
24|1919,1921
98|1922,1924
%|1924,1925
2L|1926,1928
<EOL>|1930,1931
GENERAL|1932,1939
:|1939,1940
Well|1941,1945
appearing|1946,1955
,|1955,1956
NAD|1957,1960
,|1960,1961
no|1962,1964
accessory|1965,1974
muscle|1975,1981
use|1982,1985
.|1985,1986
<EOL>|1988,1989
HEENT|1990,1995
:|1995,1996
NCAT|1997,2001
.|2001,2002
Sclera|2003,2009
anicteric|2010,2019
.|2019,2020
PERRL|2021,2026
,|2026,2027
EOMI|2028,2032
.|2032,2033
<EOL>|2035,2036
NECK|2037,2041
:|2041,2042
No|2043,2045
JVD|2046,2049
<EOL>|2051,2052
CARDIAC|2053,2060
:|2060,2061
Irregular|2062,2071
rhythm|2072,2078
,|2078,2079
normal|2080,2086
rate|2087,2091
.|2091,2092
Normal|2093,2099
S1|2100,2102
,|2102,2103
S2|2104,2106
.|2106,2107
No|2108,2110
<EOL>|2111,2112
murmurs|2112,2119
/|2119,2120
rubs|2120,2124
/|2124,2125
gallops|2125,2132
.|2132,2133
<EOL>|2135,2136
LUNGS|2137,2142
:|2142,2143
Moving|2144,2150
air|2151,2154
well|2155,2159
bilaterally|2160,2171
.|2171,2172
Trace|2173,2178
inspiratory|2179,2190
wheezing|2191,2199
<EOL>|2200,2201
and|2201,2204
louder|2205,2211
expiratory|2212,2222
wheezing|2223,2231
in|2232,2234
all|2235,2238
lung|2239,2243
fields|2244,2250
.|2250,2251
No|2252,2254
<EOL>|2255,2256
crackles|2256,2264
/|2264,2265
rhonchi|2265,2272
.|2272,2273
<EOL>|2275,2276
ABDOMEN|2277,2284
:|2284,2285
Soft|2286,2290
,|2290,2291
NTND|2292,2296
.|2296,2297
No|2298,2300
HSM|2301,2304
or|2305,2307
tenderness|2308,2318
.|2318,2319
<EOL>|2321,2322
EXTREMITIES|2323,2334
:|2334,2335
No|2336,2338
c|2339,2340
/|2340,2341
c|2341,2342
/|2342,2343
e|2343,2344
.|2344,2345
No|2346,2348
femoral|2349,2356
bruits|2357,2363
.|2363,2364
<EOL>|2366,2367
<EOL>|2367,2368
DISCHARGE|2368,2377
PHYSICAL|2378,2386
EXAM|2387,2391
:|2391,2392
<EOL>|2392,2393
VS|2393,2395
:|2395,2396
Tm|2397,2399
98.8|2400,2404
Tc|2405,2407
98.4|2408,2412
_|2413,2414
_|2414,2415
_|2415,2416
RA|2417,2419
<EOL>|2419,2420
GENERAL|2420,2427
:|2427,2428
NAD|2429,2432
<EOL>|2432,2433
HEENT|2433,2438
:|2438,2439
NCAT|2440,2444
.|2444,2445
Sclera|2446,2452
anicteric|2453,2462
.|2462,2463
Conjunctivae|2464,2476
noninjected|2477,2488
.|2488,2489
OM|2490,2492
<EOL>|2493,2494
clear|2494,2499
.|2499,2500
<EOL>|2500,2501
NECK|2501,2505
:|2505,2506
No|2507,2509
JVD|2510,2513
<EOL>|2515,2516
CARDIAC|2516,2523
:|2523,2524
RRR|2525,2528
.|2528,2529
Normal|2530,2536
S1|2537,2539
,|2539,2540
S2|2541,2543
.|2543,2544
No|2545,2547
murmurs|2548,2555
/|2555,2556
rubs|2556,2560
/|2560,2561
gallops|2561,2568
.|2568,2569
<EOL>|2571,2572
LUNGS|2572,2577
:|2577,2578
Mildly|2579,2585
reduced|2586,2593
air|2594,2597
movement|2598,2606
,|2606,2607
significant|2608,2619
wheezing|2620,2628
<EOL>|2629,2630
bilaterally|2630,2641
,|2641,2642
+|2643,2644
rhonchi|2644,2651
,|2651,2652
no|2653,2655
crackles|2656,2664
<EOL>|2666,2667
ABDOMEN|2667,2674
:|2674,2675
Soft|2676,2680
,|2680,2681
NTND|2682,2686
.|2686,2687
No|2688,2690
HSM|2691,2694
or|2695,2697
tenderness|2698,2708
.|2708,2709
<EOL>|2711,2712
EXTREMITIES|2712,2723
:|2723,2724
No|2725,2727
c|2728,2729
/|2729,2730
c|2730,2731
/|2731,2732
e|2732,2733
.|2733,2734
<EOL>|2735,2736
<EOL>|2737,2738
Pertinent|2738,2747
Results|2748,2755
:|2755,2756
<EOL>|2756,2757
ADMISSION|2757,2766
LABS|2767,2771
:|2771,2772
<EOL>|2772,2773
_|2773,2774
_|2774,2775
_|2775,2776
03|2777,2779
:|2779,2780
38PM|2780,2784
BLOOD|2785,2790
WBC|2791,2794
-|2794,2795
7.2|2795,2798
RBC|2799,2802
-|2802,2803
4.06|2803,2807
Hgb|2808,2811
-|2811,2812
9|2812,2813
.|2813,2814
4|2814,2815
*|2815,2816
Hct|2817,2820
-|2820,2821
31|2821,2823
.|2823,2824
4|2824,2825
*|2825,2826
<EOL>|2827,2828
MCV|2828,2831
-|2831,2832
77|2832,2834
*|2834,2835
MCH|2836,2839
-|2839,2840
23|2840,2842
.|2842,2843
2|2843,2844
*|2844,2845
MCHC|2846,2850
-|2850,2851
29|2851,2853
.|2853,2854
9|2854,2855
*|2855,2856
RDW|2857,2860
-|2860,2861
16|2861,2863
.|2863,2864
9|2864,2865
*|2865,2866
RDWSD|2867,2872
-|2872,2873
47|2873,2875
.|2875,2876
2|2876,2877
*|2877,2878
Plt|2879,2882
_|2883,2884
_|2884,2885
_|2885,2886
<EOL>|2886,2887
_|2887,2888
_|2888,2889
_|2889,2890
03|2891,2893
:|2893,2894
38PM|2894,2898
BLOOD|2899,2904
Neuts|2905,2910
-|2910,2911
93|2911,2913
.|2913,2914
8|2914,2915
*|2915,2916
Lymphs|2917,2923
-|2923,2924
4|2924,2925
.|2925,2926
2|2926,2927
*|2927,2928
Monos|2929,2934
-|2934,2935
1|2935,2936
.|2936,2937
3|2937,2938
*|2938,2939
<EOL>|2940,2941
Eos|2941,2944
-|2944,2945
0|2945,2946
.|2946,2947
0|2947,2948
*|2948,2949
Baso|2950,2954
-|2954,2955
0.0|2955,2958
Im|2959,2961
_|2962,2963
_|2963,2964
_|2964,2965
AbsNeut|2966,2973
-|2973,2974
6|2974,2975
.|2975,2976
74|2976,2978
*|2978,2979
#|2979,2980
AbsLymp|2981,2988
-|2988,2989
0|2989,2990
.|2990,2991
30|2991,2993
*|2993,2994
<EOL>|2995,2996
AbsMono|2996,3003
-|3003,3004
0|3004,3005
.|3005,3006
09|3006,3008
*|3008,3009
AbsEos|3010,3016
-|3016,3017
0|3017,3018
.|3018,3019
00|3019,3021
*|3021,3022
AbsBaso|3023,3030
-|3030,3031
0|3031,3032
.|3032,3033
00|3033,3035
*|3035,3036
<EOL>|3036,3037
_|3037,3038
_|3038,3039
_|3039,3040
03|3041,3043
:|3043,3044
38PM|3044,3048
BLOOD|3049,3054
_|3055,3056
_|3056,3057
_|3057,3058
PTT|3059,3062
-|3062,3063
30.3|3063,3067
_|3068,3069
_|3069,3070
_|3070,3071
<EOL>|3071,3072
_|3072,3073
_|3073,3074
_|3074,3075
03|3076,3078
:|3078,3079
38PM|3079,3083
BLOOD|3084,3089
Glucose|3090,3097
-|3097,3098
141|3098,3101
*|3101,3102
UreaN|3103,3108
-|3108,3109
20|3109,3111
Creat|3112,3117
-|3117,3118
1.0|3118,3121
Na|3122,3124
-|3124,3125
133|3125,3128
<EOL>|3129,3130
K|3130,3131
-|3131,3132
3.8|3132,3135
Cl|3136,3138
-|3138,3139
93|3139,3141
*|3141,3142
HCO3|3143,3147
-|3147,3148
30|3148,3150
AnGap|3151,3156
-|3156,3157
14|3157,3159
<EOL>|3159,3160
_|3160,3161
_|3161,3162
_|3162,3163
03|3164,3166
:|3166,3167
38PM|3167,3171
BLOOD|3172,3177
Calcium|3178,3185
-|3185,3186
9.9|3186,3189
Phos|3190,3194
-|3194,3195
2.8|3195,3198
Mg|3199,3201
-|3201,3202
2.1|3202,3205
<EOL>|3205,3206
<EOL>|3206,3207
PERTINENT|3207,3216
LABS|3217,3221
:|3221,3222
<EOL>|3222,3223
_|3223,3224
_|3224,3225
_|3225,3226
03|3227,3229
:|3229,3230
58PM|3230,3234
BLOOD|3235,3240
cTropnT|3241,3248
-|3248,3249
<|3249,3250
0|3250,3251
.|3251,3252
01|3252,3254
<EOL>|3254,3255
_|3255,3256
_|3256,3257
_|3257,3258
06|3259,3261
:|3261,3262
50AM|3262,3266
BLOOD|3267,3272
CK|3273,3275
-|3275,3276
MB|3276,3278
-|3278,3279
4|3279,3280
cTropnT|3281,3288
-|3288,3289
<|3289,3290
0|3290,3291
.|3291,3292
01|3292,3294
<EOL>|3294,3295
_|3295,3296
_|3296,3297
_|3297,3298
06|3299,3301
:|3301,3302
50AM|3302,3306
BLOOD|3307,3312
calTIBC|3313,3320
-|3320,3321
398|3321,3324
Ferritn|3325,3332
-|3332,3333
16|3333,3335
TRF|3336,3339
-|3339,3340
306|3340,3343
<EOL>|3343,3344
_|3344,3345
_|3345,3346
_|3346,3347
06|3348,3350
:|3350,3351
50AM|3351,3355
BLOOD|3356,3361
TSH|3362,3365
-|3365,3366
4|3366,3367
.|3367,3368
5|3368,3369
*|3369,3370
<EOL>|3370,3371
_|3371,3372
_|3372,3373
_|3373,3374
09|3375,3377
:|3377,3378
31AM|3378,3382
BLOOD|3383,3388
_|3389,3390
_|3390,3391
_|3391,3392
pO2|3393,3396
-|3396,3397
73|3397,3399
*|3399,3400
pCO2|3401,3405
-|3405,3406
58|3406,3408
*|3408,3409
pH|3410,3412
-|3412,3413
7.35|3413,3417
<EOL>|3418,3419
calTCO2|3419,3426
-|3426,3427
33|3427,3429
*|3429,3430
Base|3431,3435
XS|3436,3438
-|3438,3439
3|3439,3440
<EOL>|3445,3446
_|3446,3447
_|3447,3448
_|3448,3449
07|3450,3452
:|3452,3453
15AM|3453,3457
BLOOD|3458,3463
T4|3464,3466
,|3466,3467
FREE|3468,3472
,|3472,3473
DIRECT|3474,3480
DIALYSIS|3481,3489
-|3489,3490
Test|3490,3494
<EOL>|3496,3497
<EOL>|3497,3498
DISCHARGE|3498,3507
LABS|3508,3512
:|3512,3513
<EOL>|3517,3518
_|3518,3519
_|3519,3520
_|3520,3521
05|3522,3524
:|3524,3525
30AM|3525,3529
BLOOD|3530,3535
WBC|3536,3539
-|3539,3540
13|3540,3542
.|3542,3543
2|3543,3544
*|3544,3545
RBC|3546,3549
-|3549,3550
3|3550,3551
.|3551,3552
97|3552,3554
Hgb|3555,3558
-|3558,3559
9|3559,3560
.|3560,3561
0|3561,3562
*|3562,3563
Hct|3564,3567
-|3567,3568
31|3568,3570
.|3570,3571
1|3571,3572
*|3572,3573
<EOL>|3574,3575
MCV|3575,3578
-|3578,3579
78|3579,3581
*|3581,3582
MCH|3583,3586
-|3586,3587
22|3587,3589
.|3589,3590
7|3590,3591
*|3591,3592
MCHC|3593,3597
-|3597,3598
28|3598,3600
.|3600,3601
9|3601,3602
*|3602,3603
RDW|3604,3607
-|3607,3608
17|3608,3610
.|3610,3611
4|3611,3612
*|3612,3613
RDWSD|3614,3619
-|3619,3620
48|3620,3622
.|3622,3623
7|3623,3624
*|3624,3625
Plt|3626,3629
_|3630,3631
_|3631,3632
_|3632,3633
<EOL>|3633,3634
_|3634,3635
_|3635,3636
_|3636,3637
05|3638,3640
:|3640,3641
30AM|3641,3645
BLOOD|3646,3651
Glucose|3652,3659
-|3659,3660
85|3660,3662
UreaN|3663,3668
-|3668,3669
23|3669,3671
*|3671,3672
Creat|3673,3678
-|3678,3679
0.9|3679,3682
Na|3683,3685
-|3685,3686
136|3686,3689
<EOL>|3690,3691
K|3691,3692
-|3692,3693
3.9|3693,3696
Cl|3697,3699
-|3699,3700
95|3700,3702
*|3702,3703
HCO3|3704,3708
-|3708,3709
30|3709,3711
AnGap|3712,3717
-|3717,3718
15|3718,3720
<EOL>|3720,3721
_|3721,3722
_|3722,3723
_|3723,3724
06|3725,3727
:|3727,3728
30AM|3728,3732
BLOOD|3733,3738
Calcium|3739,3746
-|3746,3747
9.7|3747,3750
Phos|3751,3755
-|3755,3756
3.0|3756,3759
Mg|3760,3762
-|3762,3763
2.0|3763,3766
<EOL>|3766,3767
<EOL>|3767,3768
IMAGING|3768,3775
:|3775,3776
<EOL>|3776,3777
_|3777,3778
_|3778,3779
_|3779,3780
Chest|3781,3786
X|3787,3788
ray|3789,3792
:|3792,3793
Relative|3794,3802
increase|3803,3811
in|3812,3814
opacity|3815,3822
over|3823,3827
the|3828,3831
lung|3832,3836
<EOL>|3837,3838
bases|3838,3843
bilaterally|3844,3855
felt|3856,3860
due|3861,3864
to|3865,3867
overlying|3868,3877
soft|3878,3882
tissue|3883,3889
rather|3890,3896
than|3897,3901
<EOL>|3902,3903
consolidation|3903,3916
.|3916,3917
Lateral|3919,3926
view|3927,3931
may|3932,3935
be|3936,3938
helpful|3939,3946
for|3947,3950
confirmation|3951,3963
.|3963,3964
<EOL>|3964,3965
<EOL>|3965,3966
_|3966,3967
_|3967,3968
_|3968,3969
Chest|3970,3975
X|3976,3977
ray|3978,3981
:|3981,3982
There|3983,3988
is|3989,3991
hyperinflation|3992,4006
.|4006,4007
There|4009,4014
is|4015,4017
no|4018,4020
<EOL>|4021,4022
pneumothorax|4022,4034
,|4034,4035
effusion|4036,4044
,|4044,4045
consolidation|4046,4059
or|4060,4062
CHF|4063,4066
.|4066,4067
There|4069,4074
is|4075,4077
probable|4078,4086
<EOL>|4087,4088
osteopenia|4088,4098
.|4098,4099
<EOL>|4099,4100
<EOL>|4101,4102
Brief|4102,4107
Hospital|4108,4116
Course|4117,4123
:|4123,4124
<EOL>|4124,4125
_|4125,4126
_|4126,4127
_|4127,4128
is|4129,4131
a|4132,4133
_|4134,4135
_|4135,4136
_|4136,4137
with|4138,4142
a|4143,4144
history|4145,4152
of|4153,4155
CAD|4156,4159
,|4159,4160
PVD|4161,4164
,|4164,4165
and|4166,4169
<EOL>|4170,4171
COPD|4171,4175
and|4176,4179
history|4180,4187
of|4188,4190
recurrent|4191,4200
chest|4201,4206
pain|4207,4211
who|4212,4215
presented|4216,4225
with|4226,4230
afib|4231,4235
<EOL>|4236,4237
with|4237,4241
RVR|4242,4245
and|4246,4249
COPD|4250,4254
exacerbation|4255,4267
.|4267,4268
<EOL>|4269,4270
<EOL>|4272,4273
ACUTE|4273,4278
PROBLEMS|4279,4287
:|4287,4288
<EOL>|4288,4289
<EOL>|4289,4290
#|4290,4291
COPD|4291,4295
exacerbation|4296,4308
:|4308,4309
Ms.|4310,4313
_|4314,4315
_|4315,4316
_|4316,4317
had|4318,4321
had|4322,4325
two|4326,4329
recent|4330,4336
ED|4337,4339
visits|4340,4346
<EOL>|4347,4348
for|4348,4351
COPD|4352,4356
exacerbation|4357,4369
,|4369,4370
most|4371,4375
recently|4376,4384
_|4385,4386
_|4386,4387
_|4387,4388
when|4389,4393
she|4394,4397
was|4398,4401
started|4402,4409
<EOL>|4410,4411
on|4411,4413
prednisone|4414,4424
60|4425,4427
mg|4428,4430
.|4430,4431
She|4432,4435
presented|4436,4445
to|4446,4448
her|4449,4452
PCP|4453,4456
's|4456,4458
office|4459,4465
with|4466,4470
<EOL>|4471,4472
worsening|4472,4481
dyspnea|4482,4489
despite|4490,4497
this|4498,4502
therapy|4503,4510
and|4511,4514
was|4515,4518
also|4519,4523
complaining|4524,4535
<EOL>|4536,4537
of|4537,4539
nasal|4540,4545
congestion|4546,4556
,|4556,4557
suggesting|4558,4568
a|4569,4570
viral|4571,4576
URI|4577,4580
trigger|4581,4588
.|4588,4589
In|4590,4592
clinic|4593,4599
<EOL>|4600,4601
she|4601,4604
was|4605,4608
also|4609,4613
noted|4614,4619
to|4620,4622
be|4623,4625
in|4626,4628
afib|4629,4633
with|4634,4638
RVR|4639,4642
so|4643,4645
was|4646,4649
referred|4650,4658
to|4659,4661
the|4662,4665
<EOL>|4666,4667
ED|4667,4669
where|4670,4675
she|4676,4679
was|4680,4683
admitted|4684,4692
after|4693,4698
control|4699,4706
of|4707,4709
her|4710,4713
heart|4714,4719
rate|4720,4724
(|4725,4726
see|4726,4729
<EOL>|4730,4731
below|4731,4736
)|4736,4737
.|4737,4738
On|4739,4741
admission|4742,4751
to|4752,4754
the|4755,4758
floor|4759,4764
,|4764,4765
she|4766,4769
was|4770,4773
noted|4774,4779
to|4780,4782
have|4783,4787
<EOL>|4788,4789
wheezing|4789,4797
,|4797,4798
increased|4799,4808
work|4809,4813
of|4814,4816
breathing|4817,4826
,|4826,4827
and|4828,4831
poor|4832,4836
air|4837,4840
movement|4841,4849
.|4849,4850
<EOL>|4851,4852
She|4852,4855
was|4856,4859
treated|4860,4867
with|4868,4872
125|4873,4876
mg|4877,4879
solumedrol|4880,4890
and|4891,4894
maintained|4895,4905
on|4906,4908
60|4909,4911
mg|4912,4914
<EOL>|4915,4916
PO|4916,4918
prednisone|4919,4929
daily|4930,4935
.|4935,4936
Her|4937,4940
home|4941,4945
theophylline|4946,4958
was|4959,4962
decreased|4963,4972
from|4973,4977
<EOL>|4978,4979
400|4979,4982
mg|4983,4985
BID|4986,4989
to|4990,4992
_|4993,4994
_|4994,4995
_|4995,4996
mg|4997,4999
BID|5000,5003
due|5004,5007
to|5008,5010
concerns|5011,5019
it|5020,5022
was|5023,5026
contributing|5027,5039
to|5040,5042
<EOL>|5043,5044
her|5044,5047
tachyarrhythmia|5048,5063
.|5063,5064
She|5065,5068
was|5069,5072
placed|5073,5079
on|5080,5082
ipratropium|5083,5094
nebs|5095,5099
q6h|5100,5103
,|5103,5104
<EOL>|5105,5106
albuterol|5106,5115
nebs|5116,5120
q2h|5121,5124
,|5124,5125
and|5126,5129
fluticasone|5130,5141
-|5141,5142
salmeterol|5142,5152
.|5152,5153
Pulmonary|5154,5163
was|5164,5167
<EOL>|5168,5169
consulted|5169,5178
and|5179,5182
recommended|5183,5194
a|5195,5196
trial|5197,5202
of|5203,5205
diuresis|5206,5214
so|5215,5217
she|5218,5221
received|5222,5230
10|5231,5233
<EOL>|5234,5235
mg|5235,5237
IV|5238,5240
Lasix|5241,5246
as|5247,5249
well|5250,5254
.|5254,5255
Azithromycin|5256,5268
was|5269,5272
not|5273,5276
given|5277,5282
due|5283,5286
to|5287,5289
concerns|5290,5298
<EOL>|5299,5300
for|5300,5303
QT|5304,5306
prolongation|5307,5319
with|5320,5324
theophylline|5325,5337
and|5338,5341
amiodarone|5342,5352
(|5353,5354
QTc|5354,5357
was|5358,5361
<EOL>|5362,5363
460|5363,5366
)|5366,5367
.|5367,5368
She|5369,5372
was|5373,5376
started|5377,5384
on|5385,5387
a|5388,5389
5|5390,5391
day|5392,5395
course|5396,5402
of|5403,5405
ceftriaxone|5406,5417
instead|5418,5425
,|5425,5426
<EOL>|5427,5428
and|5428,5431
discharged|5432,5442
to|5443,5445
finish|5446,5452
the|5453,5456
course|5457,5463
with|5464,5468
cefpodoxime|5469,5480
.|5480,5481
She|5482,5485
was|5486,5489
<EOL>|5490,5491
discharged|5491,5501
with|5502,5506
a|5507,5508
prednisone|5509,5519
taper|5520,5525
(|5526,5527
10|5527,5529
mg|5530,5532
decrease|5533,5541
q3d|5542,5545
until|5546,5551
at|5552,5554
<EOL>|5555,5556
10|5556,5558
mg|5559,5561
,|5561,5562
then|5563,5567
stay|5568,5572
at|5573,5575
10|5576,5578
mg|5579,5581
until|5582,5587
pulm|5588,5592
follow|5593,5599
up|5600,5602
)|5602,5603
as|5604,5606
well|5607,5611
as|5612,5614
<EOL>|5615,5616
follow|5616,5622
up|5623,5625
with|5626,5630
pulmonary|5631,5640
rehab|5641,5646
and|5647,5650
a|5651,5652
pulmonologist|5653,5666
she|5667,5670
<EOL>|5671,5672
previously|5672,5682
followed|5683,5691
with|5692,5696
,|5696,5697
Dr.|5698,5701
_|5702,5703
_|5703,5704
_|5704,5705
.|5705,5706
She|5707,5710
was|5711,5714
also|5715,5719
discharged|5720,5730
on|5731,5733
<EOL>|5734,5735
2L|5735,5737
supplemental|5738,5750
O2|5751,5753
to|5754,5756
be|5757,5759
worn|5760,5764
at|5765,5767
all|5768,5771
times|5772,5777
.|5777,5778
<EOL>|5779,5780
<EOL>|5780,5781
#|5781,5782
Atrial|5782,5788
fibrillation|5789,5801
:|5801,5802
Ms.|5803,5806
_|5807,5808
_|5808,5809
_|5809,5810
has|5811,5814
known|5815,5820
atrial|5821,5827
<EOL>|5828,5829
fibrillation|5829,5841
for|5842,5845
which|5846,5851
she|5852,5855
was|5856,5859
on|5860,5862
amiodarone|5863,5873
and|5874,5877
apixaban|5878,5886
but|5887,5890
<EOL>|5891,5892
was|5892,5895
found|5896,5901
to|5902,5904
have|5905,5909
HR|5910,5912
in|5913,5915
the|5916,5919
120s|5920,5924
in|5925,5927
her|5928,5931
PCP|5932,5935
's|5935,5937
office|5938,5944
,|5944,5945
prompting|5946,5955
<EOL>|5956,5957
her|5957,5960
referral|5961,5969
to|5970,5972
the|5973,5976
ED|5977,5979
.|5979,5980
Her|5981,5984
COPD|5985,5989
exacerbation|5990,6002
was|6003,6006
the|6007,6010
likely|6011,6017
<EOL>|6018,6019
precipitant|6019,6030
,|6030,6031
with|6032,6036
medications|6037,6048
also|6049,6053
possibly|6054,6062
contributing|6063,6075
,|6075,6076
<EOL>|6077,6078
particularly|6078,6090
theophylline|6091,6103
.|6103,6104
She|6105,6108
was|6109,6112
started|6113,6120
on|6121,6123
a|6124,6125
diltiazem|6126,6135
gtt|6136,6139
in|6140,6142
<EOL>|6143,6144
the|6144,6147
ED|6148,6150
to|6151,6153
control|6154,6161
her|6162,6165
rates|6166,6171
than|6172,6176
transitioned|6177,6189
to|6190,6192
diltiazem|6193,6202
90|6203,6205
mg|6206,6208
<EOL>|6209,6210
q6h|6210,6213
.|6213,6214
After|6215,6220
arrival|6221,6228
to|6229,6231
the|6232,6235
floor|6236,6241
,|6241,6242
her|6243,6246
rates|6247,6252
remained|6253,6261
controlled|6262,6272
.|6272,6273
<EOL>|6274,6275
Her|6275,6278
amiodarone|6279,6289
and|6290,6293
apixaban|6294,6302
were|6303,6307
continued|6308,6317
.|6317,6318
Her|6319,6322
theophylline|6323,6335
was|6336,6339
<EOL>|6340,6341
decreased|6341,6350
to|6351,6353
200|6354,6357
mg|6358,6360
BID|6361,6364
from|6365,6369
400|6370,6373
mg|6374,6376
BID|6377,6380
.|6380,6381
<EOL>|6381,6382
<EOL>|6382,6383
#|6383,6384
Iron|6384,6388
deficiency|6389,6399
anemia|6400,6406
.|6406,6407
Patient|6408,6415
was|6416,6419
found|6420,6425
to|6426,6428
have|6429,6433
microcytic|6434,6444
<EOL>|6445,6446
anemia|6446,6452
with|6453,6457
low|6458,6461
iron|6462,6466
and|6467,6470
ferritin|6471,6479
.|6479,6480
She|6481,6484
was|6485,6488
started|6489,6496
on|6497,6499
IV|6500,6502
iron|6503,6507
<EOL>|6508,6509
125|6509,6512
mg|6513,6515
ferric|6516,6522
gluconate|6523,6532
x4|6533,6535
doses|6536,6541
and|6542,6545
wasdischarged|6546,6559
on|6560,6562
PO|6563,6565
iron|6566,6570
<EOL>|6571,6572
with|6572,6576
a|6577,6578
bowel|6579,6584
regimen|6585,6592
.|6592,6593
Her|6594,6597
H|6598,6599
/|6599,6600
H|6600,6601
was|6602,6605
stable|6606,6612
throughout|6613,6623
the|6624,6627
<EOL>|6628,6629
hospitalized|6629,6641
;|6641,6642
there|6643,6648
was|6649,6652
no|6653,6655
evidence|6656,6664
of|6665,6667
bleeding|6668,6676
.|6676,6677
<EOL>|6677,6678
<EOL>|6678,6679
Transitional|6679,6691
issues|6692,6698
:|6698,6699
<EOL>|6699,6700
-|6700,6701
patient|6702,6709
discharged|6710,6720
on|6721,6723
prednisone|6724,6734
taper|6735,6740
:|6740,6741
decrease|6742,6750
by|6751,6753
10|6754,6756
mg|6757,6759
<EOL>|6760,6761
every|6761,6766
3|6767,6768
days|6769,6773
until|6774,6779
at|6780,6782
10|6783,6785
mg|6786,6788
,|6788,6789
then|6790,6794
keep|6795,6799
at|6800,6802
10|6803,6805
mg|6806,6808
until|6809,6814
seen|6815,6819
by|6820,6822
<EOL>|6823,6824
pulmonology|6824,6835
<EOL>|6835,6836
-|6836,6837
patient|6838,6845
discharged|6846,6856
with|6857,6861
plan|6862,6866
to|6867,6869
follow|6870,6876
up|6877,6879
with|6880,6884
pulmonology|6885,6896
and|6897,6900
<EOL>|6901,6902
pulmonary|6902,6911
rehab|6912,6917
.|6917,6918
Can|6919,6922
call|6923,6927
_|6928,6929
_|6929,6930
_|6930,6931
to|6932,6934
schedule|6935,6943
appointment|6944,6955
<EOL>|6956,6957
with|6957,6961
pulmonary|6962,6971
rehab|6972,6977
.|6977,6978
<EOL>|6978,6979
-|6979,6980
patient|6981,6988
discharged|6989,6999
on|7000,7002
with|7003,7007
2|7008,7009
days|7010,7014
of|7015,7017
cefpodoxime|7018,7029
to|7030,7032
complete|7033,7041
5|7042,7043
<EOL>|7044,7045
day|7045,7048
course|7049,7055
of|7056,7058
antibiotics|7059,7070
for|7071,7074
severe|7075,7081
COPD|7082,7086
exacerbation|7087,7099
<EOL>|7099,7100
-|7100,7101
patient|7102,7109
discharged|7110,7120
with|7121,7125
O2|7126,7128
concentrator|7129,7141
for|7142,7145
continuous|7146,7156
home|7157,7161
O2|7162,7164
<EOL>|7164,7165
-|7165,7166
patient|7167,7174
's|7174,7176
theophylline|7177,7189
decreased|7190,7199
from|7200,7204
300|7205,7208
mg|7209,7211
BID|7212,7215
to|7216,7218
_|7219,7220
_|7220,7221
_|7221,7222
mg|7223,7225
BID|7226,7229
<EOL>|7230,7231
due|7231,7234
to|7235,7237
her|7238,7241
afib|7242,7246
with|7247,7251
RVR|7252,7255
;|7255,7256
may|7257,7260
want|7261,7265
to|7266,7268
consider|7269,7277
further|7278,7285
<EOL>|7286,7287
theophylline|7287,7299
wean|7300,7304
,|7304,7305
and|7306,7309
addition|7310,7318
of|7319,7321
azithromycin|7322,7334
(|7335,7336
if|7336,7338
QTc|7339,7342
is|7343,7345
<EOL>|7346,7347
decreased|7347,7356
as|7357,7359
patient|7360,7367
also|7368,7372
on|7373,7375
amiodarone|7376,7386
)|7386,7387
,|7387,7388
and|7389,7392
/|7392,7393
or|7393,7395
roflumilast|7396,7407
<EOL>|7408,7409
therapy|7409,7416
<EOL>|7416,7417
-|7417,7418
patient|7419,7426
found|7427,7432
to|7433,7435
be|7436,7438
iron|7439,7443
deficient|7444,7453
,|7453,7454
started|7455,7462
on|7463,7465
IV|7466,7468
iron|7469,7473
<EOL>|7474,7475
repletion|7475,7484
,|7484,7485
discharged|7486,7496
on|7497,7499
PO|7500,7502
iron|7503,7507
<EOL>|7507,7508
-|7508,7509
patient|7510,7517
found|7518,7523
to|7524,7526
have|7527,7531
elevated|7532,7540
TSH|7541,7544
,|7544,7545
please|7546,7552
follow|7553,7559
up|7560,7562
free|7563,7567
T4|7568,7570
<EOL>|7571,7572
which|7572,7577
was|7578,7581
pending|7582,7589
on|7590,7592
discharge|7593,7602
<EOL>|7602,7603
-|7603,7604
Code|7605,7609
:|7609,7610
full|7611,7615
<EOL>|7615,7616
-|7616,7617
Emergency|7618,7627
Contact|7628,7635
_|7636,7637
_|7637,7638
_|7638,7639
(|7640,7641
Husband|7641,7648
)|7648,7649
_|7650,7651
_|7651,7652
_|7652,7653
<EOL>|7654,7655
Daughter|7655,7663
_|7664,7665
_|7665,7666
_|7666,7667
:|7667,7668
_|7669,7670
_|7670,7671
_|7671,7672
<EOL>|7673,7674
<EOL>|7675,7676
_|7676,7677
_|7677,7678
_|7678,7679
on|7680,7682
Admission|7683,7692
:|7692,7693
<EOL>|7693,7694
The|7694,7697
Preadmission|7698,7710
Medication|7711,7721
list|7722,7726
is|7727,7729
accurate|7730,7738
and|7739,7742
complete|7743,7751
.|7751,7752
<EOL>|7752,7753
1.|7753,7755
Acetaminophen|7756,7769
650|7770,7773
mg|7774,7776
PO|7777,7779
Q6H|7780,7783
:|7783,7784
PRN|7784,7787
pain|7788,7792
<EOL>|7793,7794
2.|7794,7796
Apixaban|7797,7805
5|7806,7807
mg|7808,7810
PO|7811,7813
BID|7814,7817
<EOL>|7818,7819
3.|7819,7821
Albuterol|7822,7831
0.083|7832,7837
%|7837,7838
Neb|7839,7842
Soln|7843,7847
1|7848,7849
NEB|7850,7853
IH|7854,7856
Q6H|7857,7860
:|7860,7861
PRN|7861,7864
shortness|7865,7874
of|7875,7877
<EOL>|7878,7879
breath|7879,7885
<EOL>|7886,7887
4.|7887,7889
Amiodarone|7890,7900
200|7901,7904
mg|7905,7907
PO|7908,7910
DAILY|7911,7916
<EOL>|7917,7918
5.|7918,7920
Atorvastatin|7921,7933
10|7934,7936
mg|7937,7939
PO|7940,7942
QPM|7943,7946
<EOL>|7947,7948
6.|7948,7950
Artificial|7951,7961
Tears|7962,7967
_|7968,7969
_|7969,7970
_|7970,7971
DROP|7972,7976
BOTH|7977,7981
EYES|7982,7986
PRN|7987,7990
irritation|7991,8001
<EOL>|8002,8003
7.|8003,8005
Latanoprost|8006,8017
0.005|8018,8023
%|8023,8024
Ophth|8025,8030
.|8030,8031
Soln.|8032,8037
1|8038,8039
DROP|8040,8044
LEFT|8045,8049
EYE|8050,8053
QHS|8054,8057
<EOL>|8058,8059
8.|8059,8061
Diltiazem|8062,8071
Extended|8072,8080
-|8080,8081
Release|8081,8088
180|8089,8092
mg|8093,8095
PO|8096,8098
BID|8099,8102
<EOL>|8103,8104
9.|8104,8106
Fluticasone|8107,8118
Propionate|8119,8129
NASAL|8130,8135
1|8136,8137
SPRY|8138,8142
NU|8143,8145
BID|8146,8149
<EOL>|8150,8151
10.|8151,8154
Fluticasone|8155,8166
-|8166,8167
Salmeterol|8167,8177
Diskus|8178,8184
(|8185,8186
250|8186,8189
/|8189,8190
50|8190,8192
)|8192,8193
1|8195,8196
INH|8197,8200
IH|8201,8203
BID|8204,8207
<EOL>|8208,8209
11.|8209,8212
Hydrochlorothiazide|8213,8232
50|8233,8235
mg|8236,8238
PO|8239,8241
DAILY|8242,8247
<EOL>|8248,8249
12.|8249,8252
Isosorbide|8253,8263
Mononitrate|8264,8275
(|8276,8277
Extended|8277,8285
Release|8286,8293
)|8293,8294
240|8295,8298
mg|8299,8301
PO|8302,8304
DAILY|8305,8310
<EOL>|8311,8312
13.|8312,8315
Lorazepam|8316,8325
0.5|8326,8329
mg|8330,8332
PO|8333,8335
QHS|8336,8339
:|8339,8340
PRN|8340,8343
insomnia|8344,8352
<EOL>|8353,8354
14.|8354,8357
Theophylline|8358,8370
ER|8371,8373
300|8374,8377
mg|8378,8380
PO|8381,8383
BID|8384,8387
<EOL>|8388,8389
15.|8389,8392
Ranitidine|8393,8403
300|8404,8407
mg|8408,8410
PO|8411,8413
DAILY|8414,8419
<EOL>|8420,8421
16|8421,8423
.|8423,8424
Tiotropium|8425,8435
Bromide|8436,8443
1|8444,8445
CAP|8446,8449
IH|8450,8452
DAILY|8453,8458
<EOL>|8459,8460
17.|8460,8463
Multivitamins|8464,8477
W|8478,8479
/|8479,8480
minerals|8480,8488
1|8489,8490
TAB|8491,8494
PO|8495,8497
DAILY|8498,8503
<EOL>|8504,8505
18.|8505,8508
Aspirin|8509,8516
81|8517,8519
mg|8520,8522
PO|8523,8525
DAILY|8526,8531
<EOL>|8532,8533
19|8533,8535
.|8535,8536
Dorzolamide|8537,8548
2|8549,8550
%|8550,8551
Ophth|8552,8557
.|8557,8558
Soln.|8559,8564
1|8565,8566
DROP|8567,8571
BOTH|8572,8576
EYES|8577,8581
BID|8582,8585
<EOL>|8586,8587
<EOL>|8587,8588
<EOL>|8589,8590
Discharge|8590,8599
Medications|8600,8611
:|8611,8612
<EOL>|8612,8613
1.|8613,8615
Home|8616,8620
O2|8621,8623
<EOL>|8623,8624
2|8624,8625
Liters|8626,8632
continuous|8633,8643
nasal|8644,8649
cannula|8650,8657
with|8658,8662
exertion|8663,8671
<EOL>|8671,8672
Diagnosis|8672,8681
:|8681,8682
chronic|8683,8690
obstructive|8691,8702
pulmonary|8703,8712
disease|8713,8720
(|8721,8722
J44|8722,8725
.9|8725,8727
)|8727,8728
<EOL>|8728,8729
Length|8729,8735
of|8736,8738
Needs|8739,8744
:|8744,8745
ongoing|8746,8753
(|8754,8755
years|8755,8760
)|8760,8761
<EOL>|8761,8762
2.|8762,8764
Acetaminophen|8765,8778
650|8779,8782
mg|8783,8785
PO|8786,8788
Q6H|8789,8792
:|8792,8793
PRN|8793,8796
pain|8797,8801
<EOL>|8802,8803
3.|8803,8805
Amiodarone|8806,8816
200|8817,8820
mg|8821,8823
PO|8824,8826
DAILY|8827,8832
<EOL>|8833,8834
4.|8834,8836
Apixaban|8837,8845
5|8846,8847
mg|8848,8850
PO|8851,8853
BID|8854,8857
<EOL>|8858,8859
5.|8859,8861
Albuterol|8862,8871
0.083|8872,8877
%|8877,8878
Neb|8879,8882
Soln|8883,8887
1|8888,8889
NEB|8890,8893
IH|8894,8896
Q2H|8897,8900
:|8900,8901
PRN|8901,8904
shortness|8905,8914
of|8915,8917
<EOL>|8918,8919
breath|8919,8925
<EOL>|8926,8927
6.|8927,8929
Artificial|8930,8940
Tears|8941,8946
_|8947,8948
_|8948,8949
_|8949,8950
DROP|8951,8955
BOTH|8956,8960
EYES|8961,8965
PRN|8966,8969
irritation|8970,8980
<EOL>|8981,8982
7.|8982,8984
Aspirin|8985,8992
81|8993,8995
mg|8996,8998
PO|8999,9001
DAILY|9002,9007
<EOL>|9008,9009
8.|9009,9011
Atorvastatin|9012,9024
10|9025,9027
mg|9028,9030
PO|9031,9033
QPM|9034,9037
<EOL>|9038,9039
9.|9039,9041
Diltiazem|9042,9051
Extended|9052,9060
-|9060,9061
Release|9061,9068
180|9069,9072
mg|9073,9075
PO|9076,9078
BID|9079,9082
<EOL>|9083,9084
10.|9084,9087
Dorzolamide|9088,9099
2|9100,9101
%|9101,9102
Ophth|9103,9108
.|9108,9109
Soln.|9110,9115
1|9116,9117
DROP|9118,9122
BOTH|9123,9127
EYES|9128,9132
BID|9133,9136
<EOL>|9137,9138
11.|9138,9141
Fluticasone|9142,9153
Propionate|9154,9164
NASAL|9165,9170
1|9171,9172
SPRY|9173,9177
NU|9178,9180
BID|9181,9184
<EOL>|9185,9186
12.|9186,9189
Fluticasone|9190,9201
-|9201,9202
Salmeterol|9202,9212
Diskus|9213,9219
(|9220,9221
250|9221,9224
/|9224,9225
50|9225,9227
)|9227,9228
1|9230,9231
INH|9232,9235
IH|9236,9238
BID|9239,9242
<EOL>|9243,9244
13.|9244,9247
Hydrochlorothiazide|9248,9267
50|9268,9270
mg|9271,9273
PO|9274,9276
DAILY|9277,9282
<EOL>|9283,9284
14.|9284,9287
Isosorbide|9288,9298
Mononitrate|9299,9310
(|9311,9312
Extended|9312,9320
Release|9321,9328
)|9328,9329
240|9330,9333
mg|9334,9336
PO|9337,9339
DAILY|9340,9345
<EOL>|9346,9347
15.|9347,9350
Latanoprost|9351,9362
0.005|9363,9368
%|9368,9369
Ophth|9370,9375
.|9375,9376
Soln.|9377,9382
1|9383,9384
DROP|9385,9389
LEFT|9390,9394
EYE|9395,9398
QHS|9399,9402
<EOL>|9403,9404
16|9404,9406
.|9406,9407
Lorazepam|9408,9417
0.5|9418,9421
mg|9422,9424
PO|9425,9427
QHS|9428,9431
:|9431,9432
PRN|9432,9435
insomnia|9436,9444
<EOL>|9445,9446
17.|9446,9449
Multivitamins|9450,9463
W|9464,9465
/|9465,9466
minerals|9466,9474
1|9475,9476
TAB|9477,9480
PO|9481,9483
DAILY|9484,9489
<EOL>|9490,9491
18.|9491,9494
Ranitidine|9495,9505
300|9506,9509
mg|9510,9512
PO|9513,9515
DAILY|9516,9521
<EOL>|9522,9523
19|9523,9525
.|9525,9526
Tiotropium|9527,9537
Bromide|9538,9545
1|9546,9547
CAP|9548,9551
IH|9552,9554
DAILY|9555,9560
<EOL>|9561,9562
20|9562,9564
.|9564,9565
Theophylline|9566,9578
SR|9579,9581
200|9582,9585
mg|9586,9588
PO|9589,9591
BID|9592,9595
<EOL>|9596,9597
RX|9597,9599
*|9600,9601
theophylline|9601,9613
200|9614,9617
mg|9618,9620
1|9621,9622
tablet|9623,9629
(|9629,9630
s|9630,9631
)|9631,9632
by|9633,9635
mouth|9636,9641
twice|9642,9647
a|9648,9649
day|9650,9653
Disp|9654,9658
<EOL>|9659,9660
#|9660,9661
*|9661,9662
60|9662,9664
Tablet|9665,9671
Refills|9672,9679
:|9679,9680
*|9680,9681
0|9681,9682
<EOL>|9682,9683
21|9683,9685
.|9685,9686
Cefpodoxime|9687,9698
Proxetil|9699,9707
200|9708,9711
mg|9712,9714
PO|9715,9717
Q12H|9718,9722
Duration|9723,9731
:|9731,9732
2|9733,9734
Days|9735,9739
<EOL>|9740,9741
RX|9741,9743
*|9744,9745
cefpodoxime|9745,9756
200|9757,9760
mg|9761,9763
1|9764,9765
tablet|9766,9772
(|9772,9773
s|9773,9774
)|9774,9775
by|9776,9778
mouth|9779,9784
twice|9785,9790
a|9791,9792
day|9793,9796
Disp|9797,9801
#|9802,9803
*|9803,9804
4|9804,9805
<EOL>|9806,9807
Tablet|9807,9813
Refills|9814,9821
:|9821,9822
*|9822,9823
0|9823,9824
<EOL>|9824,9825
22.|9825,9828
Ferrous|9829,9836
Sulfate|9837,9844
325|9845,9848
mg|9849,9851
PO|9852,9854
DAILY|9855,9860
<EOL>|9861,9862
RX|9862,9864
*|9865,9866
ferrous|9866,9873
sulfate|9874,9881
325|9882,9885
mg|9886,9888
(|9889,9890
65|9890,9892
mg|9893,9895
iron|9896,9900
)|9900,9901
1|9902,9903
tablet|9904,9910
(|9910,9911
s|9911,9912
)|9912,9913
by|9914,9916
mouth|9917,9922
<EOL>|9923,9924
daily|9924,9929
Disp|9930,9934
#|9935,9936
*|9936,9937
30|9937,9939
Tablet|9940,9946
Refills|9947,9954
:|9954,9955
*|9955,9956
0|9956,9957
<EOL>|9957,9958
23|9958,9960
.|9960,9961
Docusate|9962,9970
Sodium|9971,9977
100|9978,9981
mg|9982,9984
PO|9985,9987
BID|9988,9991
<EOL>|9992,9993
RX|9993,9995
*|9996,9997
docusate|9997,10005
sodium|10006,10012
100|10013,10016
mg|10017,10019
1|10020,10021
capsule|10022,10029
(|10029,10030
s|10030,10031
)|10031,10032
by|10033,10035
mouth|10036,10041
twice|10042,10047
a|10048,10049
day|10050,10053
<EOL>|10054,10055
Disp|10055,10059
#|10060,10061
*|10061,10062
60|10062,10064
Capsule|10065,10072
Refills|10073,10080
:|10080,10081
*|10081,10082
0|10082,10083
<EOL>|10083,10084
24|10084,10086
.|10086,10087
Polyethylene|10088,10100
Glycol|10101,10107
17|10108,10110
g|10111,10112
PO|10113,10115
DAILY|10116,10121
<EOL>|10122,10123
RX|10123,10125
*|10126,10127
polyethylene|10127,10139
glycol|10140,10146
3350|10147,10151
17|10152,10154
gram|10155,10159
/|10159,10160
dose|10160,10164
1|10165,10166
powder|10167,10173
(|10173,10174
s|10174,10175
)|10175,10176
by|10177,10179
mouth|10180,10185
<EOL>|10186,10187
daily|10187,10192
Refills|10193,10200
:|10200,10201
*|10201,10202
0|10202,10203
<EOL>|10203,10204
25|10204,10206
.|10206,10207
Ipratropium|10208,10219
Bromide|10220,10227
Neb|10228,10231
1|10232,10233
NEB|10234,10237
IH|10238,10240
Q6H|10241,10244
:|10244,10245
PRN|10245,10248
dyspnea|10249,10256
,|10256,10257
wheezing|10258,10266
<EOL>|10267,10268
RX|10268,10270
*|10271,10272
ipratropium|10272,10283
bromide|10284,10291
0.2|10292,10295
mg|10296,10298
/|10298,10299
mL|10299,10301
(|10303,10304
0.02|10304,10308
%|10309,10310
)|10310,10311
1|10312,10313
neb|10314,10317
INH|10318,10321
Every|10322,10327
six|10328,10331
<EOL>|10332,10333
hours|10333,10338
Disp|10339,10343
#|10344,10345
*|10345,10346
30|10346,10348
Nebule|10349,10355
Refills|10356,10363
:|10363,10364
*|10364,10365
0|10365,10366
<EOL>|10366,10367
26|10367,10369
.|10369,10370
PredniSONE|10371,10381
10|10382,10384
mg|10385,10387
PO|10388,10390
ASDIR|10391,10396
<EOL>|10397,10398
50|10398,10400
mg|10401,10403
_|10404,10405
_|10405,10406
_|10406,10407
,|10407,10408
then|10409,10413
<EOL>|10414,10415
40|10415,10417
mg|10418,10420
_|10421,10422
_|10422,10423
_|10423,10424
,|10424,10425
then|10426,10430
<EOL>|10430,10431
30|10431,10433
mg|10434,10436
_|10437,10438
_|10438,10439
_|10439,10440
,|10440,10441
then|10442,10446
<EOL>|10446,10447
20|10447,10449
mg|10450,10452
_|10453,10454
_|10454,10455
_|10455,10456
,|10456,10457
then|10458,10462
<EOL>|10462,10463
10|10463,10465
mg|10466,10468
ongoing|10469,10476
<EOL>|10477,10478
Tapered|10478,10485
dose|10486,10490
-|10491,10492
DOWN|10493,10497
<EOL>|10498,10499
RX|10499,10501
*|10502,10503
prednisone|10503,10513
10|10514,10516
mg|10517,10519
1|10520,10521
to|10522,10524
5|10525,10526
tablet|10527,10533
(|10533,10534
s|10534,10535
)|10535,10536
by|10537,10539
mouth|10540,10545
As|10546,10548
directed|10549,10557
Disp|10558,10562
<EOL>|10563,10564
#|10564,10565
*|10565,10566
50|10566,10568
Tablet|10569,10575
Refills|10576,10583
:|10583,10584
*|10584,10585
0|10585,10586
<EOL>|10586,10587
<EOL>|10587,10588
<EOL>|10589,10590
Discharge|10590,10599
Disposition|10600,10611
:|10611,10612
<EOL>|10612,10613
Home|10613,10617
With|10618,10622
Service|10623,10630
<EOL>|10630,10631
<EOL>|10632,10633
Facility|10633,10641
:|10641,10642
<EOL>|10642,10643
_|10643,10644
_|10644,10645
_|10645,10646
<EOL>|10646,10647
<EOL>|10648,10649
Discharge|10649,10658
Diagnosis|10659,10668
:|10668,10669
<EOL>|10669,10670
Primary|10670,10677
diagnoses|10678,10687
:|10687,10688
<EOL>|10688,10689
Chronic|10689,10696
obstructive|10697,10708
pulmonary|10709,10718
disease|10719,10726
<EOL>|10726,10727
Atrial|10727,10733
fibrillation|10734,10746
with|10747,10751
rapid|10752,10757
ventricular|10758,10769
response|10770,10778
<EOL>|10778,10779
<EOL>|10779,10780
Secondary|10780,10789
diagnoses|10790,10799
:|10799,10800
<EOL>|10800,10801
Hypertension|10801,10813
<EOL>|10813,10814
Coronary|10814,10822
artery|10823,10829
disease|10830,10837
<EOL>|10837,10838
Peripheral|10838,10848
vascular|10849,10857
disease|10858,10865
<EOL>|10865,10866
<EOL>|10866,10867
<EOL>|10868,10869
Discharge|10869,10878
Condition|10879,10888
:|10888,10889
<EOL>|10889,10890
Mental|10890,10896
Status|10897,10903
:|10903,10904
Clear|10905,10910
and|10911,10914
coherent|10915,10923
.|10923,10924
<EOL>|10924,10925
Level|10925,10930
of|10931,10933
Consciousness|10934,10947
:|10947,10948
Alert|10949,10954
and|10955,10958
interactive|10959,10970
.|10970,10971
<EOL>|10971,10972
Activity|10972,10980
Status|10981,10987
:|10987,10988
Ambulatory|10989,10999
-|11000,11001
Independent|11002,11013
.|11013,11014
<EOL>|11014,11015
<EOL>|11015,11016
<EOL>|11017,11018
Discharge|11018,11027
Instructions|11028,11040
:|11040,11041
<EOL>|11041,11042
Dear|11042,11046
Ms.|11047,11050
_|11051,11052
_|11052,11053
_|11053,11054
,|11054,11055
<EOL>|11055,11056
<EOL>|11056,11057
You|11057,11060
were|11061,11065
hospitalized|11066,11078
at|11079,11081
_|11082,11083
_|11083,11084
_|11084,11085
<EOL>|11086,11087
because|11087,11094
you|11095,11098
were|11099,11103
having|11104,11110
difficulty|11111,11121
breathing|11122,11131
and|11132,11135
were|11136,11140
found|11141,11146
in|11147,11149
<EOL>|11150,11151
clinic|11151,11157
to|11158,11160
have|11161,11165
a|11166,11167
fast|11168,11172
heart|11173,11178
rate|11179,11183
.|11183,11184
Your|11185,11189
difficulty|11190,11200
breathing|11201,11210
was|11211,11214
<EOL>|11215,11216
due|11216,11219
to|11220,11222
your|11223,11227
COPD|11228,11232
flaring|11233,11240
.|11240,11241
Your|11242,11246
fast|11247,11251
heart|11252,11257
rate|11258,11262
was|11263,11266
due|11267,11270
to|11271,11273
your|11274,11278
<EOL>|11279,11280
atrial|11280,11286
fibrillation|11287,11299
,|11299,11300
which|11301,11306
is|11307,11309
an|11310,11312
irregular|11313,11322
heart|11323,11328
rate|11329,11333
that|11334,11338
can|11339,11342
<EOL>|11343,11344
sometimes|11344,11353
cause|11354,11359
the|11360,11363
heart|11364,11369
to|11370,11372
beat|11373,11377
very|11378,11382
quickly|11383,11390
.|11390,11391
Medications|11392,11403
that|11404,11408
<EOL>|11409,11410
you|11410,11413
were|11414,11418
taking|11419,11425
,|11425,11426
such|11427,11431
as|11432,11434
theophylline|11435,11447
,|11447,11448
were|11449,11453
likely|11454,11460
contributing|11461,11473
.|11473,11474
<EOL>|11475,11476
Your|11476,11480
heart|11481,11486
rate|11487,11491
was|11492,11495
lowered|11496,11503
using|11504,11509
the|11510,11513
same|11514,11518
medication|11519,11529
that|11530,11534
you|11535,11538
<EOL>|11539,11540
take|11540,11544
at|11545,11547
home|11548,11552
,|11552,11553
diltiazem|11554,11563
,|11563,11564
given|11565,11570
through|11571,11578
your|11579,11583
IV|11584,11586
.|11586,11587
<EOL>|11588,11589
<EOL>|11589,11590
Your|11590,11594
COPD|11595,11599
was|11600,11603
likely|11604,11610
worsened|11611,11619
because|11620,11627
of|11628,11630
a|11631,11632
cold|11633,11637
.|11637,11638
However|11639,11646
,|11646,11647
your|11648,11652
<EOL>|11653,11654
flare|11654,11659
was|11660,11663
very|11664,11668
serious|11669,11676
requiring|11677,11686
IV|11687,11689
steroids|11690,11698
and|11699,11702
many|11703,11707
inhaled|11708,11715
<EOL>|11716,11717
treatments|11717,11727
.|11727,11728
You|11729,11732
should|11733,11739
follow|11740,11746
up|11747,11749
with|11750,11754
the|11755,11758
lung|11759,11763
doctors|11764,11771
as|11772,11774
_|11775,11776
_|11776,11777
_|11777,11778
<EOL>|11779,11780
as|11780,11782
with|11783,11787
pulmonary|11788,11797
rehab|11798,11803
to|11804,11806
make|11807,11811
sure|11812,11816
your|11817,11821
lung|11822,11826
disease|11827,11834
is|11835,11837
being|11838,11843
<EOL>|11844,11845
treated|11845,11852
as|11853,11855
well|11856,11860
as|11861,11863
possible|11864,11872
to|11873,11875
prevent|11876,11883
you|11884,11887
from|11888,11892
coming|11893,11899
into|11900,11904
the|11905,11908
<EOL>|11909,11910
hospital|11910,11918
as|11919,11921
often|11922,11927
.|11927,11928
Please|11929,11935
call|11936,11940
_|11941,11942
_|11942,11943
_|11943,11944
to|11945,11947
schedule|11948,11956
an|11957,11959
<EOL>|11960,11961
appointment|11961,11972
with|11973,11977
them|11978,11982
.|11982,11983
<EOL>|11983,11984
<EOL>|11984,11985
It|11985,11987
was|11988,11991
a|11992,11993
pleasure|11994,12002
participating|12003,12016
in|12017,12019
your|12020,12024
care|12025,12029
.|12029,12030
We|12031,12033
wish|12034,12038
you|12039,12042
all|12043,12046
<EOL>|12047,12048
the|12048,12051
best|12052,12056
in|12057,12059
the|12060,12063
future|12064,12070
.|12070,12071
<EOL>|12071,12072
<EOL>|12072,12073
Sincerely|12073,12082
,|12082,12083
<EOL>|12083,12084
<EOL>|12084,12085
Your|12085,12089
_|12090,12091
_|12091,12092
_|12092,12093
team|12094,12098
<EOL>|12098,12099
<EOL>|12100,12101
Followup|12101,12109
Instructions|12110,12122
:|12122,12123
<EOL>|12123,12124
_|12124,12125
_|12125,12126
_|12126,12127
<EOL>|12127,12128

