 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|168,177|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|168,177|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|168,177|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Antibiotic|SIMPLE_SEGMENT|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|SIMPLE_SEGMENT|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|SIMPLE_SEGMENT|180,189|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Event|Event|SIMPLE_SEGMENT|180,189|false|false|false|||meropenem
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|210,225|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|216,225|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|216,225|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|216,225|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Functional Concept|SIMPLE_SEGMENT|227,231|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|227,235|false|false|false|C0524471|Left hip region structure|left hip
Finding|Sign or Symptom|SIMPLE_SEGMENT|227,240|false|false|false|C2141922|Pain of left hip joint|left hip pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|232,235|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|232,235|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|232,235|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|232,235|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|232,240|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|232,240|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|236,240|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|236,240|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|236,240|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|236,240|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|243,248|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|249,257|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|249,257|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|261,279|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|270,279|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|270,279|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|270,279|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|270,279|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|270,279|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|288,297|false|false|false|||reduction
Finding|Finding|SIMPLE_SEGMENT|288,297|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|288,297|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|288,297|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Finding|Functional Concept|SIMPLE_SEGMENT|302,314|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|SIMPLE_SEGMENT|315,322|false|false|false|||pinning
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|315,322|false|false|false|C0021885|Intramedullary Nailing|pinning
Event|Event|SIMPLE_SEGMENT|324,328|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|324,328|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|329,336|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|329,341|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|329,350|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|SIMPLE_SEGMENT|337,341|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|337,341|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|337,341|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|337,350|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|342,350|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|342,350|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|354,361|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|354,361|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,364|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|354,380|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|354,380|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|365,372|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|365,372|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|365,380|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|373,380|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|427,430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|427,430|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|434,446|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|434,446|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|457,466|false|false|false|||sustained
Event|Event|SIMPLE_SEGMENT|469,479|false|false|false|||mechanical
Finding|Functional Concept|SIMPLE_SEGMENT|469,479|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|469,479|false|false|false|C0699886|Mechanical Treatments|mechanical
Event|Event|SIMPLE_SEGMENT|480,484|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|480,484|false|false|false|C0085639|Falls|fall
Finding|Functional Concept|SIMPLE_SEGMENT|494,498|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|499,504|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|499,504|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|506,515|false|false|false|C0015385|Limb structure|extremity
Finding|Idea or Concept|SIMPLE_SEGMENT|521,530|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|521,530|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|immediate
Attribute|Clinical Attribute|SIMPLE_SEGMENT|531,535|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|531,535|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|531,535|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|531,535|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|537,546|false|false|false|||inability
Finding|Finding|SIMPLE_SEGMENT|537,558|false|false|false|C5436357|Inability to ambulate|inability to ambulate
Event|Event|SIMPLE_SEGMENT|550,558|false|false|false|||ambulate
Finding|Finding|SIMPLE_SEGMENT|550,558|false|false|false|C4036205|Ambulate|ambulate
Finding|Body Substance|SIMPLE_SEGMENT|566,573|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|566,573|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|566,573|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|574,580|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|581,584|true|false|false|||LOC
Event|Event|SIMPLE_SEGMENT|598,606|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|598,606|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|598,606|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|611,614|true|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|611,614|true|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|611,614|true|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|SIMPLE_SEGMENT|611,614|true|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|611,614|true|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|SIMPLE_SEGMENT|611,614|true|false|false|||ROS
Finding|Gene or Genome|SIMPLE_SEGMENT|611,614|true|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|SIMPLE_SEGMENT|611,614|true|false|false|C0489633|Review of systems (procedure)|ROS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|632,640|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|632,640|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|632,640|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|SIMPLE_SEGMENT|646,666|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|651,658|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|651,658|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|651,658|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|651,658|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|651,658|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|651,666|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|659,666|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|659,666|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|659,666|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|668,674|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|668,674|false|false|false|||Anemia
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|677,699|false|false|false|C0694540|borderline cholesterol|Borderline cholesterol
Drug|Biologically Active Substance|SIMPLE_SEGMENT|688,699|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|SIMPLE_SEGMENT|688,699|false|false|false|C0008377|cholesterol|cholesterol
Event|Event|SIMPLE_SEGMENT|688,699|false|false|false|||cholesterol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|688,699|false|false|false|C0201950|Cholesterol measurement|cholesterol
Finding|Sign or Symptom|SIMPLE_SEGMENT|722,732|false|false|false|C0016204|Flatulence|Flatulence
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|735,740|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|735,740|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|735,740|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|735,747|false|false|false|C0018808|Heart murmur|Heart Murmur
Event|Event|SIMPLE_SEGMENT|741,747|false|false|false|||Murmur
Finding|Finding|SIMPLE_SEGMENT|741,747|false|false|false|C0018808|Heart murmur|Murmur
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|750,762|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|750,762|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|765,779|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|765,779|false|false|false|||Hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|782,802|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral Regurgitation
Event|Event|SIMPLE_SEGMENT|789,802|false|false|false|||Regurgitation
Finding|Finding|SIMPLE_SEGMENT|789,802|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|789,802|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|789,802|false|false|false|C0460152|Regurgitation - mechanism|Regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|805,817|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|805,817|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|805,817|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|820,829|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|SIMPLE_SEGMENT|820,829|false|false|false|||Pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|832,841|false|false|false|C0037199|Sinusitis|Sinusitis
Event|Event|SIMPLE_SEGMENT|832,841|false|false|false|||Sinusitis
Finding|Functional Concept|SIMPLE_SEGMENT|855,861|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|855,869|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|862,869|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|862,869|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|862,869|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|862,869|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|875,881|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|875,881|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|875,881|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|875,881|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|875,889|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|882,889|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|882,889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|882,889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|882,889|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|896,903|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|896,903|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|896,906|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|896,919|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|907,919|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|907,919|false|false|false|||hypertension
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|923,933|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|923,933|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|923,933|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|927,933|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|927,933|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|936,942|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|936,942|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Classification|SIMPLE_SEGMENT|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|945,951|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|959,966|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|959,966|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|959,969|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|979,986|false|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|979,986|false|false|false|||cancers
Event|Event|SIMPLE_SEGMENT|999,1010|false|false|false|||grandfather
Event|Event|SIMPLE_SEGMENT|1019,1026|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1019,1026|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1019,1029|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1030,1037|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1030,1037|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1030,1037|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|1030,1037|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|1030,1037|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1030,1037|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1030,1044|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1038,1044|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1038,1044|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1065,1072|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1065,1072|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1065,1075|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1076,1082|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1076,1082|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1076,1082|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|SIMPLE_SEGMENT|1076,1082|false|false|false|||throat
Finding|Body Substance|SIMPLE_SEGMENT|1076,1082|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|1076,1082|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1084,1090|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1084,1090|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1096,1103|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1096,1103|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1096,1106|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1107,1112|true|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1107,1112|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1107,1112|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|1107,1112|true|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1107,1120|true|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1113,1120|true|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|1113,1120|true|false|false|||cancers
Finding|Conceptual Entity|SIMPLE_SEGMENT|1122,1128|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1122,1128|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1133,1139|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1133,1139|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1133,1139|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|SIMPLE_SEGMENT|1145,1151|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1145,1151|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1145,1151|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1145,1151|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1160,1166|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1173,1178|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1173,1178|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1173,1178|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1173,1184|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1179,1184|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|1185,1193|false|false|false|||replaced
Event|Event|SIMPLE_SEGMENT|1198,1206|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1198,1206|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1198,1206|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1198,1206|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1198,1211|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1198,1211|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1207,1211|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1207,1211|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1207,1211|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1216,1225|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1216,1225|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1228,1234|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1228,1234|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1228,1234|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|SIMPLE_SEGMENT|1228,1234|false|false|false|C0812455|Pelvis problem|Pelvis
Event|Event|SIMPLE_SEGMENT|1235,1241|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1235,1241|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|1260,1271|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|1260,1271|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1260,1271|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|1260,1271|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1260,1271|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Anatomy|Body System|SIMPLE_SEGMENT|1279,1283|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1279,1283|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1279,1283|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|1279,1283|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|1279,1283|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|SIMPLE_SEGMENT|1279,1289|false|false|false|C0574729|Skin clean|skin clean
Event|Activity|SIMPLE_SEGMENT|1284,1289|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|SIMPLE_SEGMENT|1294,1300|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|1294,1300|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|1302,1305|false|false|false|||LLE
Event|Event|SIMPLE_SEGMENT|1306,1315|false|false|false|||Shortened
Event|Event|SIMPLE_SEGMENT|1331,1338|false|false|false|||rotated
Event|Event|SIMPLE_SEGMENT|1340,1347|false|false|false|||painful
Finding|Sign or Symptom|SIMPLE_SEGMENT|1340,1347|false|false|false|C0030193|Pain|painful
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1366,1374|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|SIMPLE_SEGMENT|1366,1374|false|false|false|C0521134|External route|external
Finding|Functional Concept|SIMPLE_SEGMENT|1366,1383|false|false|false|C0231462|External rotation|external rotation
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1375,1383|false|false|false|C3669037|Rotation (malposition) (morphologic abnormality)|rotation
Event|Event|SIMPLE_SEGMENT|1375,1383|false|false|false|||rotation
Finding|Finding|SIMPLE_SEGMENT|1375,1383|false|false|false|C0035868;C0677597;C2117331|Musculoskeletal rotation;Rotation|rotation
Finding|Functional Concept|SIMPLE_SEGMENT|1375,1383|false|false|false|C0035868;C0677597;C2117331|Musculoskeletal rotation;Rotation|rotation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1391,1394|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1391,1394|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|1391,1394|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1391,1394|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1398,1404|false|false|false|C0039866|Thigh structure|Thighs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1409,1412|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|1413,1425|false|false|false|||compartments
Finding|Intellectual Product|SIMPLE_SEGMENT|1413,1425|false|false|false|C1185625|Anatomical compartments|compartments
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1413,1425|false|false|false|C1382196|Compartments [PK]|compartments
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1426,1430|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|1426,1430|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|1432,1441|false|false|false|||Saphenous
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1443,1448|false|false|false|C0626053|sural|Sural
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1450,1454|false|false|false|C4318566|Deep Resection Margin|Deep
Event|Event|SIMPLE_SEGMENT|1486,1490|false|false|false|||SILT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1496,1499|false|false|false|C0265372;C3665330|Feline hyperesthesia syndrome;Fetal hydantoin syndrome|FHS
Event|Event|SIMPLE_SEGMENT|1496,1499|false|false|false|||FHS
Finding|Finding|SIMPLE_SEGMENT|1496,1499|false|false|false|C0241889|Family Medical History|FHS
Event|Event|SIMPLE_SEGMENT|1517,1521|false|false|false|C0016141|fire disaster|Fire
Finding|Gene or Genome|SIMPLE_SEGMENT|1517,1521|false|false|false|C1426107|ADGRE4P gene|Fire
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1517,1521|false|false|false|C0000912;C0700614;C0702194|Accident caused by unspecified fire;Fire (physical force);Fire as a heat source|Fire
Drug|Food|SIMPLE_SEGMENT|1537,1543|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|1537,1543|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|1537,1543|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|1537,1543|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1545,1549|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1545,1549|false|false|false|C0562271|Examination of knee joint|Knee
Event|Event|SIMPLE_SEGMENT|1550,1556|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1550,1556|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1570,1576|false|false|false|C0042282|Valgus deformity|valgus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1577,1583|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|1577,1583|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1577,1583|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|1577,1583|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|1577,1583|false|false|false|C0038435|Stress|stress
Finding|Classification|SIMPLE_SEGMENT|1588,1596|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|1588,1596|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1588,1596|false|false|false|C5237010|Expression Negative|Negative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1597,1605|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|1597,1605|false|false|false|||anterior
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1607,1616|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|SIMPLE_SEGMENT|1624,1629|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|1624,1629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1624,1629|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|1637,1646|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1637,1646|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1637,1646|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1649,1652|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1649,1652|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1649,1652|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1649,1652|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1649,1652|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1660,1668|false|false|false|C2338258|Cranial incision point|INcision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1660,1668|false|false|false|C0332803|Surgical wound|INcision
Event|Event|SIMPLE_SEGMENT|1660,1668|false|false|false|||INcision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1660,1668|false|false|false|C0184898|Surgical incisions|INcision
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1670,1678|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|SIMPLE_SEGMENT|1670,1678|false|false|false|||dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1670,1678|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|1670,1678|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|1670,1678|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1670,1678|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|SIMPLE_SEGMENT|1679,1686|false|false|false|||changed
Event|Event|SIMPLE_SEGMENT|1715,1721|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|1715,1721|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|1732,1738|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|1732,1738|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|1740,1744|false|false|false|||SILT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1783,1788|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|1783,1788|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|1783,1788|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1783,1788|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|1783,1788|false|false|false|C0034107|Pulse taking|pulse
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1811,1814|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|Hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1811,1814|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Event|Event|SIMPLE_SEGMENT|1811,1814|false|false|false|||Hip
Finding|Gene or Genome|SIMPLE_SEGMENT|1811,1814|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|Hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1811,1814|false|false|false|C1292890|Procedure on hip|Hip
Event|Event|SIMPLE_SEGMENT|1823,1833|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|1823,1833|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|1823,1833|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1836,1844|false|false|false|C0040456|Impacted tooth|Impacted
Event|Event|SIMPLE_SEGMENT|1836,1844|false|false|false|||Impacted
Finding|Functional Concept|SIMPLE_SEGMENT|1836,1844|false|false|false|C0333125|Impacted|Impacted
Finding|Functional Concept|SIMPLE_SEGMENT|1845,1849|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1861,1868|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1861,1873|false|false|false|C0015815|Structure of neck of femur|femoral neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1869,1873|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|1869,1873|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|1869,1873|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1875,1883|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|1875,1883|false|false|false|||fracture
Finding|Intellectual Product|SIMPLE_SEGMENT|1887,1892|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|1893,1901|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1893,1908|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|1893,1908|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|1928,1936|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|1944,1949|false|false|false|C0812371|Ortho-|ortho
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1950,1956|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|1950,1956|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|1950,1956|false|false|false|C0548346|Trauma assessment and care|trauma
Event|Occupational Activity|SIMPLE_SEGMENT|1957,1964|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|1957,1964|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|SIMPLE_SEGMENT|1970,1975|false|false|false|||found
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1986,1992|false|false|false|C0042282|Valgus deformity|valgus
Event|Event|SIMPLE_SEGMENT|1993,2001|false|false|false|||impacted
Finding|Functional Concept|SIMPLE_SEGMENT|2002,2006|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2002,2019|false|false|false|C0833290|Neck of left femur|left femoral neck
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2007,2014|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2007,2019|false|false|false|C0015815|Structure of neck of femur|femoral neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2015,2019|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2015,2019|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|2015,2019|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2020,2023|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2020,2023|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|2020,2023|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2020,2023|false|false|false|C1292890|Procedure on hip|hip
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2020,2032|false|false|false|C0019557;C0149531|Fracture of pelvis;Hip Fractures|hip fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2024,2032|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|2024,2032|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|2066,2075|false|false|false|||reduction
Finding|Finding|SIMPLE_SEGMENT|2066,2075|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2066,2075|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2066,2075|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Event|Event|SIMPLE_SEGMENT|2080,2092|false|false|false|||percutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|2080,2092|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|SIMPLE_SEGMENT|2094,2101|false|false|false|||pinning
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2094,2101|false|false|false|C0021885|Intramedullary Nailing|pinning
Event|Event|SIMPLE_SEGMENT|2103,2107|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|2103,2107|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2108,2115|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2108,2120|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2108,2129|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2116,2120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2116,2120|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|2116,2120|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2116,2129|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2121,2129|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|2121,2129|false|false|false|||fracture
Finding|Body Substance|SIMPLE_SEGMENT|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2153,2160|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2165,2170|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|2177,2187|false|false|false|||recovering
Finding|Finding|SIMPLE_SEGMENT|2188,2192|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2199,2206|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2199,2206|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2199,2206|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|2212,2218|false|false|false|||became
Event|Event|SIMPLE_SEGMENT|2219,2230|false|false|false|||hypotensive
Finding|Pathologic Function|SIMPLE_SEGMENT|2219,2230|false|false|false|C0857353|Hypotensive|hypotensive
Finding|Finding|SIMPLE_SEGMENT|2236,2244|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|2236,2244|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2236,2244|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|2236,2252|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2236,2252|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|2245,2252|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|2245,2252|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|2245,2252|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2245,2252|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|2261,2271|false|false|false|||normalized
Event|Event|SIMPLE_SEGMENT|2287,2295|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|2287,2295|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2287,2295|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Body Substance|SIMPLE_SEGMENT|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2310,2317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2318,2327|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|2334,2338|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|2334,2338|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2348,2352|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|2357,2365|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|2357,2365|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2357,2365|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|2357,2373|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2357,2373|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|2366,2373|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|2366,2373|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|2366,2373|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2366,2373|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|2378,2385|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|2390,2399|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2390,2399|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2390,2399|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2405,2410|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|2411,2419|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|2411,2419|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Functional Concept|SIMPLE_SEGMENT|2422,2428|false|false|false|C0728831|Social|SOcial
Event|Event|SIMPLE_SEGMENT|2429,2433|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|2429,2433|false|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|2434,2437|false|false|false|||saw
Finding|Finding|SIMPLE_SEGMENT|2449,2459|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|SIMPLE_SEGMENT|2449,2466|false|false|false|C0582154|Difficulty coping|difficulty coping
Event|Event|SIMPLE_SEGMENT|2460,2466|false|false|false|||coping
Finding|Finding|SIMPLE_SEGMENT|2460,2466|false|true|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Finding|Individual Behavior|SIMPLE_SEGMENT|2460,2466|false|true|false|C0009967;C0517270|Child coping with hospitalization;Coping Behavior|coping
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2460,2466|false|true|false|C2700390;C3502819|COPING - Dental Restorative Procedure;COPING - Fixed Prosthodontics|coping
Event|Event|SIMPLE_SEGMENT|2472,2481|false|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|2472,2481|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2483,2491|false|false|false|C0080078|Range of Motion, Articular|mobility
Event|Event|SIMPLE_SEGMENT|2483,2491|false|false|false|||mobility
Finding|Finding|SIMPLE_SEGMENT|2483,2491|false|false|false|C0425245|Mobility finding|mobility
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2497,2501|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|2502,2508|false|false|false|||showed
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2509,2515|false|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|2509,2515|false|true|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2509,2515|false|true|false|C0337443|Sodium measurement|sodium
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2509,2521|false|false|false|C0428291|Finding of sodium level|sodium level
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2509,2521|false|false|false|C0337443|Sodium measurement|sodium level
Event|Event|SIMPLE_SEGMENT|2516,2521|false|false|false|||level
Event|Event|SIMPLE_SEGMENT|2530,2539|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|2530,2539|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|2554,2561|false|false|false|||similar
Event|Event|SIMPLE_SEGMENT|2572,2581|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2572,2581|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2597,2609|false|false|false|C3263700||instructions
Event|Event|SIMPLE_SEGMENT|2597,2609|false|false|false|||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|2597,2609|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Drug|Organic Chemical|SIMPLE_SEGMENT|2669,2676|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2669,2676|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|2669,2676|false|false|false|||lovenox
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2714,2725|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2714,2725|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|2714,2725|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2714,2725|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|2714,2738|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|2729,2738|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2729,2738|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2757,2767|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|2757,2767|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|2757,2772|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|2768,2772|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|2768,2772|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|2776,2784|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|2789,2797|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|2789,2797|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|2789,2797|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|2789,2797|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2802,2815|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|SIMPLE_SEGMENT|2802,2815|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2802,2822|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2816,2822|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|2816,2822|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|2816,2822|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2816,2822|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2843,2853|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2843,2853|false|false|false|C0065374|lisinopril|Lisinopril
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2872,2887|false|false|false|C2878629|Poisoning by, adverse effect of and underdosing of methylphenidate|MethylPHENIDATE
Drug|Organic Chemical|SIMPLE_SEGMENT|2872,2887|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2872,2887|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Event|Event|SIMPLE_SEGMENT|2872,2887|false|false|false|||MethylPHENIDATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2872,2887|false|false|false|C0524188|Methylphenidate measurement|MethylPHENIDATE
Drug|Organic Chemical|SIMPLE_SEGMENT|2889,2896|false|false|false|C0728759|Ritalin|Ritalin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2889,2896|false|false|false|C0728759|Ritalin|Ritalin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2908,2911|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2908,2911|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2908,2911|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|2908,2911|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|2908,2911|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|2916,2927|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2916,2927|false|false|false|C0049506|mirtazapine|mirtazapine
Event|Event|SIMPLE_SEGMENT|2916,2927|false|false|false|||mirtazapine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2934,2938|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2934,2938|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|2934,2938|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|2934,2938|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Event|Event|SIMPLE_SEGMENT|2939,2942|false|false|false|||QHS
Event|Event|SIMPLE_SEGMENT|2947,2956|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2947,2956|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2947,2956|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|2947,2968|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2957,2968|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2957,2968|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|2957,2968|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2957,2968|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2973,2986|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|SIMPLE_SEGMENT|2973,2986|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2973,2993|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2987,2993|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|2987,2993|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|2987,2993|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2987,2993|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3014,3024|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3014,3024|false|false|false|C0065374|lisinopril|Lisinopril
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3043,3058|false|false|false|C2878629|Poisoning by, adverse effect of and underdosing of methylphenidate|MethylPHENIDATE
Drug|Organic Chemical|SIMPLE_SEGMENT|3043,3058|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3043,3058|false|false|false|C0025810|methylphenidate|MethylPHENIDATE
Event|Event|SIMPLE_SEGMENT|3043,3058|false|false|false|||MethylPHENIDATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3043,3058|false|false|false|C0524188|Methylphenidate measurement|MethylPHENIDATE
Drug|Organic Chemical|SIMPLE_SEGMENT|3060,3067|false|false|false|C0728759|Ritalin|Ritalin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3060,3067|false|false|false|C0728759|Ritalin|Ritalin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3079,3082|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3079,3082|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3079,3082|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|3079,3082|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|3079,3082|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|3087,3098|false|false|false|C0049506|mirtazapine|mirtazapine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3087,3098|false|false|false|C0049506|mirtazapine|mirtazapine
Event|Event|SIMPLE_SEGMENT|3087,3098|false|false|false|||mirtazapine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3105,3109|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3105,3109|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|3105,3109|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|3105,3109|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Event|Event|SIMPLE_SEGMENT|3110,3113|false|false|false|||QHS
Drug|Organic Chemical|SIMPLE_SEGMENT|3118,3131|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3118,3131|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|3118,3131|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3118,3131|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Event|Event|SIMPLE_SEGMENT|3143,3146|false|false|false|||TID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3151,3159|false|false|false|C0002367|aluminum|Aluminum
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3151,3159|false|false|false|C0002367|aluminum|Aluminum
Event|Event|SIMPLE_SEGMENT|3151,3159|false|false|false|||Aluminum
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3151,3159|false|false|false|C0202311|Aluminum measurement|Aluminum
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3160,3169|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|Magnesium
Event|Event|SIMPLE_SEGMENT|3160,3169|false|false|false|||Magnesium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3160,3169|false|false|false|C0373675|Magnesium measurement|Magnesium
Drug|Organic Chemical|SIMPLE_SEGMENT|3178,3189|false|false|false|C0037138|simethicone|Simethicone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3178,3189|false|false|false|C0037138|simethicone|Simethicone
Event|Event|SIMPLE_SEGMENT|3200,3203|false|false|false|||QID
Finding|Gene or Genome|SIMPLE_SEGMENT|3204,3207|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|3209,3218|false|false|false|||Dyspepsia
Finding|Sign or Symptom|SIMPLE_SEGMENT|3209,3218|false|false|false|C0013395|Dyspepsia|Dyspepsia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3223,3239|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Event|Event|SIMPLE_SEGMENT|3234,3239|false|false|false|||Tears
Finding|Body Substance|SIMPLE_SEGMENT|3234,3239|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|SIMPLE_SEGMENT|3234,3239|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3244,3248|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|3244,3248|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|3244,3248|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3249,3258|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3254,3258|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3254,3258|false|false|false|C5848506||EYES
Event|Event|SIMPLE_SEGMENT|3259,3262|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|3259,3262|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3263,3271|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3263,3271|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3263,3271|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3267,3271|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3267,3271|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|3267,3271|false|false|false|||eyes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Enzyme|SIMPLE_SEGMENT|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3276,3283|false|false|false|C0673636|Biotene|Biotene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3276,3293|true|false|false|C5762022|Biotene Dry Mouth|Biotene Dry Mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3284,3293|true|false|false|C0043352|Xerostomia|Dry Mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3288,3293|true|false|false|C0226896;C0230028|Oral cavity;Oral region|Mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3288,3293|true|false|false|C0226896;C0230028|Oral cavity;Oral region|Mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3288,3299|true|false|false|C0026647|Mouthwash|Mouth Rinse
Finding|Body Substance|SIMPLE_SEGMENT|3288,3299|true|false|false|C5849077|Mouth Rinse Specimen|Mouth Rinse
Event|Activity|SIMPLE_SEGMENT|3294,3299|true|false|false|C1882955|Rinsing|Rinse
Event|Event|SIMPLE_SEGMENT|3294,3299|true|false|false|||Rinse
Finding|Functional Concept|SIMPLE_SEGMENT|3294,3299|true|false|false|C1701810|Rinse Dosage Form|Rinse
Finding|Body Substance|SIMPLE_SEGMENT|3301,3307|true|false|false|C0036087;C0438730;C1546769|Saliva specimen;saliva|saliva
Finding|Intellectual Product|SIMPLE_SEGMENT|3301,3307|true|false|false|C0036087;C0438730;C1546769|Saliva specimen;saliva|saliva
Event|Activity|SIMPLE_SEGMENT|3308,3320|true|false|false|C1706204|Substitution - change|substitution
Event|Event|SIMPLE_SEGMENT|3308,3320|true|false|false|||substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|3308,3320|true|false|false|C1555721|Substitution - ActClass|substitution
Event|Event|SIMPLE_SEGMENT|3321,3326|true|false|false|||combo
Event|Event|SIMPLE_SEGMENT|3336,3347|false|false|false|||application
Finding|Functional Concept|SIMPLE_SEGMENT|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|SIMPLE_SEGMENT|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|SIMPLE_SEGMENT|3336,3347|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3336,3347|false|false|false|C0185125|Application procedure|application
Finding|Body Substance|SIMPLE_SEGMENT|3348,3354|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|Mucous
Anatomy|Tissue|SIMPLE_SEGMENT|3348,3363|false|false|false|C0026724|Mucous Membrane|Mucous Membrane
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3348,3363|false|false|false|C0151785|Disease of mucous membrane|Mucous Membrane
Finding|Functional Concept|SIMPLE_SEGMENT|3348,3363|false|false|false|C1549524|Route of Administration - Mucous Membrane|Mucous Membrane
Anatomy|Cell Component|SIMPLE_SEGMENT|3355,3363|false|false|false|C0025255;C0596901|Membrane;Membrane Tissue|Membrane
Anatomy|Tissue|SIMPLE_SEGMENT|3355,3363|false|false|false|C0025255;C0596901|Membrane;Membrane Tissue|Membrane
Event|Event|SIMPLE_SEGMENT|3364,3368|false|false|false|||q2hr
Drug|Organic Chemical|SIMPLE_SEGMENT|3373,3382|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3373,3382|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|SIMPLE_SEGMENT|3401,3404|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|3405,3417|false|false|false|||Constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3405,3417|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3423,3430|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3423,3430|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3423,3430|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3423,3430|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3423,3440|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3423,3440|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3431,3440|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Event|Event|SIMPLE_SEGMENT|3452,3455|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|3461,3469|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3461,3469|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|3461,3469|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|3461,3476|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3461,3476|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3470,3476|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|3470,3476|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|3470,3476|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3470,3476|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3487,3490|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3487,3490|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3487,3490|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|3487,3490|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|3487,3490|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|3496,3506|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3496,3506|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|3496,3506|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|3496,3513|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3496,3513|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3507,3513|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|3507,3513|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|3507,3513|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3507,3513|false|false|false|C0337443|Sodium measurement|Sodium
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3529,3532|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3529,3532|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3529,3532|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3529,3544|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3533,3544|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3545,3553|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|3545,3553|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|3564,3569|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|3588,3592|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|SIMPLE_SEGMENT|3593,3600|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|3593,3600|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3593,3600|false|false|false|C1979801|Routine coag|Routine
Event|Event|SIMPLE_SEGMENT|3601,3615|false|false|false|||Administration
Event|Occupational Activity|SIMPLE_SEGMENT|3601,3615|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3601,3615|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|3617,3621|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|SIMPLE_SEGMENT|3627,3637|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3627,3637|false|false|false|C0206460|enoxaparin|enoxaparin
Event|Event|SIMPLE_SEGMENT|3627,3637|false|false|false|||enoxaparin
Event|Event|SIMPLE_SEGMENT|3687,3694|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|3687,3694|false|false|false|C0807726|refill|Refills
Drug|Food|SIMPLE_SEGMENT|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Immunologic Factor|SIMPLE_SEGMENT|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Substance|SIMPLE_SEGMENT|3702,3706|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Event|Event|SIMPLE_SEGMENT|3702,3706|false|false|false|||Milk
Finding|Body Substance|SIMPLE_SEGMENT|3702,3706|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Finding|Intellectual Product|SIMPLE_SEGMENT|3702,3706|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Drug|Clinical Drug|SIMPLE_SEGMENT|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3702,3718|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3710,3718|false|false|false|C0024477|magnesium oxide|Magnesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3710,3718|false|false|false|C0024477|magnesium oxide|Magnesia
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3728,3731|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3728,3731|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3728,3731|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|3728,3731|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|3728,3731|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|3732,3735|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|3736,3745|false|false|false|||Dyspepsia
Finding|Sign or Symptom|SIMPLE_SEGMENT|3736,3745|false|false|false|C0013395|Dyspepsia|Dyspepsia
Drug|Organic Chemical|SIMPLE_SEGMENT|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|3751,3764|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|3751,3764|false|false|false|||Multivitamins
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3767,3770|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3767,3770|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|3767,3770|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|3767,3770|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3767,3770|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|SIMPLE_SEGMENT|3771,3773|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|3785,3794|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3785,3794|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|SIMPLE_SEGMENT|3785,3794|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3785,3794|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|SIMPLE_SEGMENT|3796,3805|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|3796,3805|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3796,3813|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|SIMPLE_SEGMENT|3806,3813|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|3806,3813|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|3806,3813|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3806,3813|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|3830,3833|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3834,3838|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3834,3838|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3834,3838|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3834,3838|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3840,3842|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|3844,3853|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3844,3853|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|3844,3853|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3844,3853|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3863,3869|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|SIMPLE_SEGMENT|3863,3869|false|false|false|||tablet
Finding|Functional Concept|SIMPLE_SEGMENT|3873,3881|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3876,3881|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3876,3881|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|3899,3903|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|3899,3903|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3910,3916|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|3917,3924|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|3917,3924|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|3932,3944|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3932,3944|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|3964,3969|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3964,3969|false|false|false|C3489575|sennosides, USP|Senna
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3972,3975|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|3972,3975|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|3987,3994|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|3987,3996|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3987,3996|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|3995,3996|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|4001,4005|false|false|false|||UNIT
Event|Event|SIMPLE_SEGMENT|4019,4028|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4019,4028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4019,4028|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4019,4040|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|4019,4040|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4029,4040|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|4029,4040|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|4029,4040|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|4042,4050|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|4042,4050|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|4042,4055|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|4051,4055|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|4051,4055|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|4051,4055|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|4051,4055|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|4058,4066|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|4058,4066|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|4074,4083|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4074,4083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4074,4083|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|4074,4093|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4084,4093|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|4084,4093|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|4084,4093|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4084,4093|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4084,4093|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4095,4099|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4095,4112|false|false|false|C0833290|Neck of left femur|left femoral neck
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4100,4107|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4100,4112|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4100,4121|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4108,4112|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4108,4112|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|4108,4112|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4108,4121|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4113,4121|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|4113,4121|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|4125,4134|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4125,4134|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4125,4134|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4125,4134|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4125,4134|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4135,4144|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4135,4144|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|4135,4144|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|4135,4144|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|4146,4152|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4146,4159|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|4146,4159|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4153,4159|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4153,4159|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|4161,4166|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4161,4166|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|4171,4179|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|4171,4179|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|4181,4186|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4181,4203|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|4181,4203|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|4190,4203|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|4190,4203|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|4190,4203|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4205,4210|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|4205,4210|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4205,4210|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|4205,4210|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|4205,4210|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|4215,4226|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|4215,4226|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|4228,4236|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4228,4236|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|4228,4236|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4237,4243|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|4237,4243|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4237,4243|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4252,4255|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|4252,4255|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|4252,4255|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|4261,4271|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|4261,4271|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|4285,4295|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|4285,4295|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|4300,4309|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4300,4309|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4300,4309|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4300,4309|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4300,4309|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4300,4322|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4300,4322|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|4300,4322|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4310,4322|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|4310,4322|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4310,4322|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4324,4335|false|false|false|C0802604;C2598133||MEDICATIONS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4324,4335|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATIONS
Event|Event|SIMPLE_SEGMENT|4324,4335|false|false|false|||MEDICATIONS
Finding|Intellectual Product|SIMPLE_SEGMENT|4324,4335|false|false|false|C4284232|Medications|MEDICATIONS
Event|Event|SIMPLE_SEGMENT|4347,4351|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4356,4367|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4356,4367|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|4356,4367|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4356,4367|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|4371,4381|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|4405,4414|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4405,4414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4405,4414|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|4419,4427|false|false|false|||Continue
Finding|Idea or Concept|SIMPLE_SEGMENT|4432,4436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4432,4436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4432,4436|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4437,4448|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4437,4448|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|4437,4448|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4437,4448|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|4469,4479|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|4484,4488|false|false|false|||stop
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4497,4504|false|false|false|C5444295||surgeon
Event|Event|SIMPLE_SEGMENT|4516,4521|true|false|false|||drink
Drug|Organic Chemical|SIMPLE_SEGMENT|4522,4529|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4522,4529|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|4522,4529|true|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|4522,4529|true|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|SIMPLE_SEGMENT|4531,4536|true|false|false|||drive
Finding|Functional Concept|SIMPLE_SEGMENT|4539,4544|true|false|false|C1513492|motor movement|motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4545,4552|true|false|false|C0042444|Drug vehicle|vehicle
Event|Event|SIMPLE_SEGMENT|4545,4552|true|false|false|||vehicle
Event|Event|SIMPLE_SEGMENT|4557,4564|false|false|false|||operate
Finding|Functional Concept|SIMPLE_SEGMENT|4557,4564|false|false|false|C3242339|operate|operate
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4566,4575|false|false|false|C0337246|Contact with machinery|machinery
Event|Event|SIMPLE_SEGMENT|4566,4575|false|false|false|||machinery
Event|Event|SIMPLE_SEGMENT|4582,4588|false|false|false|||taking
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4589,4597|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4589,4597|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4598,4602|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4598,4602|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4598,4602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4598,4602|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|SIMPLE_SEGMENT|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4598,4612|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|SIMPLE_SEGMENT|4603,4612|false|false|false|||relievers
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4617,4625|false|false|false|C0027415|Narcotics|Narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4617,4625|false|false|false|C0027415|Narcotics|Narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4626,4630|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|4626,4630|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4626,4630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4626,4630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|SIMPLE_SEGMENT|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4626,4640|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|SIMPLE_SEGMENT|4631,4640|false|false|false|||relievers
Event|Event|SIMPLE_SEGMENT|4651,4663|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|4651,4663|false|false|false|C0009806|Constipation|constipation
Drug|Food|SIMPLE_SEGMENT|4680,4685|false|false|false|C0452428|Drink (dietary substance)|drink
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4707,4712|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4707,4712|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|SIMPLE_SEGMENT|4707,4712|false|false|false|||water
Finding|Intellectual Product|SIMPLE_SEGMENT|4707,4712|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4707,4712|false|false|false|C0020311|Hydrotherapy|water
Event|Event|SIMPLE_SEGMENT|4723,4727|false|false|false|||take
Finding|Body Substance|SIMPLE_SEGMENT|4730,4735|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|4730,4744|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4730,4744|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|SIMPLE_SEGMENT|4736,4744|false|false|false|||softener
Drug|Organic Chemical|SIMPLE_SEGMENT|4747,4753|false|false|false|C0282139|Colace|colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4747,4753|false|false|false|C0282139|Colace|colace
Event|Event|SIMPLE_SEGMENT|4758,4765|false|false|false|||prevent
Finding|Pathologic Function|SIMPLE_SEGMENT|4771,4782|false|false|false|C0879626|Adverse effects|side effect
Event|Event|SIMPLE_SEGMENT|4776,4782|false|false|false|||effect
Event|Event|SIMPLE_SEGMENT|4788,4803|false|false|false|||ANTICOAGULATION
Finding|Finding|SIMPLE_SEGMENT|4788,4803|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Finding|Physiologic Function|SIMPLE_SEGMENT|4788,4803|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4788,4803|false|false|false|C0003281|Anticoagulation Therapy|ANTICOAGULATION
Drug|Organic Chemical|SIMPLE_SEGMENT|4820,4827|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4820,4827|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|4828,4832|false|false|false|||40mg
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4855,4860|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|SIMPLE_SEGMENT|4855,4860|false|false|false|||WOUND
Finding|Body Substance|SIMPLE_SEGMENT|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|SIMPLE_SEGMENT|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|SIMPLE_SEGMENT|4855,4860|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4855,4865|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|SIMPLE_SEGMENT|4861,4865|false|false|false|C1947933|care activity|CARE
Event|Event|SIMPLE_SEGMENT|4861,4865|false|false|false|||CARE
Finding|Finding|SIMPLE_SEGMENT|4861,4865|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|4861,4865|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4886,4891|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|4886,4891|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|4886,4891|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4896,4909|false|false|false|C2937301|take a shower|take a shower
Event|Event|SIMPLE_SEGMENT|4910,4918|false|false|false|||starting
Event|Event|SIMPLE_SEGMENT|4938,4945|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|4938,4945|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4938,4945|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|4956,4960|false|false|false|||wash
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4973,4977|false|false|false|C1705308|Soap Dosage Form|soap
Event|Event|SIMPLE_SEGMENT|4973,4977|false|false|false|||soap
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4982,4987|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4982,4987|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|SIMPLE_SEGMENT|4982,4987|false|false|false|||water
Finding|Intellectual Product|SIMPLE_SEGMENT|4982,4987|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4982,4987|false|false|false|C0020311|Hydrotherapy|water
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4993,4996|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|SIMPLE_SEGMENT|4993,4996|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4993,4996|false|false|false|C2825250|Fenamole|pat
Event|Event|SIMPLE_SEGMENT|4993,4996|false|false|false|||pat
Finding|Molecular Function|SIMPLE_SEGMENT|4993,4996|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4993,4996|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5002,5010|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5002,5010|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|5002,5010|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5002,5010|false|false|false|C0184898|Surgical incisions|incision
Event|Event|SIMPLE_SEGMENT|5021,5030|false|false|false|||showering
Event|Event|SIMPLE_SEGMENT|5040,5045|true|false|false|||baths
Procedure|Health Care Activity|SIMPLE_SEGMENT|5040,5045|true|false|false|C0150141|Bathing|baths
Event|Event|SIMPLE_SEGMENT|5049,5057|true|false|false|||swimming
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5049,5057|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|SIMPLE_SEGMENT|5049,5057|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Event|Event|SIMPLE_SEGMENT|5087,5095|true|false|false|||stitches
Event|Event|SIMPLE_SEGMENT|5099,5106|true|false|false|||staples
Event|Event|SIMPLE_SEGMENT|5112,5116|true|false|false|||need
Event|Event|SIMPLE_SEGMENT|5123,5130|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|5146,5149|false|false|false|||out
Finding|Intellectual Product|SIMPLE_SEGMENT|5160,5164|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|5165,5171|false|false|false|||follow
Event|Activity|SIMPLE_SEGMENT|5175,5186|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|5175,5186|false|false|false|||appointment
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5194,5202|true|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|SIMPLE_SEGMENT|5194,5202|true|false|false|||dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5194,5202|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|5194,5202|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|5194,5202|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5194,5202|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|SIMPLE_SEGMENT|5206,5212|true|false|false|||needed
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5216,5221|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|5216,5221|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5216,5221|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|5222,5231|false|false|false|||continues
Event|Event|SIMPLE_SEGMENT|5238,5250|false|false|false|||non-draining
Event|Activity|SIMPLE_SEGMENT|5256,5264|false|false|false|C0441655|Activities|ACTIVITY
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5256,5264|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|SIMPLE_SEGMENT|5256,5264|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5269,5275|false|false|false|C0944911||WEIGHT
Event|Event|SIMPLE_SEGMENT|5269,5275|false|false|false|||WEIGHT
Finding|Finding|SIMPLE_SEGMENT|5269,5275|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Finding|Sign or Symptom|SIMPLE_SEGMENT|5269,5275|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Procedure|Health Care Activity|SIMPLE_SEGMENT|5269,5275|false|false|false|C1305866|Weighing patient|WEIGHT
Event|Event|SIMPLE_SEGMENT|5286,5291|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|5286,5291|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5286,5291|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5286,5291|false|false|false|C0152054|Therapeutic Touch|touch
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5297,5303|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|5297,5303|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|5297,5303|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|5297,5303|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|5297,5303|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|5312,5315|false|false|false|||LLE
Event|Event|SIMPLE_SEGMENT|5316,5324|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|5316,5324|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|5316,5324|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|5316,5324|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|SIMPLE_SEGMENT|5316,5332|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5316,5332|false|false|false|C0949766|Physical therapy|Physical Therapy
Event|Event|SIMPLE_SEGMENT|5325,5332|false|false|false|||Therapy
Finding|Finding|SIMPLE_SEGMENT|5325,5332|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|SIMPLE_SEGMENT|5325,5332|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5325,5332|false|false|false|C0087111|Therapeutic procedure|Therapy
Finding|Mental Process|SIMPLE_SEGMENT|5334,5339|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|Touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5334,5339|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|Touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5334,5339|false|false|false|C0152054|Therapeutic Touch|Touch
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5345,5351|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|5345,5351|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|5345,5351|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|5345,5351|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|5345,5351|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|5360,5363|false|false|false|||LLE
Event|Event|SIMPLE_SEGMENT|5364,5374|false|false|false|||Treatments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5364,5374|false|false|false|C0087111|Therapeutic procedure|Treatments
Event|Event|SIMPLE_SEGMENT|5375,5384|false|false|false|||Frequency
Finding|Intellectual Product|SIMPLE_SEGMENT|5375,5384|false|false|false|C3898838;C4321352|Frequency;How Often|Frequency
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5386,5391|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|SIMPLE_SEGMENT|5386,5391|false|false|false|||WOUND
Finding|Body Substance|SIMPLE_SEGMENT|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|SIMPLE_SEGMENT|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|SIMPLE_SEGMENT|5386,5391|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5386,5396|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|SIMPLE_SEGMENT|5392,5396|false|false|false|C1947933|care activity|CARE
Event|Event|SIMPLE_SEGMENT|5392,5396|false|false|false|||CARE
Finding|Finding|SIMPLE_SEGMENT|5392,5396|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|5392,5396|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5417,5422|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|5417,5422|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5417,5422|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5427,5440|false|false|false|C2937301|take a shower|take a shower
Event|Event|SIMPLE_SEGMENT|5441,5449|false|false|false|||starting
Event|Event|SIMPLE_SEGMENT|5469,5476|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|5469,5476|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5469,5476|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|5487,5491|false|false|false|||wash
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5504,5508|false|false|false|C1705308|Soap Dosage Form|soap
Event|Event|SIMPLE_SEGMENT|5504,5508|false|false|false|||soap
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5513,5518|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5513,5518|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|SIMPLE_SEGMENT|5513,5518|false|false|false|||water
Finding|Intellectual Product|SIMPLE_SEGMENT|5513,5518|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5513,5518|false|false|false|C0020311|Hydrotherapy|water
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5524,5527|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|SIMPLE_SEGMENT|5524,5527|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5524,5527|false|false|false|C2825250|Fenamole|pat
Event|Event|SIMPLE_SEGMENT|5524,5527|false|false|false|||pat
Finding|Molecular Function|SIMPLE_SEGMENT|5524,5527|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5524,5527|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5533,5541|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5533,5541|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|5533,5541|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5533,5541|false|false|false|C0184898|Surgical incisions|incision
Event|Event|SIMPLE_SEGMENT|5552,5561|false|false|false|||showering
Event|Event|SIMPLE_SEGMENT|5571,5576|true|false|false|||baths
Procedure|Health Care Activity|SIMPLE_SEGMENT|5571,5576|true|false|false|C0150141|Bathing|baths
Event|Event|SIMPLE_SEGMENT|5580,5588|true|false|false|||swimming
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5580,5588|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|SIMPLE_SEGMENT|5580,5588|true|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Event|Event|SIMPLE_SEGMENT|5618,5626|true|false|false|||stitches
Event|Event|SIMPLE_SEGMENT|5630,5637|true|false|false|||staples
Event|Event|SIMPLE_SEGMENT|5643,5647|true|false|false|||need
Event|Event|SIMPLE_SEGMENT|5654,5661|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|5677,5680|false|false|false|||out
Finding|Intellectual Product|SIMPLE_SEGMENT|5691,5695|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|5696,5702|false|false|false|||follow
Event|Activity|SIMPLE_SEGMENT|5706,5717|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|5706,5717|false|false|false|||appointment
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5725,5733|true|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|SIMPLE_SEGMENT|5725,5733|true|false|false|||dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5725,5733|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|5725,5733|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|5725,5733|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5725,5733|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|SIMPLE_SEGMENT|5737,5743|true|false|false|||needed
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5747,5752|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|5747,5752|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5747,5752|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|5753,5762|false|false|false|||continues
Event|Event|SIMPLE_SEGMENT|5769,5781|false|false|false|||non-draining
Procedure|Health Care Activity|SIMPLE_SEGMENT|5786,5794|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5795,5807|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|5795,5807|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5795,5807|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

