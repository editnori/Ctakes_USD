 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|false|false|false|C1717415||Allergies
Event|Event|Allergies|181,190|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|181,190|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|206,215|false|false|false|||Reactions
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|253,260|false|false|false|||dyspnea
Finding|Finding|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Classification|Chief Complaint|263,268|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|269,277|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|269,277|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,299|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|290,299|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|290,299|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|290,299|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|290,299|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|290,299|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|301,308|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Chief Complaint|301,308|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|Chief Complaint|301,324|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|Chief Complaint|301,324|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|Chief Complaint|301,324|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|Chief Complaint|301,324|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|Chief Complaint|309,324|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|309,324|false|false|false|C0007430|Catheterization|catheterization
Event|Event|History of Present Illness|381,388|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|381,391|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|392,400|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|History of Present Illness|392,400|false|false|false|||diabetes
Attribute|Clinical Attribute|History of Present Illness|402,411|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|History of Present Illness|402,415|false|false|false|C2183328|diastolic congestive heart failure|diastolic CHF
Anatomy|Body Space or Junction|History of Present Illness|412,415|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|412,415|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|History of Present Illness|412,415|false|false|false|||CHF
Disorder|Disease or Syndrome|History of Present Illness|418,430|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|418,430|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|433,436|false|true|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|433,436|false|true|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|433,436|false|true|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|433,436|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|433,436|false|true|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|433,436|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|433,436|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|433,436|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|438,465|false|false|false|C0085096|Peripheral Vascular Diseases|peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|449,457|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|History of Present Illness|449,465|false|true|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|History of Present Illness|458,465|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|458,465|false|false|false|||disease
Disorder|Disease or Syndrome|History of Present Illness|467,470|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|History of Present Illness|471,481|false|false|false|||presenting
Finding|Idea or Concept|History of Present Illness|471,481|false|false|false|C0449450|Presentation|presenting
Event|Event|History of Present Illness|511,518|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|511,518|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|511,518|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|History of Present Illness|538,543|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|538,543|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|538,543|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|538,543|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|550,556|false|false|false|||denies
Event|Event|History of Present Illness|557,563|false|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|557,563|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|565,571|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|565,571|false|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|History of Present Illness|573,578|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|573,578|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|573,583|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|573,583|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|579,583|false|false|false|C2598155||pain
Event|Event|History of Present Illness|579,583|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|579,583|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|579,583|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|585,591|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|585,591|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|585,591|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|593,601|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|593,601|true|false|false|C0042963|Vomiting|vomiting
Attribute|Clinical Attribute|History of Present Illness|608,614|false|false|false|C4255046||report
Event|Event|History of Present Illness|608,614|false|false|false|||report
Finding|Intellectual Product|History of Present Illness|608,614|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|608,614|false|false|false|C0700287|Reporting|report
Event|Event|History of Present Illness|615,622|false|false|false|||feeling
Finding|Finding|History of Present Illness|623,631|false|false|false|C2984079|Somewhat|somewhat
Event|Event|History of Present Illness|632,638|false|false|false|||wheezy
Finding|Sign or Symptom|History of Present Illness|632,638|false|false|false|C0043144|Wheezing|wheezy
Event|Event|History of Present Illness|640,646|false|false|false|||Denies
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|647,650|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|History of Present Illness|647,659|false|false|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|History of Present Illness|651,659|false|false|false|||swelling
Finding|Finding|History of Present Illness|651,659|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|651,659|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|History of Present Illness|666,674|false|false|false|C0332149|Possible|possibly
Attribute|Clinical Attribute|History of Present Illness|686,692|false|false|false|C0944911||weight
Finding|Finding|History of Present Illness|686,692|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|686,692|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|686,692|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|686,697|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Finding|Intellectual Product|History of Present Illness|686,697|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Event|Event|History of Present Illness|693,697|false|false|false|||gain
Event|Event|History of Present Illness|699,705|false|false|false|||Denies
Drug|Pharmacologic Substance|History of Present Illness|713,723|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|History of Present Illness|713,723|false|false|false|||medication
Finding|Intellectual Product|History of Present Illness|713,723|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|History of Present Illness|724,729|false|false|false|||doses
Attribute|Clinical Attribute|History of Present Illness|737,743|false|false|false|C4255046||report
Event|Event|History of Present Illness|737,743|false|false|false|||report
Finding|Intellectual Product|History of Present Illness|737,743|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|737,743|false|false|false|C0700287|Reporting|report
Event|Event|History of Present Illness|753,762|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|753,762|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|753,762|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|History of Present Illness|802,806|false|false|false|||sick
Finding|Sign or Symptom|History of Present Illness|802,806|false|false|false|C0221423|Illness (finding)|sick
Drug|Organic Chemical|History of Present Illness|814,819|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|814,819|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|814,819|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|814,819|false|false|false|C0010200|Coughing|cough
Finding|Idea or Concept|History of Present Illness|833,836|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|833,836|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|870,875|false|false|false|||lives
Finding|Finding|History of Present Illness|876,883|false|false|false|C4534363|At home|at home
Event|Event|History of Present Illness|879,883|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|879,883|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|879,883|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|879,883|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|907,923|false|false|false|||hospitalizations
Procedure|Health Care Activity|History of Present Illness|907,923|false|false|false|C0019993|Hospitalization|hospitalizations
Event|Event|History of Present Illness|927,934|false|false|false|||courses
Drug|Antibiotic|History of Present Illness|938,949|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|History of Present Illness|938,949|false|false|false|||antibiotics
Finding|Idea or Concept|History of Present Illness|963,970|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|971,977|false|false|false|||vitals
Event|Event|History of Present Illness|1006,1009|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1006,1009|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1010,1016|false|false|false|||showed
Finding|Finding|History of Present Illness|1018,1026|false|false|false|C0332148|Probable diagnosis|probable
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1027,1030|false|false|false|C1261074|Structure of right upper lobe of lung|RUL
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|1031,1034|false|true|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|History of Present Illness|1031,1034|false|false|false|||PNA
Anatomy|Cell|History of Present Illness|1043,1046|false|false|false|C0023516|Leukocytes|WBC
Drug|Organic Chemical|History of Present Illness|1051,1058|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|History of Present Illness|1051,1058|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|History of Present Illness|1051,1058|false|false|false|||lactate
Procedure|Laboratory Procedure|History of Present Illness|1051,1058|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|History of Present Illness|1060,1062|false|false|false|||Cr
Drug|Biomedical or Dental Material|History of Present Illness|1066,1074|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1066,1074|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1066,1074|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1078,1086|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|History of Present Illness|1078,1086|false|false|false|C0041199|Troponin|Troponin
Event|Event|History of Present Illness|1078,1086|false|false|false|||Troponin
Procedure|Laboratory Procedure|History of Present Illness|1078,1086|false|false|false|C0523952|Troponin measurement|Troponin
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1104,1109|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|History of Present Illness|1104,1109|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|History of Present Illness|1104,1109|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|History of Present Illness|1104,1109|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1111,1114|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|1111,1114|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|1111,1114|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|History of Present Illness|1111,1114|false|false|false|||BNP
Finding|Gene or Genome|History of Present Illness|1111,1114|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|1111,1114|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|History of Present Illness|1129,1136|false|false|false|||started
Event|Event|History of Present Illness|1141,1146|false|false|false|||bipap
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1141,1146|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|bipap
Event|Event|History of Present Illness|1154,1163|false|false|false|||tachypnea
Finding|Finding|History of Present Illness|1154,1163|false|false|false|C0231835|Tachypnea|tachypnea
Finding|Finding|History of Present Illness|1168,1177|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|History of Present Illness|1168,1177|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|History of Present Illness|1168,1195|false|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|History of Present Illness|1178,1182|false|false|false|||work
Event|Occupational Activity|History of Present Illness|1178,1182|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|History of Present Illness|1178,1195|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|History of Present Illness|1186,1195|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|1186,1195|false|false|false|||breathing
Finding|Finding|History of Present Illness|1186,1195|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|1186,1195|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|1186,1195|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|1186,1195|false|false|false|C1160636|respiratory system process|breathing
Drug|Organic Chemical|History of Present Illness|1220,1225|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|History of Present Illness|1220,1225|false|false|false|C0699992|Lasix|lasix
Event|Event|History of Present Illness|1220,1225|false|false|false|||lasix
Event|Event|History of Present Illness|1230,1237|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1241,1251|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|History of Present Illness|1241,1251|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|History of Present Illness|1241,1251|false|false|false|||vancomycin
Procedure|Laboratory Procedure|History of Present Illness|1241,1251|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|History of Present Illness|1253,1261|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|History of Present Illness|1253,1261|false|false|false|C0055003|cefepime|cefepime
Event|Event|History of Present Illness|1253,1261|false|false|false|||cefepime
Drug|Antibiotic|History of Present Illness|1267,1279|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|History of Present Illness|1267,1279|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|History of Present Illness|1267,1279|false|false|false|||levofloxacin
Event|Event|History of Present Illness|1286,1294|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1286,1294|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1286,1294|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1286,1294|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|History of Present Illness|1296,1302|false|false|false|||vitals
Event|Event|History of Present Illness|1328,1333|false|false|false|||bipap
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1328,1333|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|bipap
Event|Activity|History of Present Illness|1339,1346|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|1339,1346|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1339,1346|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|History of Present Illness|1354,1358|false|false|false|||MICU
Finding|Body Substance|History of Present Illness|1360,1367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1360,1367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1360,1367|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1368,1375|false|false|false|||reports
Event|Event|History of Present Illness|1376,1384|false|false|false|||improved
Attribute|Clinical Attribute|History of Present Illness|1385,1394|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|1385,1394|false|false|false|||breathing
Finding|Finding|History of Present Illness|1385,1394|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|1385,1394|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|1385,1394|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|1385,1394|false|false|false|C1160636|respiratory system process|breathing
Event|Event|History of Present Illness|1399,1404|false|false|false|||bipap
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1399,1404|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|bipap
Event|Event|History of Present Illness|1409,1415|false|false|false|||Review
Finding|Idea or Concept|History of Present Illness|1409,1415|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|1409,1415|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|1409,1418|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|1409,1426|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|History of Present Illness|1409,1426|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Event|Event|History of Present Illness|1419,1426|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|1419,1426|false|false|false|C0449913|System|systems
Disorder|Disease or Syndrome|History of Present Illness|1438,1441|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|1438,1441|false|false|false|||HPI
Finding|Finding|History of Present Illness|1438,1441|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|1438,1441|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Disorder|Disease or Syndrome|Past Medical History|1470,1482|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Past Medical History|1470,1482|false|false|false|||hypertension
Disorder|Disease or Syndrome|Past Medical History|1485,1493|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Past Medical History|1485,1493|false|false|false|||diabetes
Disorder|Disease or Syndrome|Past Medical History|1499,1502|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|1499,1502|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Past Medical History|1499,1502|false|false|false|||CVA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1504,1514|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1515,1524|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Past Medical History|1525,1531|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Past Medical History|1525,1531|false|false|false|||stroke
Finding|Finding|Past Medical History|1525,1531|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Past Medical History|1541,1544|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1541,1544|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|1541,1544|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|1541,1544|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|1541,1544|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|1541,1544|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|1541,1544|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1541,1544|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Past Medical History|1561,1567|false|false|false|||cathed
Disorder|Disease or Syndrome|Past Medical History|1587,1614|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1598,1606|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|Past Medical History|1598,1614|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|Past Medical History|1607,1614|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|1607,1614|false|false|false|||disease
Disorder|Disease or Syndrome|Past Medical History|1616,1628|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|Past Medical History|1616,1628|false|false|false|||claudication
Finding|Finding|Past Medical History|1616,1628|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1643,1651|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|Past Medical History|1653,1660|false|false|false|||managed
Attribute|Clinical Attribute|Past Medical History|1678,1683|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|1678,1686|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Past Medical History|1687,1690|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Past Medical History|1687,1690|false|false|false|||CKD
Drug|Biomedical or Dental Material|Past Medical History|1692,1700|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Past Medical History|1692,1700|false|false|false|||baseline
Finding|Idea or Concept|Past Medical History|1692,1700|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|1712,1716|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1712,1716|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|1717,1727|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|Past Medical History|1717,1733|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Event|Past Medical History|1728,1733|false|false|false|||rings
Event|Activity|Family Medical History|1787,1791|false|false|false|C1947906|Sorting|sort
Event|Event|Family Medical History|1787,1791|false|false|false|||sort
Finding|Cell Function|Family Medical History|1787,1791|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|Family Medical History|1787,1791|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|Family Medical History|1795,1801|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1795,1801|false|false|false|||cancer
Finding|Classification|Family Medical History|1817,1823|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|1817,1823|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|1817,1823|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|1817,1823|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|1817,1831|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|Family Medical History|1817,1834|true|false|false|C0241889|Family Medical History|family history of
Event|Event|Family Medical History|1824,1831|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|1824,1831|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1824,1831|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1824,1831|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1824,1834|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|1836,1842|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1836,1842|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1852,1857|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Family Medical History|1852,1857|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Family Medical History|1852,1857|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Family Medical History|1852,1865|false|false|false|C0018799|Heart Diseases|heart disease
Disorder|Disease or Syndrome|Family Medical History|1858,1865|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|1858,1865|false|false|false|||disease
Procedure|Health Care Activity|General Exam|1884,1893|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|1894,1898|false|false|false|||EXAM
Finding|Functional Concept|General Exam|1894,1898|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|1894,1898|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|1900,1907|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|1900,1907|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|1918,1929|false|false|false|||comfortable
Finding|Finding|General Exam|1918,1929|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|General Exam|1933,1938|false|false|false|||BiPap
Procedure|Therapeutic or Preventive Procedure|General Exam|1933,1938|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPap
Anatomy|Body Location or Region|General Exam|1939,1944|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1946,1951|false|false|false|||PERRL
Finding|Finding|General Exam|1946,1951|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|1953,1957|false|false|false|||EOMI
Anatomy|Body Location or Region|General Exam|1959,1963|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1959,1963|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1959,1963|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1965,1974|false|false|false|||difficult
Finding|Finding|General Exam|1965,1974|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|General Exam|1978,1984|false|false|false|||assess
Event|Event|General Exam|1985,1988|false|false|false|||JVP
Finding|Finding|General Exam|1985,1988|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|1996,2003|false|false|false|||habitus
Event|Event|General Exam|2008,2016|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|General Exam|2008,2016|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|General Exam|2008,2019|false|false|false|C0150312|Present|presence of
Procedure|Therapeutic or Preventive Procedure|General Exam|2021,2026|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPap
Event|Event|General Exam|2027,2032|false|false|false|||strap
Finding|Conceptual Entity|General Exam|2027,2032|false|false|false|C0935605;C1426138;C1539847;C1539888|SRFBP1 gene;STRAP gene;Strap muscle type;TTC5 gene|strap
Finding|Gene or Genome|General Exam|2027,2032|false|false|false|C0935605;C1426138;C1539847;C1539888|SRFBP1 gene;STRAP gene;Strap muscle type;TTC5 gene|strap
Event|Event|General Exam|2039,2042|false|false|false|||RRR
Event|Event|General Exam|2047,2054|false|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|2055,2060|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|2063,2067|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|General Exam|2068,2071|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|2068,2071|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|2068,2071|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|General Exam|2068,2071|false|false|false|||air
Finding|Finding|General Exam|2068,2071|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|2068,2071|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|2068,2071|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|General Exam|2072,2077|false|false|false|||entry
Finding|Functional Concept|General Exam|2072,2077|false|false|false|C1550548;C1705654|Entry (data);entry - ActRelationshipCheckpoint|entry
Finding|Intellectual Product|General Exam|2072,2077|false|false|false|C1550548;C1705654|Entry (data);entry - ActRelationshipCheckpoint|entry
Finding|Finding|General Exam|2087,2095|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|General Exam|2101,2108|false|false|false|||rhonchi
Finding|Finding|General Exam|2101,2108|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Part, Organ, or Organ Component|General Exam|2112,2115|false|false|false|C1261074|Structure of right upper lobe of lung|RUL
Event|Event|General Exam|2118,2127|false|false|false|||scattered
Finding|Organism Function|General Exam|2128,2139|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Sign or Symptom|General Exam|2128,2148|false|false|false|C0231874|Inspiratory wheezing|inspiratory wheezing
Event|Event|General Exam|2140,2148|false|false|false|||wheezing
Finding|Sign or Symptom|General Exam|2140,2148|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|General Exam|2149,2156|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2149,2156|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|2149,2156|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2159,2163|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|2159,2163|false|false|false|||soft
Disorder|Congenital Abnormality|General Exam|2170,2173|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|2170,2173|false|false|false|||Ext
Finding|Gene or Genome|General Exam|2170,2173|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Functional Concept|General Exam|2176,2181|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|General Exam|2182,2187|false|false|false|C1717255||edema
Event|Event|General Exam|2182,2187|false|false|false|||edema
Finding|Pathologic Function|General Exam|2182,2187|false|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|2189,2194|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|General Exam|2189,2194|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Organ or Tissue Function|General Exam|2195,2212|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|General Exam|2206,2212|false|false|false|C5890763||pulses
Event|Event|General Exam|2206,2212|false|false|false|||pulses
Finding|Physiologic Function|General Exam|2206,2212|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|2206,2212|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|2234,2240|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|2247,2258|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Finding|General Exam|2260,2276|false|false|false|C5425896|Mildly decreased|mildly decreased
Event|Event|General Exam|2267,2276|false|false|false|||decreased
Event|Event|General Exam|2278,2286|false|false|false|||strength
Finding|Idea or Concept|General Exam|2278,2286|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|2290,2293|false|false|false|C1261077|Structure of left lower lobe of lung|LLL
Finding|Body Substance|General Exam|2295,2304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2295,2304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2295,2304|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2295,2304|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|2305,2309|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2305,2309|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2305,2309|false|false|false|C0582103|Medical Examination|EXAM
Drug|Amino Acid, Peptide, or Protein|General Exam|2330,2333|false|false|false|C0069500|DBL Oncoprotein|P66
Drug|Biologically Active Substance|General Exam|2330,2333|false|false|false|C0069500|DBL Oncoprotein|P66
Event|Event|General Exam|2330,2333|false|false|false|||P66
Finding|Gene or Genome|General Exam|2330,2333|false|false|false|C1335821;C1427199;C1539553;C3814043|GATAD2B gene;POLD3 gene;POLD3 wt Allele;SHC1 gene|P66
Event|Event|General Exam|2351,2358|false|false|false|||GENERAL
Finding|Classification|General Exam|2351,2358|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2351,2358|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|2360,2366|false|false|false|||Laying
Disorder|Disease or Syndrome|General Exam|2370,2373|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|2370,2373|false|false|false|||bed
Finding|Intellectual Product|General Exam|2370,2373|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|General Exam|2375,2383|false|false|false|||sleeping
Finding|Intellectual Product|General Exam|2388,2393|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|2394,2402|false|false|false|||distress
Finding|Finding|General Exam|2394,2402|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2394,2402|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2406,2411|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2413,2435|false|false|false|C0517391|Moist mucous membranes|Moist mucous membranes
Finding|Body Substance|General Exam|2419,2425|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|General Exam|2419,2435|false|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|General Exam|2419,2435|false|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|General Exam|2426,2435|false|false|false|C0025255|Membrane Tissue|membranes
Anatomy|Body Location or Region|General Exam|2438,2442|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2438,2442|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2438,2442|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|2444,2450|false|false|false|||Supple
Finding|Functional Concept|General Exam|2444,2450|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|2452,2458|false|false|false|||unable
Finding|Finding|General Exam|2452,2458|false|false|false|C1299582|Unable|unable
Event|Event|General Exam|2462,2471|false|false|false|||visualize
Event|Event|General Exam|2472,2475|false|false|false|||JVP
Finding|Finding|General Exam|2472,2475|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|2477,2484|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|2477,2484|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|General Exam|2494,2498|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|2494,2498|false|false|false|||rate
Finding|Idea or Concept|General Exam|2494,2498|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|2503,2509|false|false|false|||rhythm
Finding|Finding|General Exam|2503,2509|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2503,2509|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Organ or Tissue Function|General Exam|2542,2550|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|2542,2557|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|General Exam|2551,2557|false|false|false|||murmur
Finding|Finding|General Exam|2551,2557|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|General Exam|2559,2564|false|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|2566,2571|false|false|false|||Clear
Finding|Idea or Concept|General Exam|2566,2571|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|2575,2587|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|2575,2587|false|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|2604,2612|false|false|false|||crackles
Finding|Finding|General Exam|2604,2612|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|General Exam|2614,2621|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|2614,2621|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|2624,2631|false|false|false|||rhonchi
Finding|Finding|General Exam|2624,2631|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|2635,2642|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|2635,2642|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|2635,2642|false|false|false|||ABDOMEN
Finding|Finding|General Exam|2635,2642|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|2649,2653|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|2649,2653|false|false|false|||soft
Event|Event|General Exam|2655,2667|false|false|false|||nondistended
Event|Event|General Exam|2669,2678|false|false|false|||nontender
Event|Event|General Exam|2682,2691|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|2682,2691|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|General Exam|2696,2707|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|2709,2713|false|false|false|||Warm
Finding|Finding|General Exam|2709,2713|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2709,2713|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2718,2722|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2723,2731|false|false|false|||perfused
Drug|Food|General Exam|2733,2739|false|false|false|C5890763||Pulses
Event|Event|General Exam|2733,2739|false|false|false|||Pulses
Finding|Physiologic Function|General Exam|2733,2739|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|General Exam|2733,2739|false|false|false|C0034107|Pulse taking|Pulses
Finding|Functional Concept|General Exam|2744,2749|false|false|false|C1883002|Sequence Chromatogram|Trace
Attribute|Clinical Attribute|General Exam|2762,2767|false|false|false|C1717255||edema
Event|Event|General Exam|2762,2767|false|false|false|||edema
Finding|Pathologic Function|General Exam|2762,2767|false|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|General Exam|2794,2803|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|General Exam|2818,2823|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2818,2823|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2818,2823|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2824,2827|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2832,2835|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2832,2835|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2832,2835|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2842,2845|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2842,2845|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2842,2845|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2842,2845|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2851,2854|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2851,2854|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2862,2865|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2862,2865|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2862,2865|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2862,2865|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2862,2865|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2869,2872|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2869,2872|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2869,2872|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2869,2872|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2869,2872|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2869,2872|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|2879,2883|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2898,2901|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2918,2923|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2918,2923|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2918,2923|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|2939,2944|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|2939,2944|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|2939,2944|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|2949,2952|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|2949,2952|false|false|false|||Eos
Finding|Gene or Genome|General Exam|2949,2952|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|2979,2984|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2979,2984|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2979,2984|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2989,2992|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|2989,2992|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|2989,2992|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3015,3020|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3015,3020|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3015,3020|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3015,3028|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3015,3028|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3015,3028|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3021,3028|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3021,3028|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3021,3028|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3021,3028|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3021,3028|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3021,3028|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3075,3079|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3075,3079|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3075,3079|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3105,3110|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3105,3110|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3105,3110|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3111,3116|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3111,3116|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3111,3116|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3111,3116|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|3114,3118|false|false|false|C4722362|MB-6|MB-6
Drug|Amino Acid, Peptide, or Protein|General Exam|3119,3125|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|3119,3125|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|3144,3149|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3144,3149|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3144,3149|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3176,3181|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3176,3181|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3176,3181|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3182,3187|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3182,3187|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3182,3187|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3182,3187|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|3216,3221|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3216,3221|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3216,3221|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3216,3229|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|3222,3229|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|3222,3229|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|General Exam|3222,3229|false|false|false|||Lactate
Procedure|Laboratory Procedure|General Exam|3222,3229|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|General Exam|3246,3251|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|3246,3251|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|3246,3251|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|3246,3257|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|3252,3257|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3252,3257|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|General Exam|3258,3263|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|General Exam|3271,3276|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|3296,3301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|3296,3301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|3296,3301|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|3296,3307|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|3302,3307|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|3302,3307|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|3308,3311|false|false|false|||NEG
Finding|Finding|General Exam|3308,3311|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|3312,3319|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|3312,3319|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|3312,3319|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|General Exam|3320,3323|false|false|false|||NEG
Finding|Finding|General Exam|3320,3323|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|3324,3331|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|3324,3331|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|3324,3331|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|3324,3331|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|3324,3331|false|false|false|C0202202|Protein measurement|Protein
Event|Event|General Exam|3332,3335|false|false|false|||NEG
Finding|Finding|General Exam|3332,3335|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|3337,3344|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3337,3344|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3337,3344|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3337,3344|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3337,3344|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3337,3344|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|3345,3348|false|false|false|||NEG
Finding|Finding|General Exam|3345,3348|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|3349,3355|false|false|false|C0022634|Ketones|Ketone
Event|Event|General Exam|3356,3359|false|false|false|||NEG
Finding|Finding|General Exam|3356,3359|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|3368,3371|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|3380,3383|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|3397,3400|false|false|false|||NEG
Finding|Finding|General Exam|3397,3400|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|3405,3414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3405,3414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3405,3414|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3405,3414|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|3429,3434|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3429,3434|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3429,3434|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3435,3438|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3443,3446|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3443,3446|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3443,3446|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3453,3456|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3453,3456|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3453,3456|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3453,3456|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3462,3465|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3462,3465|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3473,3476|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3473,3476|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3473,3476|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3473,3476|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3473,3476|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3480,3483|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3480,3483|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3480,3483|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3480,3483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3480,3483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3480,3483|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|3489,3493|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|3489,3493|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3508,3511|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3528,3533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3528,3533|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3528,3533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3528,3541|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3528,3541|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3528,3541|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3534,3541|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3534,3541|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3534,3541|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3534,3541|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3534,3541|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3534,3541|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3589,3593|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3589,3593|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3589,3593|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3618,3623|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3618,3623|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3618,3623|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3618,3631|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3624,3631|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3624,3631|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3624,3631|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3624,3631|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3624,3631|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3624,3631|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3624,3631|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3624,3631|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|General Exam|3654,3657|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|3654,3657|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Functional Concept|General Exam|3663,3668|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|3663,3679|false|false|false|C1261074|Structure of right upper lobe of lung|Right upper lobe
Disorder|Disease or Syndrome|General Exam|3663,3689|false|false|false|C0585106|Right upper zone pneumonia|Right upper lobe pneumonia
Anatomy|Body Part, Organ, or Organ Component|General Exam|3669,3679|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|3675,3679|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|3675,3679|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|General Exam|3680,3689|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|3680,3689|false|false|false|||pneumonia
Event|Event|General Exam|3693,3697|false|false|false|||mass
Finding|Finding|General Exam|3693,3697|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|3693,3697|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3693,3697|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Functional Concept|General Exam|3715,3720|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|3728,3736|false|false|false|||fullness
Finding|Finding|General Exam|3738,3744|false|false|false|C0577559|Mass of body structure|a mass
Event|Event|General Exam|3740,3744|false|false|false|||mass
Finding|Finding|General Exam|3740,3744|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|3740,3744|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3740,3744|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|General Exam|3745,3754|false|false|false|||resulting
Disorder|Disease or Syndrome|General Exam|3775,3784|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|3801,3813|false|false|false|||differential
Finding|Idea or Concept|General Exam|3801,3813|false|false|false|C1549478|Amount type - Differential|differential
Anatomy|Body Location or Region|General Exam|3826,3831|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|3826,3831|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|General Exam|3826,3834|false|false|false|C0202823|Chest CT|chest CT
Event|Event|General Exam|3832,3834|false|false|false|||CT
Procedure|Diagnostic Procedure|General Exam|3832,3860|false|false|false|C0202653|CT with intravenous contrast|CT with intravenous contrast
Finding|Functional Concept|General Exam|3840,3851|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3840,3860|false|false|false|C4072741|IV contrast|intravenous contrast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3852,3860|false|false|false|C0009924|Contrast Media|contrast
Event|Event|General Exam|3852,3860|false|false|false|||contrast
Event|Activity|General Exam|3875,3885|false|false|false|C1516048|Assessed|assessment
Event|Event|General Exam|3875,3885|false|false|false|||assessment
Finding|Intellectual Product|General Exam|3875,3885|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|General Exam|3875,3885|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|General Exam|3875,3885|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Event|Event|General Exam|3889,3892|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|3889,3892|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|General Exam|3902,3906|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3902,3913|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|General Exam|3907,3913|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|General Exam|3917,3926|false|false|false|||elongated
Finding|Intellectual Product|General Exam|3937,3941|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Conceptual Entity|General Exam|3942,3951|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3942,3951|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Functional Concept|General Exam|3952,3956|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3958,3969|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|General Exam|3958,3981|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|General Exam|3970,3981|false|false|false|||hypertrophy
Finding|Pathologic Function|General Exam|3970,3981|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Body Space or Junction|General Exam|3994,4000|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|3994,4000|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|3994,4000|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|General Exam|4001,4005|false|false|false|||size
Finding|Intellectual Product|General Exam|4016,4020|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|General Exam|4025,4033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4025,4033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|General Exam|4043,4047|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|General Exam|4043,4080|false|false|false|C1277187|Left ventricular systolic dysfunction|left ventricular systolic dysfunction
Anatomy|Body Part, Organ, or Organ Component|General Exam|4048,4059|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|4060,4068|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|4060,4080|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|4069,4080|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|4069,4080|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|4069,4080|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|4069,4080|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|4069,4080|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Social Behavior|General Exam|4108,4116|false|false|false|C0678975|inferiority|inferior
Event|Event|General Exam|4151,4159|false|false|false|||segments
Event|Event|General Exam|4175,4183|false|false|false|||segments
Event|Event|General Exam|4184,4192|false|false|false|||contract
Attribute|Clinical Attribute|General Exam|4203,4207|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|General Exam|4203,4207|false|false|false|||LVEF
Procedure|Diagnostic Procedure|General Exam|4203,4207|false|false|false|C3837267|LVEF (procedure)|LVEF
Finding|Functional Concept|General Exam|4220,4225|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4226,4237|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|4238,4245|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|General Exam|4255,4259|false|false|false|||free
Finding|Functional Concept|General Exam|4255,4259|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|General Exam|4260,4271|false|false|false|C1980023|Wall motion|wall motion
Event|Event|General Exam|4265,4271|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|General Exam|4265,4271|false|false|false|C0026597|Motion|motion
Event|Event|General Exam|4277,4283|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|4289,4295|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4289,4301|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|4296,4301|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|4302,4310|false|false|false|||leaflets
Event|Event|General Exam|4326,4335|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|General Exam|4341,4347|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|General Exam|4341,4356|true|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|General Exam|4348,4356|false|false|false|||stenosis
Finding|Pathologic Function|General Exam|4348,4356|false|false|false|C1261287|Stenosis|stenosis
Event|Event|General Exam|4364,4371|false|false|false|||present
Finding|Finding|General Exam|4364,4371|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|4364,4371|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|General Exam|4376,4382|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|General Exam|4376,4396|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|General Exam|4383,4396|false|false|false|||regurgitation
Finding|Finding|General Exam|4383,4396|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4383,4396|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4383,4396|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4400,4404|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|General Exam|4411,4423|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|4418,4423|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|4424,4432|false|false|false|||leaflets
Event|Event|General Exam|4444,4453|false|false|false|||thickened
Disorder|Disease or Syndrome|General Exam|4468,4471|false|false|false|C0039235|Tachycardia, Ectopic Junctional|jet
Event|Event|General Exam|4468,4471|false|false|false|||jet
Finding|Gene or Genome|General Exam|4468,4471|false|false|false|C1539482|FBXL15 gene|jet
Event|Event|General Exam|4476,4484|false|false|false|||moderate
Finding|Finding|General Exam|4476,4484|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4476,4484|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|General Exam|4488,4494|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|4488,4494|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|General Exam|4500,4520|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|4507,4520|false|false|false|||regurgitation
Finding|Finding|General Exam|4507,4520|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4507,4520|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4507,4520|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4524,4528|false|false|false|||seen
Finding|Finding|General Exam|4540,4548|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4540,4548|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Part, Organ, or Organ Component|General Exam|4549,4558|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|4549,4558|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|4549,4558|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4549,4565|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|4559,4565|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|4559,4565|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|4566,4574|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|General Exam|4566,4587|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|General Exam|4575,4587|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|4575,4587|false|false|false|||hypertension
Anatomy|Body Location or Region|General Exam|4602,4613|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4602,4613|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|General Exam|4602,4622|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|General Exam|4602,4622|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|General Exam|4614,4622|false|false|false|||effusion
Finding|Body Substance|General Exam|4614,4622|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|4614,4622|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|4614,4622|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|General Exam|4625,4635|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|4625,4635|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|4625,4635|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|General Exam|4637,4641|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|General Exam|4645,4653|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4645,4653|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|General Exam|4663,4667|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4668,4679|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|General Exam|4680,4688|false|false|false|||systolic
Finding|Organ or Tissue Function|General Exam|4680,4688|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|General Exam|4690,4701|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|4690,4701|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|4690,4701|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|4690,4701|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|4690,4701|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Disorder|Disease or Syndrome|General Exam|4707,4710|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|General Exam|4707,4710|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|General Exam|4707,4710|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|General Exam|4707,4710|false|false|false|||CAD
Finding|Gene or Genome|General Exam|4707,4710|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|General Exam|4707,4710|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|General Exam|4707,4710|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|General Exam|4707,4710|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|General Exam|4712,4720|false|false|false|||Moderate
Finding|Finding|General Exam|4712,4720|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|4712,4720|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Finding|General Exam|4724,4730|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|4724,4730|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|General Exam|4724,4751|false|false|false|C5393153|Severe mitral regurgitation|severe mitral regurgitation
Disorder|Disease or Syndrome|General Exam|4731,4751|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|4738,4751|false|false|false|||regurgitation
Finding|Finding|General Exam|4738,4751|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4738,4751|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4738,4751|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Finding|General Exam|4754,4762|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|4754,4762|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Pathologic Function|General Exam|4754,4785|false|false|false|C5395246|Moderate pulmonary hypertension|Moderate pulmonary hypertension
Anatomy|Body Part, Organ, or Organ Component|General Exam|4763,4772|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|4763,4772|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|4763,4772|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|4763,4785|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|General Exam|4773,4785|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|4773,4785|false|false|false|||hypertension
Event|Event|General Exam|4812,4817|false|false|false|||study
Finding|Intellectual Product|General Exam|4812,4817|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|4812,4817|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|General Exam|4826,4834|false|false|false|||reviewed
Lab|Laboratory or Test Result|General Exam|4854,4868|false|false|false|C0455816|Left ventricular wall motion|LV wall motion
Attribute|Clinical Attribute|General Exam|4857,4868|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|General Exam|4862,4868|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|General Exam|4869,4882|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|4869,4882|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|4869,4882|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|4887,4890|false|false|false|||new
Finding|Finding|General Exam|4887,4890|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|4887,4890|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|General Exam|4905,4925|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|4912,4925|false|false|false|||regurgitation
Finding|Finding|General Exam|4912,4925|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4912,4925|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4912,4925|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4930,4939|false|false|false|||increased
Anatomy|Body Part, Organ, or Organ Component|General Exam|4942,4949|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4942,4949|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Diagnostic Procedure|General Exam|4942,4954|false|false|false|C0018795|Cardiac Catheterization Procedures|CARDIAC CATH
Event|Event|General Exam|4950,4954|false|false|false|||CATH
Procedure|Therapeutic or Preventive Procedure|General Exam|4950,4954|false|false|false|C0007430|Catheterization|CATH
Anatomy|Body Part, Organ, or Organ Component|General Exam|4973,4981|false|false|false|C0018787|Heart|coronary
Procedure|Diagnostic Procedure|General Exam|4973,4993|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Procedure|Health Care Activity|General Exam|4973,4993|false|false|false|C0085532;C1548829|Consent Type - Coronary Angiography;Coronary angiography|coronary angiography
Event|Event|General Exam|4982,4993|false|false|false|||angiography
Procedure|Diagnostic Procedure|General Exam|4982,4993|false|false|false|C0002978|angiogram|angiography
Finding|Functional Concept|General Exam|5002,5007|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|General Exam|5008,5016|false|false|false|C1527180|Dominant|dominant
Drug|Biomedical or Dental Material|General Exam|5017,5023|false|false|false|C5671121|System (basic dose form)|system
Event|Event|General Exam|5017,5023|false|false|false|||system
Finding|Functional Concept|General Exam|5017,5023|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Event|General Exam|5025,5033|false|false|false|||revealed
Anatomy|Body Location or Region|General Exam|5040,5046|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|General Exam|5040,5046|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|General Exam|5040,5055|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5047,5055|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5047,5062|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|General Exam|5047,5070|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|General Exam|5056,5062|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5056,5062|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|General Exam|5056,5070|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|General Exam|5063,5070|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5063,5070|false|false|false|||disease
Drug|Organic Chemical|General Exam|5077,5081|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Pharmacologic Substance|General Exam|5077,5081|false|false|false|C2828271|levomefolate calcium|LMCA
Drug|Vitamin|General Exam|5077,5081|false|false|false|C2828271|levomefolate calcium|LMCA
Finding|Functional Concept|General Exam|5090,5101|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|General Exam|5090,5109|false|false|false|C0746982|obstructive disease|obstructive disease
Disorder|Disease or Syndrome|General Exam|5102,5109|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5102,5109|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|General Exam|5116,5119|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|5116,5119|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|5116,5119|false|false|false|||LAD
Finding|Gene or Genome|General Exam|5116,5119|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|General Exam|5126,5134|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|5126,5134|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|General Exam|5126,5142|false|false|false|C4740691|Moderate disease|moderate disease
Disorder|Disease or Syndrome|General Exam|5135,5142|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5135,5142|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|General Exam|5155,5161|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5155,5161|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Drug|Chemical Viewed Structurally|General Exam|5177,5183|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|General Exam|5177,5183|false|false|false|||branch
Attribute|Clinical Attribute|General Exam|5195,5203|false|false|false|C4489236|Proximal Resection Margin|proximal
Event|Event|General Exam|5204,5210|false|false|false|||lesion
Finding|Finding|General Exam|5204,5210|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|5204,5210|false|false|false|C0221198;C1546698|Lesion|lesion
Drug|Amino Acid, Peptide, or Protein|General Exam|5218,5221|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|Lcx
Drug|Enzyme|General Exam|5218,5221|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|Lcx
Finding|Gene or Genome|General Exam|5218,5221|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|Lcx
Attribute|Clinical Attribute|General Exam|5232,5240|false|false|false|C4489236|Proximal Resection Margin|proximal
Event|Event|General Exam|5241,5247|false|false|false|||lesion
Finding|Finding|General Exam|5241,5247|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|5241,5247|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|General Exam|5254,5257|false|false|false|||RCA
Finding|Finding|General Exam|5262,5269|false|false|false|C4699603|Totally|totally
Event|Event|General Exam|5270,5278|false|false|false|||occluded
Finding|Finding|General Exam|5270,5278|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|General Exam|5270,5278|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Anatomy|Body Location or Region|Final Diagnosis|5327,5333|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5327,5333|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5327,5342|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5334,5342|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5334,5349|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Final Diagnosis|5334,5357|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5343,5349|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Final Diagnosis|5343,5349|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Final Diagnosis|5343,5357|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Final Diagnosis|5350,5357|false|false|false|C0012634|Disease|disease
Event|Event|Final Diagnosis|5350,5357|false|false|false|||disease
Procedure|Therapeutic or Preventive Procedure|Final Diagnosis|5373,5377|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|Final Diagnosis|5378,5388|false|false|false|||evaluation
Finding|Idea or Concept|Final Diagnosis|5378,5388|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Final Diagnosis|5378,5388|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Attribute|Clinical Attribute|Final Diagnosis|5390,5398|false|false|false|C0881858||CT CHEST
Procedure|Diagnostic Procedure|Final Diagnosis|5390,5398|false|false|false|C0202823|Chest CT|CT CHEST
Anatomy|Body Location or Region|Final Diagnosis|5393,5398|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Final Diagnosis|5393,5398|false|false|false|C0741025|Chest problem|CHEST
Finding|Finding|Final Diagnosis|5426,5448|false|false|false|C5539411|Ground glass opacity|ground-glass opacities
Disorder|Disease or Syndrome|Final Diagnosis|5433,5438|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|Final Diagnosis|5433,5438|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|Final Diagnosis|5433,5438|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|Final Diagnosis|5433,5438|false|false|false|C0025611|methamphetamine|glass
Event|Event|Final Diagnosis|5439,5448|false|false|false|||opacities
Finding|Finding|Final Diagnosis|5439,5448|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|Final Diagnosis|5439,5448|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Functional Concept|Final Diagnosis|5471,5476|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5471,5487|false|false|false|C1261074|Structure of right upper lobe of lung|right upper lobe
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5477,5487|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5483,5487|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Final Diagnosis|5483,5487|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Functional Concept|Final Diagnosis|5492,5497|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5492,5508|false|false|false|C1261075|Structure of right lower lobe of lung|right lower lobe
Anatomy|Body Location or Region|Final Diagnosis|5498,5503|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Final Diagnosis|5498,5503|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5498,5508|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5504,5508|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Final Diagnosis|5504,5508|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Idea or Concept|Final Diagnosis|5509,5520|false|false|false|C0750501|most likely|most likely
Finding|Finding|Final Diagnosis|5514,5520|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Final Diagnosis|5514,5520|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Activity|Final Diagnosis|5521,5530|false|true|false|C1882932|Representation (action)|represent
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5541,5550|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Final Diagnosis|5541,5550|false|false|false|C2707265||pulmonary
Finding|Finding|Final Diagnosis|5541,5550|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Final Diagnosis|5541,5556|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Final Diagnosis|5551,5556|false|false|false|C1717255||edema
Event|Event|Final Diagnosis|5551,5556|false|false|false|||edema
Finding|Pathologic Function|Final Diagnosis|5551,5556|false|false|false|C0013604|Edema|edema
Finding|Pathologic Function|Final Diagnosis|5551,5567|false|false|false|C0013609|Localized Edema|edema, localized
Event|Event|Final Diagnosis|5558,5567|false|false|false|||localized
Finding|Functional Concept|Final Diagnosis|5575,5580|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5575,5585|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|Final Diagnosis|5581,5585|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5581,5585|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Final Diagnosis|5581,5585|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Final Diagnosis|5581,5585|false|false|false|C0740941|Lung Problem|lung
Event|Event|Final Diagnosis|5598,5607|false|false|false|||direction
Finding|Idea or Concept|Final Diagnosis|5598,5607|false|false|false|C1550715|direction - AddressPartType|direction
Disorder|Disease or Syndrome|Final Diagnosis|5611,5614|false|false|false|C0039235|Tachycardia, Ectopic Junctional|jet
Event|Event|Final Diagnosis|5611,5614|false|false|false|||jet
Finding|Gene or Genome|Final Diagnosis|5611,5614|false|false|false|C1539482|FBXL15 gene|jet
Event|Event|Final Diagnosis|5626,5639|false|false|false|||regurgitation
Finding|Finding|Final Diagnosis|5626,5639|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Final Diagnosis|5626,5639|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Final Diagnosis|5626,5639|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Finding|Final Diagnosis|5647,5655|false|false|false|C0332149|Possible|Possible
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5656,5665|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Final Diagnosis|5656,5665|false|false|false|C2707265||pulmonary
Finding|Finding|Final Diagnosis|5656,5665|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Final Diagnosis|5656,5678|false|true|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|Final Diagnosis|5666,5678|false|true|false|C0020538|Hypertensive disease|hypertension
Event|Event|Final Diagnosis|5666,5678|false|false|false|||hypertension
Finding|Finding|Final Diagnosis|5685,5693|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Final Diagnosis|5685,5693|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5694,5702|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5694,5709|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Final Diagnosis|5694,5717|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5703,5709|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Final Diagnosis|5703,5709|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Final Diagnosis|5703,5717|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Final Diagnosis|5710,5717|false|false|false|C0012634|Disease|disease
Event|Event|Final Diagnosis|5710,5717|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5721,5728|false|false|false|C0007272|Carotid Arteries|CAROTID
Event|Event|Final Diagnosis|5740,5748|false|false|false|||evidence
Finding|Idea or Concept|Final Diagnosis|5740,5748|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Final Diagnosis|5740,5751|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|Final Diagnosis|5768,5779|true|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5780,5796|false|false|false|C0741978|carotid internal|internal carotid
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5789,5796|false|false|false|C0007272|Carotid Arteries|carotid
Event|Event|Final Diagnosis|5798,5806|false|false|false|||stenosis
Finding|Pathologic Function|Final Diagnosis|5798,5806|false|false|false|C1261287|Stenosis|stenosis
Event|Event|Final Diagnosis|5825,5829|false|false|false|||ECHO
Procedure|Health Care Activity|Final Diagnosis|5825,5829|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Final Diagnosis|5825,5829|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Drug|Amino Acid, Peptide, or Protein|Final Diagnosis|5835,5838|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Final Diagnosis|5835,5838|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|Final Diagnosis|5835,5838|false|false|false|||PCI
Finding|Gene or Genome|Final Diagnosis|5835,5838|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Final Diagnosis|5835,5838|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Final Diagnosis|5835,5838|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Finding|Intellectual Product|Final Diagnosis|5849,5853|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Conceptual Entity|Final Diagnosis|5854,5863|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|Final Diagnosis|5854,5863|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Functional Concept|Final Diagnosis|5864,5868|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|Final Diagnosis|5864,5892|false|false|false|C3484363||left ventricular hypertrophy
Disorder|Disease or Syndrome|Final Diagnosis|5864,5892|false|false|false|C0149721|Left Ventricular Hypertrophy|left ventricular hypertrophy
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5869,5880|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|Final Diagnosis|5869,5892|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|Final Diagnosis|5881,5892|false|false|false|||hypertrophy
Finding|Pathologic Function|Final Diagnosis|5881,5892|false|false|false|C0020564|Hypertrophy|hypertrophy
Event|Event|Final Diagnosis|5898,5904|false|false|false|||normal
Anatomy|Body Space or Junction|Final Diagnosis|5906,5912|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Final Diagnosis|5906,5912|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Final Diagnosis|5906,5912|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|Final Diagnosis|5913,5917|false|false|false|||size
Finding|Intellectual Product|Final Diagnosis|5928,5932|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|Final Diagnosis|5942,5946|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|5947,5958|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|Final Diagnosis|5959,5967|false|false|false|||systolic
Finding|Organ or Tissue Function|Final Diagnosis|5959,5967|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Final Diagnosis|5969,5980|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Final Diagnosis|5969,5980|false|false|false|||dysfunction
Finding|Conceptual Entity|Final Diagnosis|5969,5980|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Final Diagnosis|5969,5980|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Final Diagnosis|5969,5980|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|Final Diagnosis|5986,5994|false|false|false|||inferior
Finding|Social Behavior|Final Diagnosis|5986,5994|false|false|false|C0678975|inferiority|inferior
Event|Event|Final Diagnosis|6014,6025|false|false|false|||hypokinesis
Finding|Finding|Final Diagnosis|6014,6025|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|Final Diagnosis|6031,6037|false|false|false|||masses
Event|Event|Final Diagnosis|6041,6048|false|false|false|||thrombi
Finding|Pathologic Function|Final Diagnosis|6041,6048|false|false|false|C0087086|Thrombus|thrombi
Event|Event|Final Diagnosis|6053,6057|false|false|false|||seen
Finding|Functional Concept|Final Diagnosis|6065,6069|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6065,6079|false|false|false|C0225897;C4266612|Chest>Heart.ventricle.left;Left ventricular structure|left ventricle
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6070,6079|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|Final Diagnosis|6070,6079|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6094,6105|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|Final Diagnosis|6094,6119|false|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|Final Diagnosis|6106,6119|false|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|Final Diagnosis|6106,6119|false|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|Final Diagnosis|6113,6119|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|Final Diagnosis|6113,6119|false|false|false|||defect
Finding|Functional Concept|Final Diagnosis|6113,6119|false|false|false|C1457869|Defect|defect
Finding|Functional Concept|Final Diagnosis|6121,6126|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6127,6138|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6139,6146|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|Final Diagnosis|6157,6161|false|false|false|||free
Finding|Functional Concept|Final Diagnosis|6157,6161|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|Final Diagnosis|6162,6173|false|false|false|C1980023|Wall motion|wall motion
Event|Event|Final Diagnosis|6167,6173|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|Final Diagnosis|6167,6173|false|false|false|C0026597|Motion|motion
Event|Event|Final Diagnosis|6178,6184|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6190,6202|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6197,6202|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Final Diagnosis|6203,6211|false|false|false|||leaflets
Event|Event|Final Diagnosis|6224,6233|false|false|false|||thickened
Disorder|Disease or Syndrome|Final Diagnosis|6248,6251|false|false|false|C0039235|Tachycardia, Ectopic Junctional|jet
Event|Event|Final Diagnosis|6248,6251|false|false|false|||jet
Finding|Gene or Genome|Final Diagnosis|6248,6251|false|false|false|C1539482|FBXL15 gene|jet
Finding|Intellectual Product|Final Diagnosis|6255,6259|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Final Diagnosis|6273,6286|false|false|false|||regurgitation
Finding|Finding|Final Diagnosis|6273,6286|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Final Diagnosis|6273,6286|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Final Diagnosis|6273,6286|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Final Diagnosis|6290,6294|false|false|false|||seen
Anatomy|Body Location or Region|Final Diagnosis|6308,6319|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Final Diagnosis|6308,6319|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Final Diagnosis|6308,6328|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Final Diagnosis|6308,6328|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|Final Diagnosis|6320,6328|false|false|false|||effusion
Finding|Body Substance|Final Diagnosis|6320,6328|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Final Diagnosis|6320,6328|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Final Diagnosis|6320,6328|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|Final Diagnosis|6356,6361|false|false|false|||study
Finding|Intellectual Product|Final Diagnosis|6356,6361|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Final Diagnosis|6356,6361|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|Final Diagnosis|6370,6378|false|false|false|||reviewed
Attribute|Clinical Attribute|Final Diagnosis|6393,6397|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|Final Diagnosis|6393,6397|false|false|false|||LVEF
Procedure|Diagnostic Procedure|Final Diagnosis|6393,6397|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|Final Diagnosis|6402,6411|false|false|false|||increased
Event|Event|Final Diagnosis|6417,6423|false|false|false|||degree
Finding|Intellectual Product|Final Diagnosis|6417,6423|false|false|false|C0542560|Academic degree|degree
Event|Event|Final Diagnosis|6430,6434|false|false|false|||seen
Event|Event|Final Diagnosis|6439,6448|false|false|false|||decreased
Disorder|Disease or Syndrome|Hospital Course|6498,6501|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|6498,6501|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|6503,6511|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Hospital Course|6503,6511|false|false|false|||diabetes
Disorder|Disease or Syndrome|Hospital Course|6513,6516|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Hospital Course|6513,6516|false|false|false|||CKD
Event|Event|Hospital Course|6517,6526|false|false|false|||presented
Event|Event|Hospital Course|6543,6550|false|false|false|||dyspnea
Finding|Finding|Hospital Course|6543,6550|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|6543,6550|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|Hospital Course|6570,6575|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|6570,6575|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|6570,6575|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|6570,6575|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|6584,6590|false|false|false|||fevers
Finding|Sign or Symptom|Hospital Course|6584,6590|true|false|false|C0015967|Fever|fevers
Event|Event|Hospital Course|6610,6615|false|false|false|||count
Event|Event|Hospital Course|6627,6635|false|false|false|||admitted
Event|Event|Hospital Course|6648,6655|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|6648,6655|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|6661,6670|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|6661,6670|false|false|false|||pneumonia
Event|Event|Hospital Course|6685,6690|false|false|false|||found
Event|Event|Hospital Course|6702,6709|false|false|false|||changes
Finding|Functional Concept|Hospital Course|6702,6709|false|false|false|C0392747|Changing|changes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6711,6717|false|false|false|C0014442;C5399708|Enzyme [APC];Enzymes|enzyme
Drug|Enzyme|Hospital Course|6711,6717|false|false|false|C0014442;C5399708|Enzyme [APC];Enzymes|enzyme
Event|Event|Hospital Course|6711,6717|false|false|false|||enzyme
Event|Event|Hospital Course|6719,6723|false|false|false|||leak
Finding|Functional Concept|Hospital Course|6719,6723|false|false|false|C0332234|Leaking|leak
Finding|Finding|Hospital Course|6725,6728|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6725,6728|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|Hospital Course|6729,6740|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|Hospital Course|6734,6740|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|Hospital Course|6741,6752|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Hospital Course|6741,6752|false|false|false|||abnormality
Finding|Finding|Hospital Course|6741,6752|false|false|false|C1704258|Abnormality|abnormality
Event|Event|Hospital Course|6753,6763|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|6753,6763|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|6753,6768|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6779,6786|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|6779,6786|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|Hospital Course|6779,6792|false|false|false|C0741923|Cardiac Events|cardiac event
Event|Event|Hospital Course|6787,6792|false|false|false|||event
Event|Event|Hospital Course|6787,6792|false|false|false|C0441471|Event|event
Event|Event|Hospital Course|6804,6812|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|6804,6812|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|6804,6815|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Hospital Course|6816,6825|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|6816,6825|false|false|false|||pneumonia
Event|Event|Hospital Course|6830,6836|false|false|false|||fevers
Finding|Sign or Symptom|Hospital Course|6830,6836|true|false|false|C0015967|Fever|fevers
Anatomy|Cell|Hospital Course|6838,6841|false|false|false|C0023516|Leukocytes|wbc
Drug|Organic Chemical|Hospital Course|6844,6851|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|Hospital Course|6844,6851|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|Hospital Course|6844,6851|false|false|false|||lactate
Procedure|Laboratory Procedure|Hospital Course|6844,6851|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|Hospital Course|6860,6866|false|false|false|||vitals
Event|Event|Hospital Course|6868,6871|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|6868,6871|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|Hospital Course|6877,6883|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6877,6883|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6894,6903|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6894,6903|false|true|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6894,6903|false|true|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|Hospital Course|6905,6910|false|false|false|C1717255||edema
Event|Event|Hospital Course|6905,6910|false|false|false|||edema
Finding|Pathologic Function|Hospital Course|6905,6910|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|Hospital Course|6916,6936|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Hospital Course|6923,6936|false|false|false|||regurgitation
Finding|Finding|Hospital Course|6923,6936|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|6923,6936|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|6923,6936|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Hospital Course|6947,6951|false|false|false|||seen
Anatomy|Body System|Hospital Course|6955,6965|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Hospital Course|6971,6982|false|false|false|||transferred
Finding|Body Substance|Hospital Course|6987,6994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6987,6994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6987,6994|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body System|Hospital Course|6998,7008|false|false|false|C0007226|Cardiovascular system|cardiology
Anatomy|Anatomical Structure|Hospital Course|7009,7014|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Intellectual Product|Hospital Course|7019,7024|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|7019,7037|false|false|false|C4083073|acute systolic congestive heart failure|Acute systolic CHF
Finding|Organ or Tissue Function|Hospital Course|7025,7033|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Hospital Course|7025,7037|false|false|false|C2039715|systolic congestive heart failure|systolic CHF
Anatomy|Body Space or Junction|Hospital Course|7034,7037|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|7034,7037|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|7038,7050|false|false|false|||exacerbation
Finding|Finding|Hospital Course|7038,7050|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Disease or Syndrome|Hospital Course|7051,7071|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Hospital Course|7058,7071|false|false|false|||regurgitation
Finding|Finding|Hospital Course|7058,7071|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|7058,7071|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|7058,7071|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Finding|Hospital Course|7074,7080|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|7074,7080|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Disorder|Neoplastic Process|Hospital Course|7081,7090|false|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|7081,7090|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|7081,7090|false|true|false|C1522484|metastatic qualifier|secondary
Finding|Functional Concept|Hospital Course|7094,7102|false|true|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|Hospital Course|7103,7119|false|false|false|C3258293|Valvular disease|valvular disease
Disorder|Disease or Syndrome|Hospital Course|7112,7119|false|true|false|C0012634|Disease|disease
Event|Event|Hospital Course|7112,7119|false|false|false|||disease
Event|Event|Hospital Course|7120,7129|false|false|false|||resulting
Disorder|Disease or Syndrome|Hospital Course|7144,7164|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Hospital Course|7151,7164|false|false|false|||regurgitation
Finding|Finding|Hospital Course|7151,7164|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|7151,7164|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|7151,7164|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Hospital Course|7166,7170|false|false|false|||ECHO
Procedure|Health Care Activity|Hospital Course|7166,7170|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7166,7170|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|Hospital Course|7181,7189|false|false|false|C0233568|Akinetic|akinetic
Event|Event|Hospital Course|7190,7198|false|false|false|||inferior
Finding|Social Behavior|Hospital Course|7190,7198|false|false|false|C0678975|inferiority|inferior
Event|Event|Hospital Course|7205,7213|false|false|false|||segments
Event|Event|Hospital Course|7226,7234|false|false|false|||supports
Finding|Functional Concept|Hospital Course|7238,7246|false|false|false|C0475224|Ischemic|ischemic
Event|Event|Hospital Course|7247,7252|false|false|false|C0441471|Event|event
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7254,7261|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|7254,7261|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|Hospital Course|7263,7267|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7263,7267|false|false|false|C0007430|Catheterization|cath
Event|Event|Hospital Course|7268,7276|false|false|false|||revealed
Anatomy|Body Location or Region|Hospital Course|7279,7285|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7279,7285|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|7286,7293|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|7286,7293|false|false|false|||disease
Finding|Body Substance|Hospital Course|7295,7302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7295,7302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7295,7302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7307,7314|false|false|false|||managed
Drug|Organic Chemical|Hospital Course|7331,7336|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|7331,7336|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|7331,7336|false|false|false|||lasix
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7338,7348|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|7338,7348|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|7338,7348|false|false|false|||lisinopril
Drug|Organic Chemical|Hospital Course|7354,7364|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|7354,7364|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|7354,7364|false|false|false|||metoprolol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7366,7373|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|7366,7373|false|false|false|C1314974|Cardiac attachment|Cardiac
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7366,7381|false|false|false|C0018821|Cardiac Surgery procedures|Cardiac surgery
Event|Event|Hospital Course|7374,7381|false|false|false|||surgery
Finding|Finding|Hospital Course|7374,7381|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|7374,7381|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|7374,7381|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7374,7381|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Hospital Course|7387,7396|false|false|false|||consulted
Finding|Finding|Hospital Course|7401,7409|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|7410,7414|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7410,7414|false|true|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7419,7431|false|false|false|C0026264|Mitral Valve|mitral valve
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7419,7438|false|false|false|C0396849|Mitral valvuloplasty|mitral valve repair
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7426,7431|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Hospital Course|7432,7438|false|false|false|||repair
Finding|Functional Concept|Hospital Course|7432,7438|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Hospital Course|7432,7438|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Hospital Course|7432,7438|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7432,7438|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|Hospital Course|7439,7450|false|false|false|||replacement
Finding|Functional Concept|Hospital Course|7439,7450|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Hospital Course|7439,7450|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7439,7450|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|Hospital Course|7481,7494|false|false|false|||comorbidities
Finding|Finding|Hospital Course|7481,7494|false|false|false|C0009488|Comorbidity|comorbidities
Finding|Finding|Hospital Course|7503,7517|false|false|false|C5787630|Extremely high|extremely high
Event|Event|Hospital Course|7513,7517|false|false|false|||high
Finding|Finding|Hospital Course|7513,7517|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|7513,7517|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|7513,7517|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|Hospital Course|7519,7523|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|7519,7523|false|false|false|C0035647|Risk|risk
Event|Event|Hospital Course|7528,7535|false|false|false|||surgery
Finding|Finding|Hospital Course|7528,7535|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|7528,7535|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|7528,7535|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7528,7535|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Hospital Course|7540,7548|false|false|false|||deferred
Event|Event|Hospital Course|7565,7573|false|false|false|||decision
Finding|Mental Process|Hospital Course|7565,7573|false|false|false|C0679006|Decision|decision
Event|Event|Hospital Course|7587,7600|false|false|false|||revascularize
Finding|Body Substance|Hospital Course|7605,7612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7605,7612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7605,7612|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7618,7621|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Hospital Course|7618,7621|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|Hospital Course|7618,7621|false|false|false|||PCI
Finding|Gene or Genome|Hospital Course|7618,7621|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Hospital Course|7618,7621|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7618,7621|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Event|Hospital Course|7625,7628|false|false|false|||see
Finding|Body Substance|Hospital Course|7636,7643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7636,7643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7636,7643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Food|Hospital Course|7651,7657|false|false|false|C1875723|REGAIN|regain
Event|Event|Hospital Course|7658,7666|false|false|false|||function
Finding|Finding|Hospital Course|7658,7666|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|7658,7666|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|7658,7666|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|7658,7666|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7674,7686|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7681,7686|false|false|false|C1186983|Anatomical valve|valve
Finding|Body Substance|Hospital Course|7688,7695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7688,7695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7688,7695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7696,7704|false|false|false|||received
Drug|Inorganic Chemical|Hospital Course|7713,7718|false|false|false|C0025552|Metals|metal
Event|Event|Hospital Course|7719,7724|false|false|false|||stent
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7732,7735|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|Hospital Course|7732,7735|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|Hospital Course|7732,7735|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7750,7757|false|false|false|C0004704|Balloon Dilatation|balloon
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7750,7769|false|false|false|C0002996;C0002997|Angioplasty, Balloon;Angioplasty, Balloon, Coronary|balloon angioplasty
Event|Event|Hospital Course|7758,7769|false|false|false|||angioplasty
Procedure|Health Care Activity|Hospital Course|7758,7769|false|false|false|C0162577;C1548817|Angioplasty;Angioplasty - Consent Type|angioplasty
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7758,7769|false|false|false|C0162577;C1548817|Angioplasty;Angioplasty - Consent Type|angioplasty
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7787,7793|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|7787,7793|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|Hospital Course|7795,7801|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|Hospital Course|7802,7806|false|false|false|||echo
Procedure|Health Care Activity|Hospital Course|7802,7806|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7802,7806|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|Hospital Course|7807,7813|false|false|false|||showed
Event|Event|Hospital Course|7814,7825|false|false|false|||improvement
Finding|Conceptual Entity|Hospital Course|7814,7825|false|false|false|C2986411|Improvement|improvement
Disorder|Disease or Syndrome|Hospital Course|7834,7854|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Hospital Course|7841,7854|false|false|false|||regurgitation
Finding|Finding|Hospital Course|7841,7854|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|7841,7854|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|7841,7854|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Disorder|Disease or Syndrome|Hospital Course|7860,7866|false|false|false|C4255010||NSTEMI
Event|Event|Hospital Course|7860,7866|false|false|false|||NSTEMI
Finding|Finding|Hospital Course|7860,7866|false|false|false|C3537184||NSTEMI
Disorder|Disease or Syndrome|Hospital Course|7867,7870|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7867,7870|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7867,7870|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7867,7870|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7867,7870|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7867,7870|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7867,7870|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7867,7870|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|7875,7884|false|false|false|||evidenced
Finding|Intellectual Product|Hospital Course|7888,7891|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|7888,7891|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|7892,7899|false|false|false|||changes
Finding|Functional Concept|Hospital Course|7892,7899|false|false|false|C0392747|Changing|changes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7904,7912|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|7904,7912|false|false|false|C0041199|Troponin|troponin
Event|Event|Hospital Course|7904,7912|false|false|false|||troponin
Procedure|Laboratory Procedure|Hospital Course|7904,7912|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|Hospital Course|7913,7917|false|false|false|||leak
Finding|Functional Concept|Hospital Course|7913,7917|false|false|false|C0332234|Leaking|leak
Finding|Body Substance|Hospital Course|7919,7926|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7919,7926|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7919,7926|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7940,7947|false|false|false|||started
Drug|Biologically Active Substance|Hospital Course|7953,7960|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7953,7960|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|7953,7960|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|7961,7965|false|false|false|||drip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7985,7992|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|7985,7992|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Hospital Course|7994,8009|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7994,8009|false|false|false|C0007430|Catheterization|catheterization
Finding|Idea or Concept|Hospital Course|8014,8019|false|false|false|C1552828|Table Frame - above|above
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8021,8028|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|8021,8028|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|Hospital Course|8021,8044|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|Hospital Course|8021,8044|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|Hospital Course|8021,8044|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|Hospital Course|8021,8044|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|Hospital Course|8029,8044|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8029,8044|false|false|false|C0007430|Catheterization|catheterization
Event|Event|Hospital Course|8045,8053|false|false|false|||revealed
Anatomy|Body Location or Region|Hospital Course|8057,8063|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8057,8063|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|8064,8071|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|8064,8071|false|false|false|||disease
Finding|Body Substance|Hospital Course|8073,8080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8073,8080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8073,8080|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8105,8112|false|false|false|||managed
Drug|Organic Chemical|Hospital Course|8119,8126|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|8119,8126|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|8119,8126|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|8128,8134|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|8128,8134|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|8128,8134|false|false|false|||plavix
Drug|Organic Chemical|Hospital Course|8136,8146|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8136,8146|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|8136,8146|false|false|false|||metoprolol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8148,8158|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|8148,8158|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|8148,8158|false|false|false|||lisinopril
Drug|Organic Chemical|Hospital Course|8164,8176|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8164,8176|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|8164,8176|false|false|false|||atorvastatin
Finding|Body Substance|Hospital Course|8186,8193|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8186,8193|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8186,8193|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|8203,8211|false|false|false|C4036058|Too high|too high
Finding|Finding|Hospital Course|8207,8211|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|8207,8211|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|8207,8211|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Hospital Course|8207,8216|false|false|false|C0332167;C4050568;C4319571;C5202937;C5238223|Disease Risk Index High Risk;High Risk Acute Leukemia;High risk;High risk of;International Prognostic Index High Risk Group|high risk
Finding|Intellectual Product|Hospital Course|8207,8216|false|false|false|C0332167;C4050568;C4319571;C5202937;C5238223|Disease Risk Index High Risk;High Risk Acute Leukemia;High risk;High risk of;International Prognostic Index High Risk Group|high risk
Event|Event|Hospital Course|8212,8216|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|8212,8216|false|false|false|C0035647|Risk|risk
Event|Event|Hospital Course|8221,8225|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8221,8225|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Body Substance|Hospital Course|8227,8234|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8227,8234|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8227,8234|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|8235,8243|false|false|false|||returned
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8252,8256|false|false|false|C0007430|Catheterization|cath
Finding|Gene or Genome|Hospital Course|8257,8260|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|Hospital Course|8257,8260|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Drug|Inorganic Chemical|Hospital Course|8276,8281|false|false|false|C0025552|Metals|metal
Event|Event|Hospital Course|8282,8287|false|false|false|||stent
Event|Event|Hospital Course|8292,8296|false|false|false|||POBA
Drug|Organic Chemical|Hospital Course|8316,8322|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|8316,8322|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|8316,8322|false|false|false|||plavix
Finding|Idea or Concept|Hospital Course|8338,8343|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|8338,8343|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Disorder|Disease or Syndrome|Hospital Course|8348,8360|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|8348,8360|false|false|false|||Hypertension
Finding|Body Substance|Hospital Course|8362,8369|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8362,8369|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8362,8369|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8370,8378|false|false|false|||remained
Event|Event|Hospital Course|8379,8391|false|false|false|||normotensive
Event|Event|Hospital Course|8393,8402|false|false|false|||Continued
Drug|Organic Chemical|Hospital Course|8404,8414|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|8404,8414|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|8404,8414|false|false|false|||nifedipine
Finding|Idea or Concept|Hospital Course|8430,8434|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8430,8434|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8430,8434|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8435,8439|false|false|false|||dose
Event|Event|Hospital Course|8441,8450|false|false|false|||Continued
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8454,8464|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|8454,8464|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|8454,8464|false|false|false|||lisinopril
Event|Event|Hospital Course|8480,8487|false|false|false|||started
Drug|Organic Chemical|Hospital Course|8491,8501|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8491,8501|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|8491,8501|false|false|false|||metoprolol
Finding|Idea or Concept|Hospital Course|8505,8510|false|false|false|C1552828|Table Frame - above|above
Anatomy|Body Space or Junction|Hospital Course|8515,8518|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|8515,8518|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|8515,8518|false|false|false|||CHF
Disorder|Disease or Syndrome|Hospital Course|8523,8531|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Hospital Course|8523,8531|false|false|false|||Diabetes
Event|Event|Hospital Course|8533,8542|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|8543,8547|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8543,8547|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8543,8547|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8548,8555|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|8548,8555|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|8548,8555|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|8548,8555|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|8548,8555|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|8548,8555|false|false|false|C0202098|Insulin measurement|insulin
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8548,8562|false|false|false|C0557978|Insulin regime|insulin regime
Event|Event|Hospital Course|8556,8562|false|false|false|||regime
Disorder|Disease or Syndrome|Hospital Course|8569,8572|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Hospital Course|8569,8572|false|false|false|||CKD
Attribute|Clinical Attribute|Hospital Course|8573,8578|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|8573,8581|false|false|false|C0441772|Stage level 4|stage IV
Drug|Biomedical or Dental Material|Hospital Course|8583,8591|false|false|false|C0168634|BaseLine dental cement|Baseline
Finding|Idea or Concept|Hospital Course|8583,8591|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8607,8612|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|8607,8612|false|false|false|C0042075|Urologic Diseases|renal
Event|Event|Hospital Course|8613,8618|false|false|false|||notes
Drug|Biomedical or Dental Material|Hospital Course|8634,8642|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|8634,8642|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|8634,8642|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|8648,8655|false|false|false|||History
Finding|Conceptual Entity|Hospital Course|8648,8655|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|8648,8655|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|8648,8655|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|8648,8658|false|false|false|C0262926|Medical History|History of
Disorder|Disease or Syndrome|Hospital Course|8659,8662|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Hospital Course|8659,8662|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Hospital Course|8659,8662|false|false|false|||CVA
Event|Event|Hospital Course|8664,8673|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|8674,8678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8674,8678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8674,8678|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|8679,8686|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|8679,8686|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|8679,8686|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|8691,8702|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|8691,8702|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|Hospital Course|8691,8702|false|false|false|||clopidogrel
Disorder|Disease or Syndrome|Hospital Course|8708,8712|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Hospital Course|8708,8712|false|false|false|||GERD
Event|Event|Hospital Course|8714,8723|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|8724,8728|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8724,8728|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8724,8728|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|8729,8739|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|8729,8739|false|false|false|C0034665|ranitidine|ranitidine
Event|Event|Hospital Course|8729,8739|false|false|false|||ranitidine
Finding|Idea or Concept|Hospital Course|8742,8754|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|8755,8761|false|false|false|||ISSUES
Event|Event|Hospital Course|8771,8775|false|false|false|||need
Event|Event|Hospital Course|8776,8782|false|false|false|||follow
Finding|Body Substance|Hospital Course|8807,8814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8807,8814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8807,8814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8824,8833|false|false|false|||scheduled
Event|Event|Hospital Course|8837,8843|false|false|false|||follow
Finding|Functional Concept|Hospital Course|8862,8871|false|false|false|C0470187|Availability of|available
Event|Event|Hospital Course|8872,8876|false|false|false|||CMED
Event|Event|Hospital Course|8878,8890|false|false|false|||cardiologist
Event|Event|Hospital Course|8900,8904|false|false|false|||need
Drug|Organic Chemical|Hospital Course|8905,8911|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|8905,8911|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|8905,8911|false|false|false|||plavix
Finding|Idea or Concept|Hospital Course|8929,8934|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|8929,8934|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Idea or Concept|Hospital Course|8936,8939|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8936,8939|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Inorganic Chemical|Hospital Course|8948,8953|false|false|false|C0025552|Metals|metal
Event|Event|Hospital Course|8948,8953|false|false|false|||metal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8955,8970|false|false|false|C2348535|Stenting|stent placement
Event|Event|Hospital Course|8961,8970|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|8961,8970|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8961,8970|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Drug|Organic Chemical|Hospital Course|8980,8992|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8980,8992|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|8993,8997|false|false|false|||dose
Event|Event|Hospital Course|8998,9007|false|false|false|||increased
Event|Event|Hospital Course|9021,9029|false|false|false|||pharmacy
Finding|Intellectual Product|Hospital Course|9021,9029|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Hospital Course|9021,9029|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|Hospital Course|9036,9045|false|false|false|||insurance
Finding|Idea or Concept|Hospital Course|9036,9045|false|false|false|C0021672|Insurance|insurance
Event|Event|Hospital Course|9051,9056|false|false|false|||cover
Finding|Idea or Concept|Hospital Course|9081,9086|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|9081,9086|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Drug|Organic Chemical|Hospital Course|9110,9120|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|9110,9120|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|9121,9125|false|false|false|||dose
Disorder|Disease or Syndrome|Hospital Course|9143,9148|false|false|false|C1410088|Still|still
Event|Event|Hospital Course|9150,9162|false|false|false|||hypertensive
Finding|Finding|Hospital Course|9150,9162|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Event|Event|Hospital Course|9174,9181|false|false|false|||recheck
Finding|Idea or Concept|Hospital Course|9191,9195|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Finding|Hospital Course|9191,9207|false|false|false|C1272171|Next appointment|next appointment
Event|Activity|Hospital Course|9196,9207|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|9196,9207|false|false|false|||appointment
Event|Event|Hospital Course|9211,9219|false|false|false|||evaluate
Disorder|Neoplastic Process|Hospital Course|9229,9238|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|9229,9238|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|9229,9238|false|false|false|C1522484|metastatic qualifier|secondary
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|9242,9245|false|false|false|C0013343|Dyes|dye
Event|Event|Hospital Course|9242,9245|false|false|false|||dye
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9262,9269|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|9262,9269|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|Hospital Course|9262,9285|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|Hospital Course|9262,9285|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|Hospital Course|9262,9285|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|Hospital Course|9262,9285|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|Hospital Course|9270,9285|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9270,9285|false|false|false|C0007430|Catheterization|catheterization
Attribute|Clinical Attribute|Hospital Course|9289,9300|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9289,9300|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9289,9300|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9289,9300|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|9289,9313|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|9304,9313|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|9304,9313|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|9332,9342|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|9332,9342|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|9332,9347|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|9343,9347|false|false|false|||list
Finding|Intellectual Product|Hospital Course|9343,9347|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|9351,9359|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|9364,9372|false|false|false|||complete
Finding|Functional Concept|Hospital Course|9364,9372|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|9364,9372|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9377,9387|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|9377,9387|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|9407,9417|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|9407,9417|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|9407,9417|false|false|false|||NIFEdipine
Drug|Organic Chemical|Hospital Course|9440,9450|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|9440,9450|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|9471,9482|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|Hospital Course|9471,9482|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9502,9509|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|9502,9509|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|9502,9509|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9502,9515|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|9502,9515|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|9502,9515|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9517,9524|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|9517,9524|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|9517,9524|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|9517,9524|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|9517,9524|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|9517,9524|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9517,9528|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|9517,9528|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|9517,9528|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9525,9528|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|9525,9528|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|9525,9528|false|false|false|||NPH
Finding|Functional Concept|Hospital Course|9558,9570|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Element, Ion, or Isotope|Hospital Course|9581,9588|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|9581,9596|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|9581,9596|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9589,9596|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|9589,9596|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|9589,9596|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|9589,9596|false|false|false|||Sulfate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9607,9610|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9607,9610|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9607,9610|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9607,9610|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9607,9610|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9615,9625|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|9615,9625|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|Hospital Course|9645,9658|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9645,9658|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9645,9658|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|9645,9658|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9661,9664|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9661,9664|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|9678,9691|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|9678,9691|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|9678,9694|false|false|false|||Nitroglycerin SL
Finding|Gene or Genome|Hospital Course|9705,9708|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|9709,9714|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9709,9714|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9709,9719|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9709,9719|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9715,9719|false|true|false|C2598155||pain
Event|Event|Hospital Course|9715,9719|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9715,9719|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9715,9719|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|9725,9740|false|false|false|C0012522|diphenhydramine|DiphenhydrAMINE
Drug|Pharmacologic Substance|Hospital Course|9725,9740|false|false|false|C0012522|diphenhydramine|DiphenhydrAMINE
Finding|Gene or Genome|Hospital Course|9753,9756|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|9757,9765|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|9757,9765|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|9757,9765|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|9771,9780|false|false|false|C0718050|sevelamer|sevelamer
Drug|Pharmacologic Substance|Hospital Course|9771,9780|false|false|false|C0718050|sevelamer|sevelamer
Event|Event|Hospital Course|9771,9780|false|false|false|||sevelamer
Drug|Organic Chemical|Hospital Course|9771,9790|false|false|false|C1721288|sevelamer carbonate|sevelamer CARBONATE
Drug|Pharmacologic Substance|Hospital Course|9771,9790|false|false|false|C1721288|sevelamer carbonate|sevelamer CARBONATE
Drug|Element, Ion, or Isotope|Hospital Course|9781,9790|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Drug|Organic Chemical|Hospital Course|9781,9790|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Drug|Pharmacologic Substance|Hospital Course|9781,9790|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Event|Event|Hospital Course|9801,9804|false|false|false|||TID
Event|Event|Hospital Course|9807,9812|false|false|false|||MEALS
Finding|Daily or Recreational Activity|Hospital Course|9807,9812|false|false|false|C1998602|Meal (occasion for eating)|MEALS
Drug|Organic Chemical|Hospital Course|9818,9829|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|9818,9829|false|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|Hospital Course|9854,9860|false|false|false|||taking
Drug|Organic Chemical|Hospital Course|9876,9883|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9876,9883|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9904,9911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9904,9911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9904,9911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|9904,9913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9904,9913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9904,9913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9904,9913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9904,9913|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|9912,9913|false|false|false|||D
Event|Event|Hospital Course|9918,9922|false|false|false|||UNIT
Event|Event|Hospital Course|9936,9945|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9936,9945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9936,9945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9936,9945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9936,9945|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9936,9957|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9946,9957|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9946,9957|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9946,9957|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9946,9957|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9962,9969|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9962,9969|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9989,10000|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|9989,10000|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|10020,10030|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|10020,10030|false|false|false|C0016860|furosemide|Furosemide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10050,10060|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|10050,10060|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|10080,10093|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|10080,10093|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|10080,10093|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|10080,10093|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|10096,10099|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|10096,10099|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|10113,10123|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|10113,10123|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|10144,10153|false|false|false|C0718050|sevelamer|sevelamer
Drug|Pharmacologic Substance|Hospital Course|10144,10153|false|false|false|C0718050|sevelamer|sevelamer
Event|Event|Hospital Course|10144,10153|false|false|false|||sevelamer
Drug|Organic Chemical|Hospital Course|10144,10163|false|false|false|C1721288|sevelamer carbonate|sevelamer CARBONATE
Drug|Pharmacologic Substance|Hospital Course|10144,10163|false|false|false|C1721288|sevelamer carbonate|sevelamer CARBONATE
Drug|Element, Ion, or Isotope|Hospital Course|10154,10163|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Drug|Organic Chemical|Hospital Course|10154,10163|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Drug|Pharmacologic Substance|Hospital Course|10154,10163|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|CARBONATE
Event|Event|Hospital Course|10154,10163|false|false|false|||CARBONATE
Event|Event|Hospital Course|10174,10177|false|false|false|||TID
Event|Event|Hospital Course|10180,10185|false|false|false|||MEALS
Finding|Daily or Recreational Activity|Hospital Course|10180,10185|false|false|false|C1998602|Meal (occasion for eating)|MEALS
Drug|Organic Chemical|Hospital Course|10190,10202|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|10190,10202|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|10223,10235|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|10223,10235|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|10223,10235|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|10244,10250|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10254,10262|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10257,10262|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10257,10262|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|10280,10286|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10287,10294|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10287,10294|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10301,10311|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|10301,10311|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|10301,10321|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|10301,10321|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|10312,10321|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|Hospital Course|10312,10321|false|false|false|||Succinate
Drug|Organic Chemical|Hospital Course|10345,10355|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|10345,10355|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|10345,10365|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|Hospital Course|10345,10365|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|Hospital Course|10356,10365|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|Hospital Course|10356,10365|false|false|false|||succinate
Drug|Biomedical or Dental Material|Hospital Course|10374,10380|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Finding|Hospital Course|10381,10389|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|Hospital Course|10381,10389|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Event|Event|Hospital Course|10390,10397|false|false|false|||release
Finding|Functional Concept|Hospital Course|10390,10397|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|10390,10397|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10390,10397|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Functional Concept|Hospital Course|10408,10416|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10411,10416|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10411,10416|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|10433,10439|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10440,10447|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10440,10447|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10455,10470|false|false|false|C0012522|diphenhydramine|DiphenhydrAMINE
Drug|Pharmacologic Substance|Hospital Course|10455,10470|false|false|false|C0012522|diphenhydramine|DiphenhydrAMINE
Finding|Gene or Genome|Hospital Course|10483,10486|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|10487,10495|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|10487,10495|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|10487,10495|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10501,10508|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|10501,10508|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|10501,10508|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10501,10514|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|10501,10514|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|10501,10514|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10516,10523|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|10516,10523|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|10516,10523|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|10516,10523|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|10516,10523|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|10516,10523|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10516,10527|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|10516,10527|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|10516,10527|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10524,10527|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|10524,10527|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|10524,10527|false|false|false|||NPH
Finding|Functional Concept|Hospital Course|10557,10569|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|Hospital Course|10581,10594|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|10581,10594|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|10581,10594|false|false|false|||Nitroglycerin
Finding|Gene or Genome|Hospital Course|10608,10611|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|10612,10617|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10612,10617|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|10612,10622|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|10612,10622|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|10618,10622|false|true|false|C2598155||pain
Event|Event|Hospital Course|10618,10622|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10618,10622|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10618,10622|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|10628,10635|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|10628,10635|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|10628,10635|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|10628,10637|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|10628,10637|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|10628,10637|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|10628,10637|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|10628,10637|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|10642,10646|false|false|false|||UNIT
Drug|Organic Chemical|Hospital Course|10661,10671|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|10661,10671|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|10661,10671|false|false|false|||NIFEdipine
Event|Event|Hospital Course|10672,10674|false|false|false|||CR
Event|Event|Hospital Course|10694,10703|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10694,10703|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10694,10703|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10694,10703|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10694,10703|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10694,10715|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10694,10715|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10704,10715|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|10704,10715|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|10704,10715|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|10717,10721|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|10717,10721|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|10717,10721|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|10717,10721|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|10727,10734|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|10727,10734|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|10737,10745|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|10737,10745|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|10753,10762|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10753,10762|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10753,10762|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10753,10762|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10753,10762|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10753,10772|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10763,10772|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|10763,10772|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|10763,10772|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10763,10772|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10763,10772|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Principle Diagnosis|10793,10799|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Principle Diagnosis|10793,10799|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Finding|Principle Diagnosis|10793,10820|false|false|false|C5393153|Severe mitral regurgitation|Severe mitral regurgitation
Disorder|Disease or Syndrome|Principle Diagnosis|10800,10820|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Principle Diagnosis|10807,10820|false|false|false|||regurgitation
Finding|Finding|Principle Diagnosis|10807,10820|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Principle Diagnosis|10807,10820|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Principle Diagnosis|10807,10820|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10821,10829|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10821,10836|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Principle Diagnosis|10821,10844|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10830,10836|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Principle Diagnosis|10830,10836|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Principle Diagnosis|10830,10844|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Principle Diagnosis|10837,10844|false|false|false|C0012634|Disease|disease
Event|Event|Principle Diagnosis|10837,10844|false|false|false|||disease
Disorder|Neoplastic Process|Principle Diagnosis|10846,10855|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Event|Event|Principle Diagnosis|10846,10855|false|false|false|||SECONDARY
Finding|Functional Concept|Principle Diagnosis|10846,10855|false|false|false|C1522484|metastatic qualifier|SECONDARY
Attribute|Clinical Attribute|Principle Diagnosis|10846,10865|false|false|false|C4255018||SECONDARY DIAGNOSIS
Finding|Finding|Principle Diagnosis|10846,10865|false|false|false|C0332138|Secondary diagnosis|SECONDARY DIAGNOSIS
Attribute|Clinical Attribute|Principle Diagnosis|10856,10865|false|false|false|C0945731||DIAGNOSIS
Finding|Classification|Principle Diagnosis|10856,10865|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|Principle Diagnosis|10856,10865|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|Principle Diagnosis|10856,10865|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Disorder|Disease or Syndrome|Principle Diagnosis|10867,10879|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Principle Diagnosis|10867,10879|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Principle Diagnosis|10880,10888|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Principle Diagnosis|10880,10888|false|false|false|||Diabetes
Finding|Mental Process|Discharge Condition|10913,10919|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10913,10926|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10913,10926|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10920,10926|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10920,10926|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10928,10933|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|10928,10933|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|10938,10946|false|false|false|||coherent
Finding|Finding|Discharge Condition|10938,10946|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|10948,10953|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|10948,10970|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10948,10970|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|10957,10970|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|10957,10970|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10957,10970|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10972,10977|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10972,10977|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10972,10977|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|10972,10977|false|false|false|||Alert
Finding|Finding|Discharge Condition|10972,10977|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10972,10977|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10972,10977|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|10982,10993|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|10982,10993|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10995,11003|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10995,11003|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10995,11003|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11004,11010|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11004,11010|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11004,11010|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11012,11022|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|11012,11022|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11012,11022|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11012,11022|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11012,11022|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11025,11036|false|false|false|||Independent
Finding|Finding|Discharge Condition|11025,11036|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|11025,11036|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|11065,11069|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|11089,11097|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|11089,11097|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|11089,11097|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|Discharge Instructions|11098,11104|false|false|false|||caring
Event|Event|Discharge Instructions|11133,11139|false|false|false|||recall
Event|Event|Discharge Instructions|11150,11158|false|false|false|||admitted
Event|Event|Discharge Instructions|11163,11172|false|false|false|||shortness
Finding|Body Substance|Discharge Instructions|11177,11183|false|false|false|C0225386|Breath|breath
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11214,11219|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11214,11219|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11214,11219|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11214,11226|false|false|false|C0018826|Heart Valves|heart valves
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11220,11226|false|false|false|C1186983|Anatomical valve|valves
Event|Event|Discharge Instructions|11231,11235|false|false|false|||weak
Finding|Intellectual Product|Discharge Instructions|11231,11235|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|11231,11235|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|Discharge Instructions|11244,11250|false|false|false|||caused
Drug|Substance|Discharge Instructions|11251,11256|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|11251,11256|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|11251,11256|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|11260,11265|false|false|false|||build
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11277,11282|false|false|false|C0024109|Lung|lungs
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11289,11294|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11289,11294|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|11289,11294|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11289,11300|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11295,11300|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Discharge Instructions|11306,11310|false|false|false|||weak
Finding|Intellectual Product|Discharge Instructions|11306,11310|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|11306,11310|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|Discharge Instructions|11331,11339|false|false|false|||blockage
Finding|Finding|Discharge Instructions|11331,11339|false|false|false|C1706968;C1879887;C2237319|Blockage (obstruction - finding);Partial Blockage within Medical Device|blockage
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11355,11360|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11355,11360|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Discharge Instructions|11355,11360|false|false|false|||heart
Finding|Sign or Symptom|Discharge Instructions|11355,11360|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11362,11370|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|Discharge Instructions|11362,11370|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|Discharge Instructions|11362,11370|false|false|false|||arteries
Procedure|Health Care Activity|Discharge Instructions|11362,11370|false|false|false|C0397581|Procedure on artery|arteries
Attribute|Clinical Attribute|Discharge Instructions|11388,11397|false|false|false|C0945766||procedure
Event|Event|Discharge Instructions|11388,11397|false|false|false|||procedure
Event|Occupational Activity|Discharge Instructions|11388,11397|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Discharge Instructions|11388,11397|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11388,11397|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Discharge Instructions|11399,11405|false|false|false|||called
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11406,11413|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Discharge Instructions|11406,11413|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Discharge Instructions|11415,11430|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11415,11430|false|false|false|C0007430|Catheterization|catheterization
Event|Event|Discharge Instructions|11438,11444|false|false|false|||opened
Finding|Finding|Discharge Instructions|11452,11459|false|false|false|C0028778;C0332206|Blocking;Obstruction|blocked
Finding|Functional Concept|Discharge Instructions|11452,11459|false|false|false|C0028778;C0332206|Blocking;Obstruction|blocked
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11460,11468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|Discharge Instructions|11460,11468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|Discharge Instructions|11460,11468|false|false|false|C0397581|Procedure on artery|arteries
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11476,11481|false|false|false|C1186983|Anatomical valve|valve
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11486,11491|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|11486,11491|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Discharge Instructions|11486,11491|false|false|false|||heart
Finding|Sign or Symptom|Discharge Instructions|11486,11491|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Discharge Instructions|11496,11503|false|false|false|||pumping
Finding|Finding|Discharge Instructions|11504,11508|false|false|false|C4281574|Much|much
Event|Event|Discharge Instructions|11552,11559|false|false|false|||feeling
Finding|Finding|Discharge Instructions|11552,11566|false|false|false|C0424578|Psychological Well Being|feeling better
Event|Event|Discharge Instructions|11560,11566|false|false|false|||better
Finding|Idea or Concept|Discharge Instructions|11560,11566|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|11575,11580|false|false|false|||weigh
Finding|Intellectual Product|Discharge Instructions|11590,11595|false|false|false|C1720374|Every - dosing instruction fragment|every
Event|Event|Discharge Instructions|11610,11614|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|11631,11637|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|11631,11637|false|false|false|||weight
Finding|Finding|Discharge Instructions|11631,11637|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|11631,11637|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|11631,11637|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|11638,11642|false|false|false|||goes
Procedure|Laboratory Procedure|Discharge Instructions|11658,11661|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Procedure|Health Care Activity|Discharge Instructions|11680,11688|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11689,11701|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|11689,11701|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|11689,11701|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

