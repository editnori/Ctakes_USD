 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
ORTHOPAEDICS|155,167
<EOL>|167,168
<EOL>|169,170
Codeine|182,189
/|190,191
Augmentin|192,201
/|202,203
Topamax|204,211
<EOL>|211,212
<EOL>|213,214
Attending|214,223
:|223,224
_|225,226
_|226,227
_|227,228
.|228,229
<EOL>|229,230
<EOL>|231,232
left|249,253
knee|254,258
osteoarthritis|259,273
/|273,274
pain|274,278
<EOL>|278,279
<EOL>|280,281
Major|281,286
Surgical|287,295
or|296,298
Invasive|299,307
Procedure|308,317
:|317,318
<EOL>|318,319
_|319,320
_|320,321
_|321,322
:|322,323
left|324,328
total|329,334
knee|335,339
arthroplasty|340,352
<EOL>|352,353
<EOL>|353,354
<EOL>|355,356
_|384,385
_|385,386
_|386,387
year|388,392
old|393,396
female|397,403
w|404,405
/|405,406
left|406,410
knee|411,415
osteoarthritis|416,430
/|430,431
pain|431,435
who|436,439
failed|440,446
<EOL>|447,448
conservative|448,460
measures|461,469
,|469,470
now|471,474
admitted|475,483
for|484,487
left|488,492
total|493,498
knee|499,503
<EOL>|504,505
arthroplasty|505,517
.|517,518
<EOL>|519,520
<EOL>|521,522
Dyslipidemia|544,556
,|556,557
varicose|558,566
veins|567,572
(|573,574
R|574,575
>|575,576
L|576,577
)|577,578
s|579,580
/|580,581
p|581,582
ligation|583,591
,|591,592
COPD|593,597
,|597,598
OSA|599,602
<EOL>|603,604
(|604,605
+|605,606
CPap|606,610
)|610,611
,|611,612
recent|613,619
URI|620,623
(|624,625
received|625,633
course|634,640
of|641,643
Zithromax|644,653
)|653,654
,|654,655
bilateral|656,665
<EOL>|666,667
PEs|667,670
(|671,672
_|672,673
_|673,674
_|674,675
)|675,676
,|676,677
antiphospholipid|678,694
antibody|695,703
syndrome|704,712
(|713,714
on|714,716
lifelong|717,725
<EOL>|726,727
anticoagulation|727,742
)|742,743
,|743,744
T2DM|745,749
(|750,751
last|751,755
A1C|756,759
6.2|760,763
on|764,766
_|767,768
_|768,769
_|769,770
,|770,771
cerebral|772,780
<EOL>|781,782
aneurysm|782,790
(|791,792
followed|792,800
by|801,803
Dr.|804,807
_|808,809
_|809,810
_|810,811
,|811,812
unchanged|813,822
)|822,823
,|823,824
GERD|825,829
,|829,830
<EOL>|831,832
diverticulosis|832,846
,|846,847
h|848,849
/|849,850
o|850,851
colon|852,857
polyps|858,864
,|864,865
depression|866,876
,|876,877
s|878,879
/|879,880
p|880,881
right|882,887
CMC|888,891
<EOL>|892,893
joint|893,898
arthroplasty|899,911
,|911,912
b|913,914
/|914,915
l|915,916
rotator|917,924
cuff|925,929
repair|930,936
,|936,937
excision|938,946
right|947,952
_|953,954
_|954,955
_|955,956
<EOL>|957,958
digit|958,963
mass|964,968
,|968,969
CCY|970,973
w|974,975
/|975,976
stone|976,981
&|982,983
pancreatic|984,994
duct|995,999
exploration|1000,1011
(|1012,1013
_|1013,1014
_|1014,1015
_|1015,1016
)|1016,1017
,|1017,1018
<EOL>|1019,1020
hysterectomy|1020,1032
,|1032,1033
tonsillectomy|1034,1047
<EOL>|1048,1049
<EOL>|1050,1051
:|1065,1066
<EOL>|1066,1067
_|1067,1068
_|1068,1069
_|1069,1070
<EOL>|1070,1071
:|1085,1086
<EOL>|1086,1087
No|1087,1089
family|1090,1096
hx|1097,1099
of|1100,1102
DVT|1103,1106
or|1107,1109
PE|1110,1112
,|1112,1113
two|1114,1117
sisters|1118,1125
have|1126,1130
atrial|1131,1137
fibrillation|1138,1150
.|1150,1151
<EOL>|1152,1153
<EOL>|1154,1155
<EOL>|1155,1156
<EOL>|1157,1158
Well|1173,1177
appearing|1178,1187
in|1188,1190
no|1191,1193
acute|1194,1199
distress|1200,1208
<EOL>|1210,1211
Afebrile|1212,1220
with|1221,1225
stable|1226,1232
vital|1233,1238
signs|1239,1244
<EOL>|1246,1247
Pain|1248,1252
well|1253,1257
-|1257,1258
controlled|1258,1268
<EOL>|1270,1271
Respiratory|1272,1283
:|1283,1284
CTAB|1285,1289
<EOL>|1291,1292
Cardiovascular|1293,1307
:|1307,1308
RRR|1309,1312
<EOL>|1314,1315
Gastrointestinal|1316,1332
:|1332,1333
NT|1334,1336
/|1336,1337
ND|1337,1339
<EOL>|1341,1342
Genitourinary|1343,1356
:|1356,1357
Voiding|1358,1365
independently|1366,1379
<EOL>|1381,1382
Neurologic|1383,1393
:|1393,1394
Intact|1395,1401
with|1402,1406
no|1407,1409
focal|1410,1415
deficits|1416,1424
<EOL>|1426,1427
Psychiatric|1428,1439
:|1439,1440
Pleasant|1441,1449
,|1449,1450
A|1451,1452
&|1452,1453
O|1453,1454
x3|1455,1457
<EOL>|1459,1460
Musculoskeletal|1461,1476
Lower|1477,1482
Extremity|1483,1492
:|1492,1493
<EOL>|1495,1496
*|1497,1498
Aquacel|1499,1506
dressing|1507,1515
with|1516,1520
scant|1521,1526
serosanguinous|1527,1541
drainage|1542,1550
<EOL>|1552,1553
*|1554,1555
Thigh|1556,1561
full|1562,1566
but|1567,1570
soft|1571,1575
<EOL>|1577,1578
*|1579,1580
No|1581,1583
calf|1584,1588
tenderness|1589,1599
<EOL>|1601,1602
*|1603,1604
_|1605,1606
_|1606,1607
_|1607,1608
strength|1609,1617
<EOL>|1619,1620
*|1621,1622
SILT|1623,1627
,|1627,1628
NVI|1629,1632
distally|1633,1641
<EOL>|1643,1644
*|1645,1646
Toes|1647,1651
warm|1652,1656
<EOL>|1657,1658
<EOL>|1659,1660
Pertinent|1660,1669
Results|1670,1677
:|1677,1678
<EOL>|1678,1679
_|1679,1680
_|1680,1681
_|1681,1682
06|1683,1685
:|1685,1686
30AM|1686,1690
BLOOD|1691,1696
WBC|1697,1700
-|1700,1701
6.8|1701,1704
RBC|1705,1708
-|1708,1709
2|1709,1710
.|1710,1711
69|1711,1713
*|1713,1714
Hgb|1715,1718
-|1718,1719
8|1719,1720
.|1720,1721
3|1721,1722
*|1722,1723
Hct|1724,1727
-|1727,1728
25|1728,1730
.|1730,1731
3|1731,1732
*|1732,1733
<EOL>|1734,1735
MCV|1735,1738
-|1738,1739
94|1739,1741
MCH|1742,1745
-|1745,1746
30.9|1746,1750
MCHC|1751,1755
-|1755,1756
32.8|1756,1760
RDW|1761,1764
-|1764,1765
13.0|1765,1769
RDWSD|1770,1775
-|1775,1776
44.0|1776,1780
Plt|1781,1784
_|1785,1786
_|1786,1787
_|1787,1788
<EOL>|1788,1789
_|1789,1790
_|1790,1791
_|1791,1792
06|1793,1795
:|1795,1796
10AM|1796,1800
BLOOD|1801,1806
WBC|1807,1810
-|1810,1811
6.4|1811,1814
RBC|1815,1818
-|1818,1819
2|1819,1820
.|1820,1821
77|1821,1823
*|1823,1824
Hgb|1825,1828
-|1828,1829
8|1829,1830
.|1830,1831
6|1831,1832
*|1832,1833
Hct|1834,1837
-|1837,1838
26|1838,1840
.|1840,1841
0|1841,1842
*|1842,1843
<EOL>|1844,1845
MCV|1845,1848
-|1848,1849
94|1849,1851
MCH|1852,1855
-|1855,1856
31.0|1856,1860
MCHC|1861,1865
-|1865,1866
33.1|1866,1870
RDW|1871,1874
-|1874,1875
13.1|1875,1879
RDWSD|1880,1885
-|1885,1886
44.7|1886,1890
Plt|1891,1894
_|1895,1896
_|1896,1897
_|1897,1898
<EOL>|1898,1899
_|1899,1900
_|1900,1901
_|1901,1902
06|1903,1905
:|1905,1906
22AM|1906,1910
BLOOD|1911,1916
WBC|1917,1920
-|1920,1921
7.6|1921,1924
RBC|1925,1928
-|1928,1929
3|1929,1930
.|1930,1931
31|1931,1933
*|1933,1934
Hgb|1935,1938
-|1938,1939
10|1939,1941
.|1941,1942
2|1942,1943
*|1943,1944
#|1944,1945
Hct|1946,1949
-|1949,1950
30|1950,1952
.|1952,1953
5|1953,1954
*|1954,1955
#|1955,1956
<EOL>|1957,1958
MCV|1958,1961
-|1961,1962
92|1962,1964
MCH|1965,1968
-|1968,1969
30.8|1969,1973
MCHC|1974,1978
-|1978,1979
33.4|1979,1983
RDW|1984,1987
-|1987,1988
12.8|1988,1992
RDWSD|1993,1998
-|1998,1999
42.6|1999,2003
Plt|2004,2007
_|2008,2009
_|2009,2010
_|2010,2011
<EOL>|2011,2012
_|2012,2013
_|2013,2014
_|2014,2015
06|2016,2018
:|2018,2019
30AM|2019,2023
BLOOD|2024,2029
Plt|2030,2033
_|2034,2035
_|2035,2036
_|2036,2037
<EOL>|2037,2038
_|2038,2039
_|2039,2040
_|2040,2041
06|2042,2044
:|2044,2045
30AM|2045,2049
BLOOD|2050,2055
_|2056,2057
_|2057,2058
_|2058,2059
<EOL>|2059,2060
_|2060,2061
_|2061,2062
_|2062,2063
06|2064,2066
:|2066,2067
10AM|2067,2071
BLOOD|2072,2077
Plt|2078,2081
_|2082,2083
_|2083,2084
_|2084,2085
<EOL>|2085,2086
_|2086,2087
_|2087,2088
_|2088,2089
06|2090,2092
:|2092,2093
10AM|2093,2097
BLOOD|2098,2103
_|2104,2105
_|2105,2106
_|2106,2107
<EOL>|2107,2108
_|2108,2109
_|2109,2110
_|2110,2111
06|2112,2114
:|2114,2115
22AM|2115,2119
BLOOD|2120,2125
Plt|2126,2129
_|2130,2131
_|2131,2132
_|2132,2133
<EOL>|2133,2134
_|2134,2135
_|2135,2136
_|2136,2137
06|2138,2140
:|2140,2141
22AM|2141,2145
BLOOD|2146,2151
_|2152,2153
_|2153,2154
_|2154,2155
<EOL>|2155,2156
_|2156,2157
_|2157,2158
_|2158,2159
10|2160,2162
:|2162,2163
55AM|2163,2167
BLOOD|2168,2173
_|2174,2175
_|2175,2176
_|2176,2177
<EOL>|2177,2178
_|2178,2179
_|2179,2180
_|2180,2181
06|2182,2184
:|2184,2185
22AM|2185,2189
BLOOD|2190,2195
Glucose|2196,2203
-|2203,2204
136|2204,2207
*|2207,2208
UreaN|2209,2214
-|2214,2215
8|2215,2216
Creat|2217,2222
-|2222,2223
0.7|2223,2226
Na|2227,2229
-|2229,2230
138|2230,2233
<EOL>|2234,2235
K|2235,2236
-|2236,2237
3.7|2237,2240
Cl|2241,2243
-|2243,2244
96|2244,2246
HCO3|2247,2251
-|2251,2252
27|2252,2254
AnGap|2255,2260
-|2260,2261
15|2261,2263
<EOL>|2263,2264
_|2264,2265
_|2265,2266
_|2266,2267
06|2268,2270
:|2270,2271
22AM|2271,2275
BLOOD|2276,2281
Calcium|2282,2289
-|2289,2290
8.4|2290,2293
Phos|2294,2298
-|2298,2299
3.1|2299,2302
Mg|2303,2305
-|2305,2306
1.7|2306,2309
<EOL>|2309,2310
<EOL>|2311,2312
The|2335,2338
patient|2339,2346
was|2347,2350
admitted|2351,2359
to|2360,2362
the|2363,2366
Orthopaedic|2367,2378
surgery|2379,2386
service|2387,2394
and|2395,2398
<EOL>|2399,2400
was|2400,2403
taken|2404,2409
to|2410,2412
the|2413,2416
operating|2417,2426
room|2427,2431
for|2432,2435
above|2436,2441
described|2442,2451
procedure|2452,2461
.|2461,2462
<EOL>|2463,2464
Please|2464,2470
see|2471,2474
separately|2475,2485
dictated|2486,2494
operative|2495,2504
report|2505,2511
for|2512,2515
details|2516,2523
.|2523,2524
The|2525,2528
<EOL>|2529,2530
surgery|2530,2537
was|2538,2541
uncomplicated|2542,2555
and|2556,2559
the|2560,2563
patient|2564,2571
tolerated|2572,2581
the|2582,2585
<EOL>|2586,2587
procedure|2587,2596
well|2597,2601
.|2601,2602
Patient|2603,2610
received|2611,2619
perioperative|2620,2633
IV|2634,2636
antibiotics|2637,2648
.|2648,2649
<EOL>|2649,2650
<EOL>|2650,2651
Postoperative|2651,2664
course|2665,2671
was|2672,2675
remarkable|2676,2686
for|2687,2690
the|2691,2694
following|2695,2704
:|2704,2705
<EOL>|2705,2706
POD|2706,2709
#|2710,2711
1|2711,2712
,|2712,2713
patient|2714,2721
was|2722,2725
administered|2726,2738
500ml|2739,2744
bolus|2745,2750
of|2751,2753
IV|2754,2756
fluids|2757,2763
for|2764,2767
<EOL>|2768,2769
hypotension|2769,2780
_|2781,2782
_|2782,2783
_|2783,2784
,|2784,2785
which|2786,2791
she|2792,2795
responded|2796,2805
to|2806,2808
appropriately|2809,2822
.|2822,2823
She|2824,2827
<EOL>|2828,2829
reported|2829,2837
nausea|2838,2844
on|2845,2847
oxycodone|2848,2857
and|2858,2861
was|2862,2865
switched|2866,2874
to|2875,2877
dilaudid|2878,2886
with|2887,2891
<EOL>|2892,2893
no|2893,2895
reported|2896,2904
adverse|2905,2912
effects|2913,2920
.|2920,2921
<EOL>|2921,2922
POD|2922,2925
#|2926,2927
2|2927,2928
,|2928,2929
patient|2930,2937
had|2938,2941
INR|2942,2945
of|2946,2948
1.8|2949,2952
and|2953,2956
lovenox|2957,2964
was|2965,2968
discontinued|2969,2981
.|2981,2982
<EOL>|2983,2984
Patient|2984,2991
will|2992,2996
continue|2997,3005
Coumadin|3006,3014
5mg|3015,3018
daily|3019,3024
.|3024,3025
Next|3026,3030
INR|3031,3034
check|3035,3040
day|3041,3044
<EOL>|3045,3046
after|3046,3051
discharge|3052,3061
.|3061,3062
Please|3063,3069
direct|3070,3076
results|3077,3084
and|3085,3088
all|3089,3092
questions|3093,3102
to|3103,3105
PCP|3106,3109
<EOL>|3110,3111
for|3111,3114
INR|3115,3118
monitoring|3119,3129
/|3129,3130
Coumadin|3130,3138
dosing|3139,3145
.|3145,3146
<EOL>|3146,3147
POD|3147,3150
#|3151,3152
3|3152,3153
,|3153,3154
INR|3155,3158
2.0|3159,3162
and|3163,3166
patient|3167,3174
will|3175,3179
be|3180,3182
due|3183,3186
for|3187,3190
5mg|3191,3194
Coumadin|3195,3203
upon|3204,3208
<EOL>|3209,3210
arrival|3210,3217
to|3218,3220
rehab|3221,3226
facility|3227,3235
.|3235,3236
<EOL>|3236,3237
<EOL>|3237,3238
Otherwise|3238,3247
,|3247,3248
pain|3249,3253
was|3254,3257
controlled|3258,3268
with|3269,3273
a|3274,3275
combination|3276,3287
of|3288,3290
IV|3291,3293
and|3294,3297
oral|3298,3302
<EOL>|3303,3304
pain|3304,3308
medications|3309,3320
.|3320,3321
The|3323,3326
patient|3327,3334
received|3335,3343
Coumadin|3344,3352
starting|3353,3361
on|3362,3364
<EOL>|3365,3366
POD|3366,3369
#|3369,3370
0|3370,3371
with|3372,3376
a|3377,3378
Lovenox|3379,3386
bridge|3387,3393
starting|3394,3402
on|3403,3405
POD|3406,3409
#|3409,3410
1|3410,3411
.|3411,3412
Lovenox|3414,3421
to|3422,3424
be|3425,3427
<EOL>|3428,3429
continued|3429,3438
until|3439,3444
INR|3445,3448
>|3449,3450
1.5|3451,3454
and|3455,3458
discontinued|3459,3471
on|3472,3474
POD|3475,3478
#|3479,3480
2|3480,3481
with|3482,3486
INR|3487,3490
<EOL>|3491,3492
1.8|3492,3495
.|3495,3496
Coumadin|3497,3505
was|3506,3509
dosed|3510,3515
daily|3516,3521
based|3522,3527
on|3528,3530
her|3531,3534
INR|3535,3538
levels|3539,3545
.|3545,3546
The|3548,3551
<EOL>|3552,3553
surgical|3553,3561
dressing|3562,3570
will|3571,3575
remain|3576,3582
on|3583,3585
until|3586,3591
POD|3592,3595
#|3595,3596
7|3596,3597
after|3598,3603
surgery|3604,3611
.|3611,3612
The|3613,3616
<EOL>|3617,3618
patient|3618,3625
was|3626,3629
seen|3630,3634
daily|3635,3640
by|3641,3643
physical|3644,3652
therapy|3653,3660
.|3660,3661
Labs|3662,3666
were|3667,3671
checked|3672,3679
<EOL>|3680,3681
throughout|3681,3691
the|3692,3695
hospital|3696,3704
course|3705,3711
and|3712,3715
repleted|3716,3724
accordingly|3725,3736
.|3736,3737
At|3738,3740
the|3741,3744
<EOL>|3745,3746
time|3746,3750
of|3751,3753
discharge|3754,3763
the|3764,3767
patient|3768,3775
was|3776,3779
tolerating|3780,3790
a|3791,3792
regular|3793,3800
diet|3801,3805
and|3806,3809
<EOL>|3810,3811
feeling|3811,3818
well|3819,3823
.|3823,3824
The|3826,3829
patient|3830,3837
was|3838,3841
afebrile|3842,3850
with|3851,3855
stable|3856,3862
vital|3863,3868
signs|3869,3874
.|3874,3875
<EOL>|3876,3877
The|3878,3881
patient|3882,3889
's|3889,3891
hematocrit|3892,3902
was|3903,3906
acceptable|3907,3917
and|3918,3921
pain|3922,3926
was|3927,3930
adequately|3931,3941
<EOL>|3942,3943
controlled|3943,3953
on|3954,3956
an|3957,3959
oral|3960,3964
regimen|3965,3972
.|3972,3973
The|3974,3977
operative|3978,3987
extremity|3988,3997
was|3998,4001
<EOL>|4002,4003
neurovascularly|4003,4018
intact|4019,4025
and|4026,4029
the|4030,4033
dressing|4034,4042
was|4043,4046
intact|4047,4053
.|4053,4054
<EOL>|4054,4055
<EOL>|4055,4056
The|4056,4059
patient|4060,4067
's|4067,4069
weight|4070,4076
-|4076,4077
bearing|4077,4084
status|4085,4091
is|4092,4094
weight|4095,4101
bearing|4102,4109
as|4110,4112
<EOL>|4113,4114
tolerated|4114,4123
on|4124,4126
the|4127,4130
operative|4131,4140
extremity|4141,4150
.|4150,4151
Please|4152,4158
use|4159,4162
walker|4163,4169
or|4170,4172
2|4173,4174
<EOL>|4175,4176
crutches|4176,4184
,|4184,4185
wean|4186,4190
as|4191,4193
able|4194,4198
.|4198,4199
<EOL>|4199,4200
<EOL>|4200,4201
Ms.|4201,4204
_|4205,4206
_|4206,4207
_|4207,4208
is|4209,4211
discharged|4212,4222
to|4223,4225
rehab|4226,4231
in|4232,4234
stable|4235,4241
condition|4242,4251
.|4251,4252
<EOL>|4252,4253
<EOL>|4253,4254
*|4254,4255
*|4255,4256
Patient|4256,4263
will|4264,4268
be|4269,4271
in|4272,4274
rehab|4275,4280
facility|4281,4289
for|4290,4293
less|4294,4298
than|4299,4303
30|4304,4306
days|4307,4311
*|4311,4312
*|4312,4313
<EOL>|4313,4314
<EOL>|4315,4316
Medications|4316,4327
on|4328,4330
Admission|4331,4340
:|4340,4341
<EOL>|4341,4342
1.|4342,4344
Albuterol|4345,4354
0.083|4355,4360
%|4360,4361
Neb|4362,4365
Soln|4366,4370
2|4371,4372
NEB|4373,4376
IH|4377,4379
Q4H|4380,4383
:|4383,4384
PRN|4384,4387
wheezing|4388,4396
,|4396,4397
cough|4398,4403
<EOL>|4404,4405
2.|4405,4407
Atorvastatin|4408,4420
40|4421,4423
mg|4424,4426
PO|4427,4429
QPM|4430,4433
<EOL>|4434,4435
3.|4435,4437
econazole|4438,4447
1|4448,4449
%|4450,4451
topical|4452,4459
BID|4460,4463
<EOL>|4464,4465
4.|4465,4467
Enoxaparin|4468,4478
Sodium|4479,4485
110|4486,4489
mg|4490,4492
SC|4493,4495
Q12H|4496,4500
<EOL>|4501,4502
Start|4502,4507
:|4507,4508
Today|4509,4514
-|4515,4516
_|4517,4518
_|4518,4519
_|4519,4520
,|4520,4521
First|4522,4527
Dose|4528,4532
:|4532,4533
Next|4534,4538
Routine|4539,4546
Administration|4547,4561
<EOL>|4562,4563
Time|4563,4567
<EOL>|4568,4569
5.|4569,4571
Furosemide|4572,4582
_|4583,4584
_|4584,4585
_|4585,4586
mg|4587,4589
PO|4590,4592
DAILY|4593,4598
:|4598,4599
PRN|4599,4602
leg|4603,4606
swelling|4607,4615
<EOL>|4616,4617
6.|4617,4619
MetFORMIN|4620,4629
(|4630,4631
Glucophage|4631,4641
)|4641,4642
500|4643,4646
mg|4647,4649
PO|4650,4652
QPM|4653,4656
<EOL>|4657,4658
7.|4658,4660
Omeprazole|4661,4671
20|4672,4674
mg|4675,4677
PO|4678,4680
BID|4681,4684
<EOL>|4685,4686
8.|4686,4688
Sertraline|4689,4699
100|4700,4703
mg|4704,4706
PO|4707,4709
DAILY|4710,4715
<EOL>|4716,4717
9.|4717,4719
TraZODone|4720,4729
50|4730,4732
mg|4733,4735
PO|4736,4738
QHS|4739,4742
:|4742,4743
PRN|4743,4746
insomnia|4747,4755
<EOL>|4756,4757
10.|4757,4760
Triamcinolone|4761,4774
Acetonide|4775,4784
0.1|4785,4788
%|4788,4789
Ointment|4790,4798
1|4799,4800
Appl|4801,4805
TP|4806,4808
BID|4809,4812
:|4812,4813
PRN|4813,4816
<EOL>|4817,4818
rash|4818,4822
/|4822,4823
itching|4823,4830
<EOL>|4831,4832
11|4832,4834
.|4834,4835
Warfarin|4836,4844
_|4845,4846
_|4846,4847
_|4847,4848
mg|4849,4851
PO|4852,4854
DAILY16|4855,4862
<EOL>|4863,4864
12.|4864,4867
Aspirin|4868,4875
81|4876,4878
mg|4879,4881
PO|4882,4884
DAILY|4885,4890
<EOL>|4891,4892
13|4892,4894
.|4894,4895
Vitamin|4896,4903
D|4904,4905
_|4906,4907
_|4907,4908
_|4908,4909
UNIT|4910,4914
PO|4915,4917
DAILY|4918,4923
<EOL>|4924,4925
<EOL>|4925,4926
<EOL>|4927,4928
Discharge|4928,4937
Medications|4938,4949
:|4949,4950
<EOL>|4950,4951
1.|4951,4953
Docusate|4955,4963
Sodium|4964,4970
100|4971,4974
mg|4975,4977
PO|4978,4980
BID|4981,4984
<EOL>|4985,4986
2.|4986,4988
Gabapentin|4990,5000
100|5001,5004
mg|5005,5007
PO|5008,5010
TID|5011,5014
<EOL>|5015,5016
3.|5016,5018
HYDROmorphone|5020,5033
(|5034,5035
Dilaudid|5035,5043
)|5043,5044
_|5045,5046
_|5046,5047
_|5047,5048
mg|5049,5051
PO|5052,5054
Q4H|5055,5058
:|5058,5059
PRN|5059,5062
Pain|5063,5067
-|5068,5069
Moderate|5070,5078
<EOL>|5079,5080
do|5080,5082
NOT|5083,5086
drink|5087,5092
alcohol|5093,5100
or|5101,5103
drive|5104,5109
while|5110,5115
taking|5116,5122
med|5123,5126
<EOL>|5127,5128
4.|5128,5130
Senna|5132,5137
8.6|5138,5141
mg|5142,5144
PO|5145,5147
BID|5148,5151
<EOL>|5152,5153
5.|5153,5155
Acetaminophen|5157,5170
1000|5171,5175
mg|5176,5178
PO|5179,5181
Q8H|5182,5185
<EOL>|5186,5187
6.|5187,5189
Warfarin|5191,5199
5|5200,5201
mg|5202,5204
PO|5205,5207
TO|5208,5210
BE|5211,5213
DOSED|5214,5219
DAILY|5220,5225
PER|5226,5229
PCP|5230,5233
<EOL>|5234,5235
DOSED|5235,5240
DAILY|5241,5246
PER|5247,5250
PCP|5251,5254
,|5254,5255
GOAL|5256,5260
INR|5261,5264
1.8|5265,5268
-|5268,5269
2.2|5269,5272
<EOL>|5273,5274
7.|5274,5276
Albuterol|5278,5287
Inhaler|5288,5295
_|5296,5297
_|5297,5298
_|5298,5299
PUFF|5300,5304
IH|5305,5307
Q6H|5308,5311
:|5311,5312
PRN|5312,5315
shortness|5316,5325
of|5326,5328
breath|5329,5335
<EOL>|5337,5338
8.|5338,5340
Aspirin|5342,5349
81|5350,5352
mg|5353,5355
PO|5356,5358
DAILY|5359,5364
<EOL>|5366,5367
9.|5367,5369
Atorvastatin|5371,5383
40|5384,5386
mg|5387,5389
PO|5390,5392
QPM|5393,5396
<EOL>|5398,5399
10.|5399,5402
econazole|5404,5413
1|5414,5415
%|5416,5417
topical|5418,5425
BID|5426,5429
<EOL>|5431,5432
11.|5432,5435
Furosemide|5437,5447
_|5448,5449
_|5449,5450
_|5450,5451
mg|5452,5454
PO|5455,5457
DAILY|5458,5463
:|5463,5464
PRN|5464,5467
leg|5468,5471
swelling|5472,5480
<EOL>|5482,5483
12.|5483,5486
MetFORMIN|5488,5497
XR|5498,5500
(|5501,5502
Glucophage|5502,5512
XR|5513,5515
)|5515,5516
500|5517,5520
mg|5521,5523
PO|5524,5526
DAILY|5527,5532
<EOL>|5534,5535
13.|5535,5538
Omeprazole|5540,5550
20|5551,5553
mg|5554,5556
PO|5557,5559
BID|5560,5563
<EOL>|5565,5566
14.|5566,5569
Sertraline|5571,5581
100|5582,5585
mg|5586,5588
PO|5589,5591
DAILY|5592,5597
<EOL>|5599,5600
15.|5600,5603
TraZODone|5605,5614
50|5615,5617
mg|5618,5620
PO|5621,5623
QHS|5624,5627
:|5627,5628
PRN|5628,5631
insomnia|5632,5640
<EOL>|5642,5643
16|5643,5645
.|5645,5646
Triamcinolone|5648,5661
Acetonide|5662,5671
0.1|5672,5675
%|5675,5676
Ointment|5677,5685
1|5686,5687
Appl|5688,5692
TP|5693,5695
BID|5696,5699
:|5699,5700
PRN|5700,5703
<EOL>|5704,5705
rash|5705,5709
/|5709,5710
itching|5710,5717
<EOL>|5719,5720
17.|5720,5723
Vitamin|5725,5732
D|5733,5734
_|5735,5736
_|5736,5737
_|5737,5738
UNIT|5739,5743
PO|5744,5746
DAILY|5747,5752
<EOL>|5754,5755
<EOL>|5755,5756
<EOL>|5757,5758
Discharge|5758,5767
Disposition|5768,5779
:|5779,5780
<EOL>|5780,5781
Extended|5781,5789
Care|5790,5794
<EOL>|5794,5795
<EOL>|5796,5797
Facility|5797,5805
:|5805,5806
<EOL>|5806,5807
_|5807,5808
_|5808,5809
_|5809,5810
<EOL>|5810,5811
<EOL>|5812,5813
Discharge|5813,5822
Diagnosis|5823,5832
:|5832,5833
<EOL>|5833,5834
left|5834,5838
knee|5839,5843
osteoarthritis|5844,5858
/|5858,5859
pain|5859,5863
<EOL>|5864,5865
<EOL>|5865,5866
<EOL>|5867,5868
Mental|5889,5895
Status|5896,5902
:|5902,5903
Clear|5904,5909
and|5910,5913
coherent|5914,5922
.|5922,5923
<EOL>|5923,5924
Level|5924,5929
of|5930,5932
Consciousness|5933,5946
:|5946,5947
Alert|5948,5953
and|5954,5957
interactive|5958,5969
.|5969,5970
<EOL>|5970,5971
Activity|5971,5979
Status|5980,5986
:|5986,5987
Ambulatory|5988,5998
-|5999,6000
requires|6001,6009
assistance|6010,6020
or|6021,6023
aid|6024,6027
(|6028,6029
walker|6029,6035
<EOL>|6036,6037
or|6037,6039
cane|6040,6044
)|6044,6045
.|6045,6046
<EOL>|6046,6047
<EOL>|6047,6048
<EOL>|6049,6050
1|6074,6075
.|6075,6076
Please|6077,6083
return|6084,6090
to|6091,6093
the|6094,6097
emergency|6098,6107
department|6108,6118
or|6119,6121
notify|6122,6128
your|6129,6133
<EOL>|6134,6135
physician|6135,6144
if|6145,6147
you|6148,6151
experience|6152,6162
any|6163,6166
of|6167,6169
the|6170,6173
following|6174,6183
:|6183,6184
severe|6185,6191
pain|6192,6196
<EOL>|6197,6198
not|6198,6201
relieved|6202,6210
by|6211,6213
medication|6214,6224
,|6224,6225
increased|6226,6235
swelling|6236,6244
,|6244,6245
decreased|6246,6255
<EOL>|6256,6257
sensation|6257,6266
,|6266,6267
difficulty|6268,6278
with|6279,6283
movement|6284,6292
,|6292,6293
fevers|6294,6300
greater|6301,6308
than|6309,6313
101.5|6314,6319
,|6319,6320
<EOL>|6321,6322
shaking|6322,6329
chills|6330,6336
,|6336,6337
increasing|6338,6348
redness|6349,6356
or|6357,6359
drainage|6360,6368
from|6369,6373
the|6374,6377
incision|6378,6386
<EOL>|6387,6388
site|6388,6392
,|6392,6393
chest|6394,6399
pain|6400,6404
,|6404,6405
shortness|6406,6415
of|6416,6418
breath|6419,6425
or|6426,6428
any|6429,6432
other|6433,6438
concerns|6439,6447
.|6447,6448
<EOL>|6448,6449
<EOL>|6451,6452
2.|6452,6454
Please|6455,6461
follow|6462,6468
up|6469,6471
with|6472,6476
your|6477,6481
primary|6482,6489
physician|6490,6499
regarding|6500,6509
this|6510,6514
<EOL>|6515,6516
admission|6516,6525
and|6526,6529
any|6530,6533
new|6534,6537
medications|6538,6549
and|6550,6553
refills|6554,6561
.|6561,6562
<EOL>|6563,6564
<EOL>|6566,6567
3.|6567,6569
Resume|6570,6576
your|6577,6581
home|6582,6586
medications|6587,6598
unless|6599,6605
otherwise|6606,6615
instructed|6616,6626
.|6626,6627
<EOL>|6627,6628
<EOL>|6630,6631
4|6631,6632
.|6632,6633
You|6634,6637
have|6638,6642
been|6643,6647
given|6648,6653
medications|6654,6665
for|6666,6669
pain|6670,6674
control|6675,6682
.|6682,6683
Please|6684,6690
do|6691,6693
<EOL>|6694,6695
not|6695,6698
drive|6699,6704
,|6704,6705
operate|6706,6713
heavy|6714,6719
machinery|6720,6729
,|6729,6730
or|6731,6733
drink|6734,6739
alcohol|6740,6747
while|6748,6753
<EOL>|6754,6755
taking|6755,6761
these|6762,6767
medications|6768,6779
.|6779,6780
As|6781,6783
your|6784,6788
pain|6789,6793
decreases|6794,6803
,|6803,6804
take|6805,6809
fewer|6810,6815
<EOL>|6816,6817
tablets|6817,6824
and|6825,6828
increase|6829,6837
the|6838,6841
time|6842,6846
between|6847,6854
doses|6855,6860
.|6860,6861
This|6862,6866
medication|6867,6877
can|6878,6881
<EOL>|6882,6883
cause|6883,6888
constipation|6889,6901
,|6901,6902
so|6903,6905
you|6906,6909
should|6910,6916
drink|6917,6922
plenty|6923,6929
of|6930,6932
water|6933,6938
daily|6939,6944
<EOL>|6945,6946
and|6946,6949
take|6950,6954
a|6955,6956
stool|6957,6962
softener|6963,6971
(|6972,6973
such|6973,6977
as|6978,6980
Colace|6981,6987
)|6987,6988
as|6989,6991
needed|6992,6998
to|6999,7001
prevent|7002,7009
<EOL>|7010,7011
this|7011,7015
side|7016,7020
effect|7021,7027
.|7027,7028
Call|7030,7034
your|7035,7039
surgeons|7040,7048
office|7049,7055
3|7056,7057
days|7058,7062
before|7063,7069
you|7070,7073
<EOL>|7074,7075
are|7075,7078
out|7079,7082
of|7083,7085
medication|7086,7096
so|7097,7099
that|7100,7104
it|7105,7107
can|7108,7111
be|7112,7114
refilled|7115,7123
.|7123,7124
These|7126,7131
<EOL>|7132,7133
medications|7133,7144
can|7145,7148
not|7148,7151
be|7152,7154
called|7155,7161
into|7162,7166
your|7167,7171
pharmacy|7172,7180
and|7181,7184
must|7185,7189
be|7190,7192
<EOL>|7193,7194
picked|7194,7200
up|7201,7203
in|7204,7206
the|7207,7210
clinic|7211,7217
or|7218,7220
mailed|7221,7227
to|7228,7230
your|7231,7235
house|7236,7241
.|7241,7242
Please|7244,7250
allow|7251,7256
<EOL>|7257,7258
an|7258,7260
extra|7261,7266
2|7267,7268
days|7269,7273
if|7274,7276
you|7277,7280
would|7281,7286
like|7287,7291
your|7292,7296
medication|7297,7307
mailed|7308,7314
to|7315,7317
your|7318,7322
<EOL>|7323,7324
home|7324,7328
.|7328,7329
<EOL>|7329,7330
<EOL>|7332,7333
5|7333,7334
.|7334,7335
You|7336,7339
may|7340,7343
not|7344,7347
drive|7348,7353
a|7354,7355
car|7356,7359
until|7360,7365
cleared|7366,7373
to|7374,7376
do|7377,7379
so|7380,7382
by|7383,7385
your|7386,7390
<EOL>|7391,7392
surgeon|7392,7399
.|7399,7400
<EOL>|7400,7401
<EOL>|7403,7404
6.|7404,7406
Please|7407,7413
call|7414,7418
your|7419,7423
surgeon|7424,7431
's|7431,7433
office|7434,7440
to|7441,7443
schedule|7444,7452
or|7453,7455
confirm|7456,7463
your|7464,7468
<EOL>|7469,7470
follow|7470,7476
-|7476,7477
up|7477,7479
appointment|7480,7491
.|7491,7492
<EOL>|7492,7493
<EOL>|7495,7496
7.|7496,7498
SWELLING|7499,7507
:|7507,7508
Ice|7509,7512
the|7513,7516
operative|7517,7526
joint|7527,7532
20|7533,7535
minutes|7536,7543
at|7544,7546
a|7547,7548
time|7549,7553
,|7553,7554
<EOL>|7555,7556
especially|7556,7566
after|7567,7572
activity|7573,7581
or|7582,7584
physical|7585,7593
therapy|7594,7601
.|7601,7602
Do|7603,7605
not|7606,7609
place|7610,7615
ice|7616,7619
<EOL>|7620,7621
directly|7621,7629
on|7630,7632
the|7633,7636
skin|7637,7641
.|7641,7642
You|7643,7646
may|7647,7650
wrap|7651,7655
the|7656,7659
knee|7660,7664
with|7665,7669
an|7670,7672
ace|7673,7676
bandage|7677,7684
<EOL>|7685,7686
for|7686,7689
added|7690,7695
compression|7696,7707
.|7707,7708
Please|7709,7715
DO|7716,7718
NOT|7719,7722
take|7723,7727
any|7728,7731
non-steroidal|7732,7745
<EOL>|7746,7747
anti-inflammatory|7747,7764
medications|7765,7776
(|7777,7778
NSAIDs|7778,7784
such|7785,7789
as|7790,7792
Celebrex|7793,7801
,|7801,7802
<EOL>|7803,7804
ibuprofen|7804,7813
,|7813,7814
Advil|7815,7820
,|7820,7821
Aleve|7822,7827
,|7827,7828
Motrin|7829,7835
,|7835,7836
naproxen|7837,7845
etc|7846,7849
)|7849,7850
until|7851,7856
cleared|7857,7864
by|7865,7867
<EOL>|7868,7869
your|7869,7873
physician|7874,7883
.|7883,7884
<EOL>|7884,7885
<EOL>|7887,7888
8.|7888,7890
ANTICOAGULATION|7891,7906
:|7906,7907
Lovenox|7908,7915
discontinued|7916,7928
on|7929,7931
_|7932,7933
_|7933,7934
_|7934,7935
due|7936,7939
to|7940,7942
INR|7943,7946
<EOL>|7947,7948
1.8|7948,7951
.|7951,7952
INR|7953,7956
goal|7957,7961
is|7962,7964
1.8|7965,7968
-|7968,7969
2.2|7969,7972
.|7972,7973
Please|7974,7980
continue|7981,7989
Coumadin|7990,7998
5mg|7999,8002
daily|8003,8008
.|8008,8009
<EOL>|8010,8011
INR|8011,8014
to|8015,8017
be|8018,8020
checked|8021,8028
day|8029,8032
after|8033,8038
discharge|8039,8048
.|8048,8049
Please|8050,8056
direct|8057,8063
all|8064,8067
INR|8068,8071
<EOL>|8072,8073
results|8073,8080
to|8081,8083
patient|8084,8091
's|8091,8093
PCP|8094,8097
.|8097,8098
You|8099,8102
may|8103,8106
continue|8107,8115
your|8116,8120
dose|8121,8125
of|8126,8128
Aspirin|8129,8136
<EOL>|8137,8138
81mg|8138,8142
daily|8143,8148
.|8148,8149
<EOL>|8149,8150
<EOL>|8152,8153
9.|8153,8155
WOUND|8156,8161
CARE|8162,8166
:|8166,8167
Please|8168,8174
remove|8175,8181
Aquacel|8182,8189
dressing|8190,8198
on|8199,8201
POD|8202,8205
#|8205,8206
7|8206,8207
after|8208,8213
<EOL>|8214,8215
surgery|8215,8222
.|8222,8223
It|8224,8226
is|8227,8229
okay|8230,8234
to|8235,8237
shower|8238,8244
after|8245,8250
surgery|8251,8258
after|8259,8264
5|8265,8266
days|8267,8271
but|8272,8275
no|8276,8278
<EOL>|8279,8280
tub|8280,8283
baths|8284,8289
,|8289,8290
swimming|8291,8299
,|8299,8300
or|8301,8303
submerging|8304,8314
your|8315,8319
incision|8320,8328
until|8329,8334
after|8335,8340
<EOL>|8341,8342
your|8342,8346
four|8347,8351
(|8352,8353
4|8353,8354
)|8354,8355
week|8356,8360
checkup|8361,8368
.|8368,8369
Please|8370,8376
place|8377,8382
a|8383,8384
dry|8385,8388
sterile|8389,8396
dressing|8397,8405
<EOL>|8406,8407
on|8407,8409
the|8410,8413
wound|8414,8419
after|8420,8425
aqaucel|8426,8433
is|8434,8436
removed|8437,8444
each|8445,8449
day|8450,8453
if|8454,8456
there|8457,8462
is|8463,8465
<EOL>|8466,8467
drainage|8467,8475
,|8475,8476
otherwise|8477,8486
leave|8487,8492
it|8493,8495
open|8496,8500
to|8501,8503
air|8504,8507
.|8507,8508
Check|8509,8514
wound|8515,8520
regularly|8521,8530
<EOL>|8531,8532
for|8532,8535
signs|8536,8541
of|8542,8544
infection|8545,8554
such|8555,8559
as|8560,8562
redness|8563,8570
or|8571,8573
thick|8574,8579
yellow|8580,8586
drainage|8587,8595
.|8595,8596
<EOL>|8597,8598
<EOL>|8599,8600
<EOL>|8600,8601
10.|8601,8604
_|8605,8606
_|8606,8607
_|8607,8608
(|8609,8610
once|8610,8614
at|8615,8617
home|8618,8622
)|8622,8623
:|8623,8624
Home|8625,8629
_|8630,8631
_|8631,8632
_|8632,8633
,|8633,8634
dressing|8635,8643
changes|8644,8651
as|8652,8654
<EOL>|8655,8656
instructed|8656,8666
,|8666,8667
and|8668,8671
wound|8672,8677
checks|8678,8684
.|8684,8685
<EOL>|8685,8686
<EOL>|8688,8689
11|8689,8691
.|8691,8692
ACTIVITY|8693,8701
:|8701,8702
Weight|8703,8709
bearing|8710,8717
as|8718,8720
tolerated|8721,8730
on|8731,8733
the|8734,8737
operative|8738,8747
<EOL>|8748,8749
extremity|8749,8758
.|8758,8759
Two|8760,8763
crutches|8764,8772
or|8773,8775
walker|8776,8782
.|8782,8783
Wean|8785,8789
assistive|8790,8799
device|8800,8806
as|8807,8809
<EOL>|8810,8811
able|8811,8815
.|8815,8816
Mobilize|8817,8825
.|8825,8826
ROM|8828,8831
as|8832,8834
tolerated|8835,8844
.|8844,8845
No|8846,8848
strenuous|8849,8858
exercise|8859,8867
or|8868,8870
<EOL>|8871,8872
heavy|8872,8877
lifting|8878,8885
until|8886,8891
follow|8892,8898
up|8899,8901
appointment|8902,8913
.|8913,8914
<EOL>|8915,8916
<EOL>|8916,8917
Physical|8917,8925
Therapy|8926,8933
:|8933,8934
<EOL>|8934,8935
WBAT|8935,8939
LLE|8940,8943
<EOL>|8943,8944
No|8944,8946
range|8947,8952
of|8953,8955
motion|8956,8962
restrictions|8963,8975
<EOL>|8975,8976
Wean|8976,8980
assistive|8981,8990
devices|8991,8998
as|8999,9001
able|9002,9006
<EOL>|9006,9007
Mobilize|9007,9015
frequently|9016,9026
<EOL>|9026,9027
Treatments|9027,9037
Frequency|9038,9047
:|9047,9048
<EOL>|9048,9049
remove|9049,9055
aquacel|9056,9063
POD|9064,9067
#|9067,9068
7|9068,9069
after|9070,9075
surgery|9076,9083
<EOL>|9083,9084
apply|9084,9089
dry|9090,9093
sterile|9094,9101
dressing|9102,9110
daily|9111,9116
if|9117,9119
needed|9120,9126
after|9127,9132
aquacel|9133,9140
<EOL>|9141,9142
dressing|9142,9150
is|9151,9153
removed|9154,9161
<EOL>|9161,9162
wound|9162,9167
checks|9168,9174
daily|9175,9180
after|9181,9186
aquacel|9187,9194
removed|9195,9202
<EOL>|9202,9203
<EOL>|9203,9204
<EOL>|9205,9206
Followup|9206,9214
Instructions|9215,9227
:|9227,9228
<EOL>|9228,9229
_|9229,9230
_|9230,9231
_|9231,9232
<EOL>|9232,9233

