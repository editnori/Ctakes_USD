 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
M|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
Corgard|176,183
/|184,185
Vasotec|186,193
<EOL>|193,194
<EOL>|195,196
Attending|196,205
:|205,206
_|207,208
_|208,209
_|209,210
.|210,211
<EOL>|211,212
<EOL>|213,214
Chief|214,219
Complaint|220,229
:|229,230
<EOL>|230,231
Dyspnea|231,238
on|239,241
Exertion|242,250
<EOL>|250,251
<EOL>|252,253
Major|253,258
Surgical|259,267
or|268,270
Invasive|271,279
Procedure|280,289
:|289,290
<EOL>|290,291
None|291,295
<EOL>|295,296
<EOL>|296,297
<EOL>|298,299
History|299,306
of|307,309
Present|310,317
Illness|318,325
:|325,326
<EOL>|326,327
=|328,329
=|329,330
=|330,331
=|331,332
=|332,333
=|333,334
=|334,335
=|335,336
=|336,337
=|337,338
=|338,339
=|339,340
=|340,341
=|341,342
=|342,343
=|343,344
=|344,345
=|345,346
=|346,347
=|347,348
=|348,349
=|349,350
=|350,351
=|351,352
=|352,353
=|353,354
=|354,355
=|355,356
=|356,357
=|357,358
=|358,359
=|359,360
=|360,361
=|361,362
=|362,363
=|363,364
=|364,365
=|365,366
=|366,367
=|367,368
=|368,369
=|369,370
=|370,371
=|371,372
=|372,373
=|373,374
=|374,375
=|375,376
=|376,377
=|377,378
=|378,379
=|379,380
=|380,381
=|381,382
=|382,383
<EOL>|385,386
_|387,388
_|388,389
_|389,390
FAILURE|391,398
ADMISSION|399,408
NOTE|409,413
<EOL>|415,416
=|417,418
=|418,419
=|419,420
=|420,421
=|421,422
=|422,423
=|423,424
=|424,425
=|425,426
=|426,427
=|427,428
=|428,429
=|429,430
=|430,431
=|431,432
=|432,433
=|433,434
=|434,435
=|435,436
=|436,437
=|437,438
=|438,439
=|439,440
=|440,441
=|441,442
=|442,443
=|443,444
=|444,445
=|445,446
=|446,447
=|447,448
=|448,449
=|449,450
=|450,451
=|451,452
=|452,453
=|453,454
=|454,455
=|455,456
=|456,457
=|457,458
=|458,459
=|459,460
=|460,461
=|461,462
=|462,463
=|463,464
=|464,465
=|465,466
=|466,467
=|467,468
=|468,469
=|469,470
=|470,471
=|471,472
<EOL>|474,475
OUTPATIENT|475,485
CARDIOLOGIST|486,498
:|498,499
_|501,502
_|502,503
_|503,504
.|504,505
,|505,506
MD|507,509
_|510,511
_|511,512
_|512,513
<EOL>|513,514
cardiology|514,524
)|524,525
,|525,526
_|527,528
_|528,529
_|529,530
_|532,533
_|533,534
_|534,535
.|535,536
,|536,537
MD|538,540
(|540,541
CHF|541,544
)|544,545
<EOL>|545,546
PCP|546,549
:|549,550
_|551,552
_|552,553
_|553,554
.|554,555
,|555,556
MD|557,559
<EOL>|560,561
<EOL>|561,562
CHIEF|562,567
COMPLAINT|568,577
:|577,578
Dyspnea|580,587
on|588,590
Exertion|591,599
<EOL>|599,600
HISTORY|600,607
OF|608,610
PRESENTING|611,621
ILLNESS|622,629
:|629,630
<EOL>|632,633
Mr.|633,636
_|637,638
_|638,639
_|639,640
is|641,643
a|644,645
_|646,647
_|647,648
_|648,649
gentleman|650,659
with|660,664
a|665,666
past|667,671
medical|672,679
<EOL>|679,680
history|680,687
pertinent|688,697
for|698,701
HFrEF|702,707
(|708,709
35|709,711
%|711,712
_|713,714
_|714,715
_|715,716
CAD|717,720
s|721,722
/|722,723
p|723,724
CABG|725,729
and|730,733
<EOL>|733,734
subsequent|734,744
PCI|745,748
,|748,749
moderate|750,758
tricuspid|759,768
regurgitation|769,782
,|782,783
right|784,789
<EOL>|789,790
ventricular|790,801
dysfunction|802,813
,|813,814
moderate|815,823
pulmonary|824,833
hypertension|834,846
,|846,847
and|848,851
<EOL>|851,852
paroxysmal|852,862
atrial|863,869
fibrillation|870,882
on|883,885
apixaban|886,894
,|894,895
stage|896,901
III|902,905
chronic|906,913
<EOL>|913,914
kidney|914,920
disease|921,928
(|929,930
Baseline|930,938
Cr|939,941
2.0|942,945
-|945,946
2.1|946,949
)|949,950
,|950,951
cerebrovascular|952,967
disease|968,975
,|975,976
<EOL>|976,977
and|977,980
metastatic|981,991
melanoma|992,1000
of|1001,1003
unknown|1004,1011
primary|1012,1019
on|1020,1022
checkpoint|1023,1033
<EOL>|1033,1034
inhibitor|1034,1043
pembrolizumab|1044,1057
who|1058,1061
was|1062,1065
found|1066,1071
volume|1072,1078
overloaded|1079,1089
with|1090,1094
<EOL>|1094,1095
increased|1095,1104
DOE|1105,1108
,|1108,1109
admitted|1110,1118
to|1119,1121
_|1122,1123
_|1123,1124
_|1124,1125
for|1126,1129
IV|1130,1132
diuresis|1133,1141
.|1141,1142
<EOL>|1143,1144
<EOL>|1144,1145
Per|1145,1148
most|1149,1153
recent|1154,1160
outpatient|1161,1171
CHF|1172,1175
notes|1176,1181
:|1181,1182
<EOL>|1182,1183
<EOL>|1183,1184
He|1184,1186
was|1187,1190
seen|1191,1195
by|1196,1198
his|1199,1202
primary|1203,1210
car|1211,1214
primary|1215,1222
Cardiologist|1223,1235
,|1235,1236
Dr.|1237,1240
_|1241,1242
_|1242,1243
_|1243,1244
increased|1245,1254
fatigue|1255,1262
and|1263,1266
exertional|1267,1277
dyspnea|1278,1285
.|1285,1286
Dr.|1287,1290
_|1291,1292
_|1292,1293
_|1293,1294
<EOL>|1295,1296
a|1296,1297
<EOL>|1297,1298
_|1298,1299
_|1299,1300
_|1300,1301
and|1302,1305
felt|1306,1310
his|1311,1314
LVEF|1315,1319
was|1320,1323
~|1324,1325
30|1325,1327
%|1327,1328
and|1329,1332
reduced|1333,1340
from|1341,1345
prior|1346,1351
.|1351,1352
He|1353,1355
was|1356,1359
<EOL>|1359,1360
started|1360,1367
on|1368,1370
low|1371,1374
-|1374,1375
dose|1375,1379
Entresto|1380,1388
,|1388,1389
but|1390,1393
could|1394,1399
n't|1399,1402
tolerate|1403,1411
it|1412,1414
from|1415,1419
a|1420,1421
BP|1422,1424
<EOL>|1424,1425
prospective|1425,1436
.|1436,1437
He|1438,1440
was|1441,1444
previously|1445,1455
on|1456,1458
losartan|1459,1467
which|1468,1473
was|1474,1477
stopped|1478,1485
<EOL>|1485,1486
due|1486,1489
to|1490,1492
this|1493,1497
lightheadedness|1498,1513
,|1513,1514
dizziness|1515,1524
and|1525,1528
worsening|1529,1538
renal|1539,1544
<EOL>|1544,1545
function|1545,1553
.|1553,1554
Dr.|1555,1558
_|1559,1560
_|1560,1561
_|1561,1562
concern|1563,1570
about|1571,1576
the|1577,1580
possibility|1581,1592
of|1593,1595
<EOL>|1595,1596
myocarditis|1596,1607
secondary|1608,1617
to|1618,1620
the|1621,1624
checkpoint|1625,1635
inhibitor|1636,1645
.|1645,1646
When|1647,1651
he|1652,1654
<EOL>|1654,1655
followed|1655,1663
up|1664,1666
with|1667,1671
the|1672,1675
Oncology|1676,1684
team|1685,1689
on|1690,1692
_|1693,1694
_|1694,1695
_|1695,1696
,|1696,1697
his|1698,1701
symptoms|1702,1710
were|1711,1715
<EOL>|1715,1716
somewhat|1716,1724
improved|1725,1733
.|1733,1734
Cardiac|1735,1742
biomarkers|1743,1753
were|1754,1758
notable|1759,1766
for|1767,1770
a|1771,1772
rising|1773,1779
<EOL>|1779,1780
NTproBNP|1780,1788
to|1789,1791
>|1792,1793
10K|1793,1796
but|1797,1800
normal|1801,1807
CK|1808,1810
-|1810,1811
MB|1811,1813
and|1814,1817
minimally|1818,1827
elevated|1828,1836
<EOL>|1837,1838
troponin|1838,1846
<EOL>|1846,1847
T|1847,1848
of|1849,1851
0.03|1852,1856
,|1856,1857
which|1858,1863
is|1864,1866
not|1867,1870
unexpected|1871,1881
in|1882,1884
the|1885,1888
setting|1889,1896
<EOL>|1896,1897
of|1897,1899
decompensated|1900,1913
_|1914,1915
_|1915,1916
_|1916,1917
failure|1918,1925
and|1926,1929
chronic|1930,1937
kidney|1938,1944
disease|1945,1952
.|1952,1953
He|1954,1956
<EOL>|1957,1958
was|1958,1961
<EOL>|1961,1962
planned|1962,1969
to|1970,1972
receive|1973,1980
immunotherapy|1981,1994
on|1995,1997
_|1998,1999
_|1999,2000
_|2000,2001
,|2001,2002
but|2003,2006
treatment|2007,2016
was|2017,2020
<EOL>|2020,2021
held|2021,2025
due|2026,2029
to|2030,2032
elevated|2033,2041
Cr|2042,2044
.|2044,2045
Recheck|2046,2053
showed|2054,2060
improvement|2061,2072
.|2072,2073
The|2074,2077
patient|2078,2085
<EOL>|2085,2086
restarted|2086,2095
pembrolizumab|2096,2109
on|2110,2112
_|2113,2114
_|2114,2115
_|2115,2116
.|2116,2117
Pembrolizumab|2118,2131
was|2132,2135
again|2136,2141
<EOL>|2142,2143
held|2143,2147
<EOL>|2147,2148
in|2148,2150
_|2151,2152
_|2152,2153
_|2153,2154
for|2155,2158
diarrhea|2159,2167
and|2168,2171
elevated|2172,2180
LFTs|2181,2185
<EOL>|2186,2187
<EOL>|2187,2188
In|2188,2190
addition|2191,2199
,|2199,2200
he|2201,2203
also|2204,2208
received|2209,2217
intravenous|2218,2229
hydration|2230,2239
.|2239,2240
<EOL>|2240,2241
Subsequently|2241,2253
,|2253,2254
he|2255,2257
was|2258,2261
noted|2262,2267
to|2268,2270
be|2271,2273
more|2274,2278
volume|2279,2285
overloaded|2286,2296
,|2296,2297
at|2298,2300
<EOL>|2301,2302
which|2302,2307
<EOL>|2307,2308
time|2308,2312
Torsemide|2313,2322
from|2323,2327
20|2328,2330
mg|2331,2333
daily|2334,2339
to|2340,2342
30|2343,2345
mg|2346,2348
daily|2349,2354
then|2355,2359
40|2360,2362
mg|2363,2365
daily|2366,2371
.|2371,2372
<EOL>|2372,2373
Troponin|2373,2381
testing|2382,2389
showed|2390,2396
Trop|2397,2401
-|2401,2402
T|2402,2403
of|2404,2406
0.04|2407,2411
,|2411,2412
attributed|2413,2423
to|2424,2426
renal|2427,2432
<EOL>|2432,2433
insufficiency|2433,2446
.|2446,2447
The|2448,2451
patient|2452,2459
was|2460,2463
also|2464,2468
noted|2469,2474
to|2475,2477
have|2478,2482
mild|2483,2487
<EOL>|2487,2488
hyperkalemia|2488,2500
(|2501,2502
K|2502,2503
5.7|2504,2507
)|2507,2508
for|2509,2512
which|2513,2518
potassium|2519,2528
supplementation|2529,2544
was|2545,2548
<EOL>|2548,2549
stopped|2549,2556
and|2557,2560
torsemide|2561,2570
dose|2571,2575
increased|2576,2585
.|2585,2586
He|2587,2589
was|2590,2593
also|2594,2598
seen|2599,2603
in|2604,2606
the|2607,2610
<EOL>|2610,2611
Emergency|2611,2620
room|2621,2625
in|2626,2628
the|2629,2632
_|2633,2634
_|2634,2635
_|2635,2636
_|2637,2638
_|2638,2639
_|2639,2640
due|2641,2644
to|2645,2647
a|2648,2649
<EOL>|2649,2650
fall|2650,2654
with|2655,2659
resultant|2660,2669
scalp|2670,2675
laceration|2676,2686
.|2686,2687
CT|2688,2690
head|2691,2695
and|2696,2699
neck|2700,2704
was|2705,2708
<EOL>|2708,2709
unremarkable|2709,2721
.|2721,2722
<EOL>|2723,2724
<EOL>|2724,2725
He|2725,2727
presented|2728,2737
this|2738,2742
morning|2743,2750
_|2751,2752
_|2752,2753
_|2753,2754
for|2755,2758
his|2759,2762
scheduled|2763,2772
visit|2773,2778
at|2779,2781
<EOL>|2781,2782
_|2782,2783
_|2783,2784
_|2784,2785
clinic|2786,2792
where|2793,2798
he|2799,2801
noted|2802,2807
that|2808,2812
his|2813,2816
weight|2817,2823
had|2824,2827
been|2828,2832
126|2833,2836
lbs|2837,2840
most|2841,2845
<EOL>|2845,2846
recently|2846,2854
on|2855,2857
his|2858,2861
home|2862,2866
scale|2867,2872
.|2872,2873
He|2874,2876
also|2877,2881
reported|2882,2890
decreased|2891,2900
appetite|2901,2909
<EOL>|2909,2910
that|2910,2914
he|2915,2917
attributes|2918,2928
to|2929,2931
eating|2932,2938
a|2939,2940
different|2941,2950
diet|2951,2955
.|2955,2956
He|2957,2959
currently|2960,2969
has|2970,2973
<EOL>|2974,2975
a|2975,2976
<EOL>|2976,2977
_|2977,2978
_|2978,2979
_|2979,2980
care|2981,2985
taker|2986,2991
that|2992,2996
makes|2997,3002
_|3003,3004
_|3004,3005
_|3005,3006
food|3007,3011
for|3012,3015
him|3016,3019
,|3019,3020
adhering|3021,3029
<EOL>|3029,3030
to|3030,3032
a|3033,3034
low|3035,3038
sodium|3039,3045
diet|3046,3050
,|3050,3051
that|3052,3056
he|3057,3059
does|3060,3064
not|3065,3068
like|3069,3073
as|3074,3076
much|3077,3081
as|3082,3084
his|3085,3088
<EOL>|3088,3089
regular|3089,3096
diet|3097,3101
.|3101,3102
He|3103,3105
drinks|3106,3112
_|3113,3114
_|3114,3115
_|3115,3116
glasses|3117,3124
of|3125,3127
water|3128,3133
or|3134,3136
juice|3137,3142
daily|3143,3148
.|3148,3149
He|3150,3152
<EOL>|3152,3153
was|3153,3156
taking|3157,3163
torsemide|3164,3173
40|3174,3176
mg|3177,3179
daily|3180,3185
,|3185,3186
that|3187,3191
he|3192,3194
decreased|3195,3204
to|3205,3207
30|3208,3210
mg|3211,3213
<EOL>|3213,3214
daily|3214,3219
several|3220,3227
days|3228,3232
ago|3233,3236
as|3237,3239
he|3240,3242
felt|3243,3247
he|3248,3250
was|3251,3254
urinating|3255,3264
too|3265,3268
<EOL>|3268,3269
frequently|3269,3279
.|3279,3280
He|3281,3283
also|3284,3288
ran|3289,3292
out|3293,3296
of|3297,3299
tamsulosin|3300,3310
several|3311,3318
days|3319,3323
ago|3324,3327
so|3328,3330
<EOL>|3330,3331
stopped|3331,3338
taking|3339,3345
this|3346,3350
around|3351,3357
the|3358,3361
same|3362,3366
time|3367,3371
.|3371,3372
He|3373,3375
noted|3376,3381
becoming|3382,3390
<EOL>|3391,3392
short|3392,3397
<EOL>|3397,3398
of|3398,3400
breath|3401,3407
after|3408,3413
taking|3414,3420
20|3421,3423
steps|3424,3429
or|3430,3432
less|3433,3437
.|3437,3438
Due|3439,3442
to|3443,3445
his|3446,3449
volume|3450,3456
<EOL>|3456,3457
overloaded|3457,3467
noted|3468,3473
on|3474,3476
exam|3477,3481
he|3482,3484
was|3485,3488
recommended|3489,3500
for|3501,3504
admission|3505,3514
to|3515,3517
_|3518,3519
_|3519,3520
_|3520,3521
<EOL>|3521,3522
for|3522,3525
IV|3526,3528
diuresis|3529,3537
<EOL>|3537,3538
<EOL>|3538,3539
On|3539,3541
the|3542,3545
floor|3546,3551
,|3551,3552
he|3553,3555
endorses|3556,3564
the|3565,3568
above|3569,3574
history|3575,3582
.|3582,3583
He|3584,3586
noted|3587,3592
that|3593,3597
his|3598,3601
<EOL>|3601,3602
SOB|3602,3605
has|3606,3609
progressive|3610,3621
gotten|3622,3628
worse|3629,3634
.|3634,3635
Mostly|3636,3642
occurs|3643,3649
with|3650,3654
activity|3655,3663
.|3663,3664
<EOL>|3664,3665
None|3665,3669
at|3670,3672
rest|3673,3677
.|3677,3678
He|3679,3681
noted|3682,3687
that|3688,3692
his|3693,3696
weight|3697,3703
has|3704,3707
been|3708,3712
slowly|3713,3719
<EOL>|3720,3721
decreasing|3721,3731
<EOL>|3731,3732
due|3732,3735
lack|3736,3740
of|3741,3743
appetite|3744,3752
and|3753,3756
him|3757,3760
being|3761,3766
to|3767,3769
lazy|3770,3774
.|3774,3775
He|3776,3778
has|3779,3782
a|3783,3784
home|3785,3789
health|3790,3796
<EOL>|3796,3797
aid|3797,3800
everyday|3801,3809
from|3810,3814
11am|3815,3819
-|3819,3820
7pm|3820,3823
,|3823,3824
who|3825,3828
helps|3829,3834
him|3835,3838
with|3839,3843
ADL|3844,3847
.|3847,3848
He|3850,3852
endorses|3853,3861
<EOL>|3861,3862
abdominal|3862,3871
bloading|3872,3880
.|3880,3881
<EOL>|3882,3883
<EOL>|3883,3884
Cardiac|3884,3891
review|3892,3898
of|3899,3901
systems|3902,3909
is|3910,3912
notable|3913,3920
for|3921,3924
absence|3925,3932
of|3933,3935
chest|3936,3941
pain|3942,3946
,|3946,3947
<EOL>|3947,3948
paroxysmal|3948,3958
nocturnal|3959,3968
dyspnea|3969,3976
,|3976,3977
orthopnea|3978,3987
,|3987,3988
palpitations|3989,4001
,|4001,4002
syncope|4003,4010
,|4010,4011
<EOL>|4011,4012
or|4012,4014
presyncope|4015,4025
.|4025,4026
<EOL>|4026,4027
<EOL>|4027,4028
ROS|4028,4031
otherwise|4032,4041
negative|4042,4050
,|4050,4051
unless|4052,4058
otherwise|4059,4068
noted|4069,4074
above|4075,4080
<EOL>|4081,4082
<EOL>|4082,4083
<EOL>|4084,4085
Past|4085,4089
Medical|4090,4097
History|4098,4105
:|4105,4106
<EOL>|4106,4107
Past|4107,4111
Medical|4112,4119
History|4120,4127
:|4127,4128
<EOL>|4128,4129
BILATERAL|4129,4138
MODERATE|4139,4147
CAROTID|4148,4155
DISEASE|4156,4163
<EOL>|4164,4165
CONGESTIVE|4165,4175
_|4176,4177
_|4177,4178
_|4178,4179
FAILURE|4180,4187
<EOL>|4188,4189
CORONARY|4189,4197
ARTERY|4198,4204
DISEASE|4205,4212
<EOL>|4213,4214
GASTROESOPHAGEAL|4214,4230
REFLUX|4231,4237
<EOL>|4238,4239
HYPERTENSION|4239,4251
<EOL>|4252,4253
SEVERE|4253,4259
EMPHYSEMA|4260,4269
<EOL>|4270,4271
PULMONARY|4271,4280
HYPERTENSION|4281,4293
<EOL>|4294,4295
RIGHT|4295,4300
BUNDLE|4301,4307
BRANCH|4308,4314
BLOCK|4315,4320
<EOL>|4321,4322
BENIGN|4322,4328
PROSTATIC|4329,4338
HYPERTROPHY|4339,4350
<EOL>|4351,4352
HYPERLIPIDEMIA|4352,4366
<EOL>|4367,4368
PAROXYSMAL|4368,4378
ATRIAL|4379,4385
FIBRILLATION|4386,4398
<EOL>|4399,4400
H|4400,4401
/|4401,4402
O|4402,4403
HISTIOPLASMOSIS|4404,4419
<EOL>|4420,4421
<EOL>|4421,4422
Past|4422,4426
Surgical|4427,4435
History|4436,4443
:|4443,4444
<EOL>|4444,4445
CARDIOVERSION|4445,4458
_|4459,4460
_|4460,4461
_|4461,4462
<EOL>|4463,4464
RIGHT|4464,4469
LOWER|4470,4475
LOBE|4476,4480
LOBECTOMY|4481,4490
_|4491,4492
_|4492,4493
_|4493,4494
<EOL>|4495,4496
CORONARY|4496,4504
BYPASS|4505,4511
SURGERY|4512,4519
_|4520,4521
_|4521,4522
_|4522,4523
<EOL>|4524,4525
<EOL>|4525,4526
<EOL>|4527,4528
Social|4528,4534
History|4535,4542
:|4542,4543
<EOL>|4543,4544
_|4544,4545
_|4545,4546
_|4546,4547
<EOL>|4547,4548
Family|4548,4554
History|4555,4562
:|4562,4563
<EOL>|4563,4564
Non-contributory|4564,4580
<EOL>|4580,4581
<EOL>|4582,4583
Physical|4583,4591
Exam|4592,4596
:|4596,4597
<EOL>|4597,4598
ADMISSION|4598,4607
PHYSICAL|4608,4616
EXAMINATION|4617,4628
:|4628,4629
<EOL>|4629,4630
=|4630,4631
=|4631,4632
=|4632,4633
=|4633,4634
=|4634,4635
=|4635,4636
=|4636,4637
=|4637,4638
=|4638,4639
=|4639,4640
=|4640,4641
=|4641,4642
=|4642,4643
=|4643,4644
=|4644,4645
=|4645,4646
=|4646,4647
=|4647,4648
=|4648,4649
=|4649,4650
=|4650,4651
=|4651,4652
=|4652,4653
=|4653,4654
=|4654,4655
=|4655,4656
=|4656,4657
=|4657,4658
=|4658,4659
=|4659,4660
=|4660,4661
<EOL>|4661,4662
24|4662,4664
HR|4665,4667
Data|4668,4672
(|4673,4674
last|4674,4678
updated|4679,4686
_|4687,4688
_|4688,4689
_|4689,4690
@|4691,4692
1335|4693,4697
)|4697,4698
<EOL>|4698,4699
Temp|4703,4707
:|4707,4708
97.4|4709,4713
(|4714,4715
Tm|4715,4717
97.4|4718,4722
)|4722,4723
,|4723,4724
BP|4725,4727
:|4727,4728
115|4729,4732
/|4732,4733
66|4733,4735
,|4735,4736
HR|4737,4739
:|4739,4740
61|4741,4743
,|4743,4744
RR|4745,4747
:|4747,4748
18|4749,4751
,|4751,4752
O2|4753,4755
sat|4756,4759
:|4759,4760
<EOL>|4760,4761
99|4761,4763
%|4763,4764
,|4764,4765
O2|4766,4768
delivery|4769,4777
:|4777,4778
ra|4779,4781
,|4781,4782
Wt|4783,4785
:|4785,4786
130.73|4787,4793
lb|4794,4796
/|4796,4797
59.3|4797,4801
kg|4802,4804
<EOL>|4806,4807
<EOL>|4807,4808
GENERAL|4808,4815
:|4815,4816
Well|4817,4821
developed|4822,4831
,|4831,4832
well|4833,4837
nourished|4838,4847
male|4848,4852
in|4853,4855
NAD|4856,4859
.|4859,4860
Oriented|4861,4869
<EOL>|4870,4871
x3|4871,4873
.|4873,4874
<EOL>|4874,4875
Mood|4875,4879
,|4879,4880
affect|4881,4887
appropriate|4888,4899
.|4899,4900
<EOL>|4902,4903
HEENT|4903,4908
:|4908,4909
Scalp|4910,4915
laceration|4916,4926
noted|4927,4932
.|4932,4933
Sclera|4934,4940
slightly|4941,4949
icteric|4950,4957
.|4957,4958
PERRL|4959,4964
.|4964,4965
<EOL>|4965,4966
EOMI|4966,4970
.|4970,4971
Conjunctiva|4972,4983
were|4984,4988
pink|4989,4993
.|4993,4994
No|4995,4997
pallor|4998,5004
or|5005,5007
cyanosis|5008,5016
of|5017,5019
the|5020,5023
oral|5024,5028
<EOL>|5028,5029
mucosa|5029,5035
.|5035,5036
No|5037,5039
xanthelasma|5040,5051
.|5051,5052
<EOL>|5054,5055
NECK|5055,5059
:|5059,5060
Supple|5061,5067
.|5067,5068
JVP|5069,5072
~|5073,5074
20|5075,5077
cm|5078,5080
with|5081,5085
positive|5086,5094
hepatojugular|5095,5108
reflex|5109,5115
.|5115,5116
<EOL>|5117,5118
CARDIAC|5118,5125
:|5125,5126
Regular|5127,5134
rate|5135,5139
and|5140,5143
rhythm|5144,5150
.|5150,5151
Normal|5152,5158
S1|5159,5161
,|5161,5162
S2|5163,5165
.|5165,5166
_|5167,5168
_|5168,5169
_|5169,5170
<EOL>|5171,5172
holosystolic|5172,5184
<EOL>|5184,5185
murmur|5185,5191
at|5192,5194
the|5195,5198
LLSB|5199,5203
and|5204,5207
the|5208,5211
apex|5212,5216
,|5216,5217
no|5218,5220
rubs|5221,5225
,|5225,5226
or|5227,5229
gallops|5230,5237
.|5237,5238
No|5239,5241
thrills|5242,5249
<EOL>|5249,5250
or|5250,5252
lifts|5253,5258
.|5258,5259
<EOL>|5261,5262
LUNGS|5262,5267
:|5267,5268
No|5269,5271
chest|5272,5277
wall|5278,5282
deformities|5283,5294
or|5295,5297
tenderness|5298,5308
.|5308,5309
Respiration|5310,5321
is|5322,5324
<EOL>|5324,5325
unlabored|5325,5334
with|5335,5339
no|5340,5342
accessory|5343,5352
muscle|5353,5359
use|5360,5363
.|5363,5364
Bibasilar|5365,5374
crackles|5375,5383
<EOL>|5384,5385
ABDOMEN|5385,5392
:|5392,5393
mildly|5394,5400
distended|5401,5410
;|5410,5411
normoactive|5412,5423
bowel|5424,5429
sounds|5430,5436
;|5436,5437
soft|5438,5442
and|5443,5446
<EOL>|5446,5447
non-tender|5447,5457
to|5458,5460
palpation|5461,5470
;|5470,5471
there|5472,5477
is|5478,5480
no|5481,5483
appreciable|5484,5495
organomegaly|5496,5508
or|5509,5511
<EOL>|5511,5512
mass|5512,5516
<EOL>|5516,5517
EXTREMITIES|5517,5528
:|5528,5529
Cool|5530,5534
,|5534,5535
1|5536,5537
+|5537,5538
pitting|5539,5546
edema|5547,5552
to|5553,5555
knee|5556,5560
caps|5561,5565
.|5565,5566
bilateral|5567,5576
<EOL>|5576,5577
status|5577,5583
dermatitis|5584,5594
.|5594,5595
<EOL>|5596,5597
SKIN|5597,5601
:|5601,5602
Eccymosis|5603,5612
noted|5613,5618
on|5619,5621
left|5622,5626
hand|5627,5631
,|5631,5632
Multiple|5633,5641
open|5642,5646
biopsy|5647,5653
<EOL>|5654,5655
excision|5655,5663
<EOL>|5663,5664
sites|5664,5669
on|5670,5672
left|5673,5677
shin|5678,5682
and|5683,5686
right|5687,5692
calf|5693,5697
<EOL>|5697,5698
PULSES|5698,5704
:|5704,5705
Distal|5706,5712
pulses|5713,5719
palpable|5720,5728
and|5729,5732
symmetric|5733,5742
.|5742,5743
<EOL>|5744,5745
<EOL>|5745,5746
Discharge|5746,5755
Physical|5756,5764
exam|5765,5769
<EOL>|5769,5770
=|5770,5771
=|5771,5772
=|5772,5773
=|5773,5774
=|5774,5775
=|5775,5776
=|5776,5777
=|5777,5778
=|5778,5779
=|5779,5780
=|5780,5781
=|5781,5782
=|5782,5783
=|5783,5784
=|5784,5785
=|5785,5786
=|5786,5787
=|5787,5788
=|5788,5789
=|5789,5790
=|5790,5791
=|5791,5792
=|5792,5793
<EOL>|5793,5794
24|5794,5796
HR|5797,5799
Data|5800,5804
(|5805,5806
last|5806,5810
updated|5811,5818
_|5819,5820
_|5820,5821
_|5821,5822
@|5823,5824
751|5825,5828
)|5828,5829
<EOL>|5829,5830
Temp|5834,5838
:|5838,5839
98.2|5840,5844
(|5845,5846
Tm|5846,5848
98.6|5849,5853
)|5853,5854
,|5854,5855
BP|5856,5858
:|5858,5859
110|5860,5863
/|5863,5864
61|5864,5866
(|5867,5868
100|5868,5871
-|5871,5872
121|5872,5875
/|5875,5876
54|5876,5878
-|5878,5879
63|5879,5881
)|5881,5882
,|5882,5883
HR|5884,5886
:|5886,5887
72|5888,5890
<EOL>|5890,5891
(|5891,5892
60|5892,5894
-|5894,5895
99|5895,5897
)|5897,5898
,|5898,5899
RR|5900,5902
:|5902,5903
16|5904,5906
(|5907,5908
_|5908,5909
_|5909,5910
_|5910,5911
)|5911,5912
,|5912,5913
O2|5914,5916
sat|5917,5920
:|5920,5921
91|5922,5924
%|5924,5925
(|5926,5927
91|5927,5929
-|5929,5930
95|5930,5932
)|5932,5933
,|5933,5934
O2|5935,5937
delivery|5938,5946
:|5946,5947
Ra|5948,5950
<EOL>|5952,5953
<EOL>|5953,5954
General|5954,5961
:|5961,5962
elderly|5963,5970
gentleman|5971,5980
in|5981,5983
NAD|5984,5987
<EOL>|5987,5988
HEENT|5988,5993
:|5993,5994
dressing|5995,6003
in|6004,6006
place|6007,6012
on|6013,6015
scalp|6016,6021
from|6022,6026
recent|6027,6033
fall|6034,6038
/|6038,6039
scalp|6039,6044
<EOL>|6044,6045
laceration|6045,6055
/|6055,6056
c|6056,6057
/|6057,6058
d|6058,6059
/|6059,6060
i|6060,6061
.|6061,6062
Sclera|6063,6069
mildly|6070,6076
icteric|6077,6084
,|6084,6085
pupils|6086,6092
equally|6093,6100
round|6101,6106
,|6106,6107
<EOL>|6107,6108
MMM|6108,6111
<EOL>|6112,6113
NECK|6113,6117
:|6117,6118
JVP|6119,6122
~|6122,6123
10cm|6123,6127
,|6127,6128
with|6129,6133
positive|6134,6142
hepatojugular|6143,6156
reflex|6157,6163
<EOL>|6163,6164
CV|6164,6166
:|6166,6167
irregularly|6169,6180
irregular|6181,6190
;|6191,6192
the|6193,6196
precordium|6197,6207
is|6208,6210
quiet|6211,6216
without|6217,6224
RV|6225,6227
<EOL>|6227,6228
heave|6228,6233
;|6233,6234
normal|6235,6241
S1|6242,6244
with|6245,6249
fixed|6250,6255
split|6256,6261
S2|6262,6264
;|6264,6265
there|6266,6271
is|6272,6274
a|6275,6276
soft|6277,6281
_|6282,6283
_|6283,6284
_|6284,6285
<EOL>|6285,6286
holosystolic|6286,6298
<EOL>|6298,6299
murmur|6299,6305
at|6306,6308
the|6309,6312
LLSB|6313,6317
and|6318,6321
the|6322,6325
apex|6326,6330
;|6330,6331
<EOL>|6331,6332
LUNGS|6332,6337
:|6337,6338
Normal|6339,6345
effort|6346,6352
.|6352,6353
Fine|6354,6358
Bibasilar|6359,6368
crackles|6369,6377
<EOL>|6377,6378
Abd|6378,6381
:|6381,6382
soft|6383,6387
,|6387,6388
mildy|6389,6394
distended|6395,6404
,|6404,6405
no|6406,6408
guarding|6409,6417
/|6418,6419
rebound|6420,6427
.|6427,6428
<EOL>|6429,6430
EXT|6430,6433
:|6433,6434
1|6436,6437
+|6437,6438
pitting|6439,6446
edema|6447,6452
to|6453,6455
the|6456,6459
mid-calf|6460,6468
L|6469,6470
leg|6471,6474
>|6475,6476
R|6477,6478
leg|6479,6482
<EOL>|6482,6483
SKIN|6483,6487
:|6487,6488
Multiple|6490,6498
excision|6499,6507
biopsy|6508,6514
wounds|6515,6521
on|6522,6524
legs|6525,6529
,|6529,6530
covered|6531,6538
with|6539,6543
<EOL>|6543,6544
dressing|6544,6552
c|6553,6554
/|6554,6555
d|6555,6556
/|6556,6557
i|6557,6558
<EOL>|6558,6559
NEURO|6559,6564
:|6564,6565
Speech|6567,6573
fluent|6574,6580
,|6580,6581
strength|6582,6590
grossly|6591,6598
intact|6599,6605
<EOL>|6606,6607
<EOL>|6607,6608
<EOL>|6609,6610
Pertinent|6610,6619
Results|6620,6627
:|6627,6628
<EOL>|6628,6629
_|6629,6630
_|6630,6631
_|6631,6632
01|6633,6635
:|6635,6636
00PM|6636,6640
_|6643,6644
_|6644,6645
_|6645,6646
PTT|6647,6650
-|6650,6651
34.4|6651,6655
_|6656,6657
_|6657,6658
_|6658,6659
<EOL>|6659,6660
_|6660,6661
_|6661,6662
_|6662,6663
01|6664,6666
:|6666,6667
00PM|6667,6671
PLT|6674,6677
COUNT|6678,6683
-|6683,6684
169|6684,6687
<EOL>|6687,6688
_|6688,6689
_|6689,6690
_|6690,6691
01|6692,6694
:|6694,6695
00PM|6695,6699
NEUTS|6702,6707
-|6707,6708
81|6708,6710
.|6710,6711
6|6711,6712
*|6712,6713
LYMPHS|6714,6720
-|6720,6721
6|6721,6722
.|6722,6723
6|6723,6724
*|6724,6725
MONOS|6726,6731
-|6731,6732
10.4|6732,6736
EOS|6737,6740
-|6740,6741
0|6741,6742
.|6742,6743
1|6743,6744
*|6744,6745
<EOL>|6746,6747
BASOS|6747,6752
-|6752,6753
0.1|6753,6756
IM|6757,6759
_|6760,6761
_|6761,6762
_|6762,6763
AbsNeut|6764,6771
-|6771,6772
6.00|6772,6776
AbsLymp|6777,6784
-|6784,6785
0|6785,6786
.|6786,6787
49|6787,6789
*|6789,6790
AbsMono|6791,6798
-|6798,6799
0|6799,6800
.|6800,6801
77|6801,6803
<EOL>|6804,6805
AbsEos|6805,6811
-|6811,6812
0|6812,6813
.|6813,6814
01|6814,6816
*|6816,6817
AbsBaso|6818,6825
-|6825,6826
0.01|6826,6830
<EOL>|6830,6831
_|6831,6832
_|6832,6833
_|6833,6834
01|6835,6837
:|6837,6838
00PM|6838,6842
WBC|6845,6848
-|6848,6849
7.4|6849,6852
RBC|6853,6856
-|6856,6857
3|6857,6858
.|6858,6859
02|6859,6861
*|6861,6862
HGB|6863,6866
-|6866,6867
9|6867,6868
.|6868,6869
1|6869,6870
*|6870,6871
HCT|6872,6875
-|6875,6876
30|6876,6878
.|6878,6879
2|6879,6880
*|6880,6881
MCV|6882,6885
-|6885,6886
100|6886,6889
*|6889,6890
<EOL>|6891,6892
MCH|6892,6895
-|6895,6896
30.1|6896,6900
MCHC|6901,6905
-|6905,6906
30|6906,6908
.|6908,6909
1|6909,6910
*|6910,6911
RDW|6912,6915
-|6915,6916
16|6916,6918
.|6918,6919
4|6919,6920
*|6920,6921
RDWSD|6922,6927
-|6927,6928
59|6928,6930
.|6930,6931
2|6931,6932
*|6932,6933
<EOL>|6933,6934
_|6934,6935
_|6935,6936
_|6936,6937
01|6938,6940
:|6940,6941
00PM|6941,6945
calTIBC|6948,6955
-|6955,6956
352|6956,6959
FERRITIN|6960,6968
-|6968,6969
111|6969,6972
TRF|6973,6976
-|6976,6977
271|6977,6980
<EOL>|6980,6981
_|6981,6982
_|6982,6983
_|6983,6984
01|6985,6987
:|6987,6988
00PM|6988,6992
CALCIUM|6995,7002
-|7002,7003
9.2|7003,7006
PHOSPHATE|7007,7016
-|7016,7017
3.7|7017,7020
MAGNESIUM|7021,7030
-|7030,7031
2|7031,7032
.|7032,7033
8|7033,7034
*|7034,7035
<EOL>|7036,7037
IRON|7037,7041
-|7041,7042
88|7042,7044
<EOL>|7044,7045
_|7045,7046
_|7046,7047
_|7047,7048
01|7049,7051
:|7051,7052
00PM|7052,7056
CK|7059,7061
-|7061,7062
MB|7062,7064
-|7064,7065
4|7065,7066
cTropnT|7067,7074
-|7074,7075
0|7075,7076
.|7076,7077
01|7077,7079
_|7080,7081
_|7081,7082
_|7082,7083
<EOL>|7083,7084
_|7084,7085
_|7085,7086
_|7086,7087
01|7088,7090
:|7090,7091
00PM|7091,7095
ALT|7098,7101
(|7101,7102
SGPT|7102,7106
)|7106,7107
-|7107,7108
56|7108,7110
*|7110,7111
AST|7112,7115
(|7115,7116
SGOT|7116,7120
)|7120,7121
-|7121,7122
52|7122,7124
*|7124,7125
LD|7126,7128
(|7128,7129
LDH|7129,7132
)|7132,7133
-|7133,7134
277|7134,7137
*|7137,7138
ALK|7139,7142
<EOL>|7143,7144
PHOS|7144,7148
-|7148,7149
135|7149,7152
*|7152,7153
TOT|7154,7157
BILI|7158,7162
-|7162,7163
0.7|7163,7166
<EOL>|7166,7167
_|7167,7168
_|7168,7169
_|7169,7170
01|7171,7173
:|7173,7174
00PM|7174,7178
estGFR|7181,7187
-|7187,7188
Using|7188,7193
this|7194,7198
<EOL>|7198,7199
_|7199,7200
_|7200,7201
_|7201,7202
01|7203,7205
:|7205,7206
00PM|7206,7210
GLUCOSE|7213,7220
-|7220,7221
100|7221,7224
UREA|7225,7229
N|7230,7231
-|7231,7232
52|7232,7234
*|7234,7235
CREAT|7236,7241
-|7241,7242
2|7242,7243
.|7243,7244
1|7244,7245
*|7245,7246
SODIUM|7247,7253
-|7253,7254
135|7254,7257
<EOL>|7258,7259
POTASSIUM|7259,7268
-|7268,7269
5.4|7269,7272
CHLORIDE|7273,7281
-|7281,7282
100|7282,7285
TOTAL|7286,7291
CO2|7292,7295
-|7295,7296
24|7296,7298
ANION|7299,7304
GAP|7305,7308
-|7308,7309
11|7309,7311
<EOL>|7311,7312
_|7312,7313
_|7313,7314
_|7314,7315
04|7316,7318
:|7318,7319
54PM|7319,7323
URINE|7324,7329
HYALINE|7331,7338
-|7338,7339
1|7339,7340
*|7340,7341
<EOL>|7341,7342
_|7342,7343
_|7343,7344
_|7344,7345
04|7346,7348
:|7348,7349
54PM|7349,7353
URINE|7354,7359
RBC|7361,7364
-|7364,7365
0|7365,7366
WBC|7367,7370
-|7370,7371
<|7371,7372
1|7372,7373
BACTERIA|7374,7382
-|7382,7383
NONE|7383,7387
YEAST|7388,7393
-|7393,7394
NONE|7394,7398
<EOL>|7399,7400
EPI|7400,7403
-|7403,7404
<|7404,7405
1|7405,7406
<EOL>|7406,7407
_|7407,7408
_|7408,7409
_|7409,7410
04|7411,7413
:|7413,7414
54PM|7414,7418
URINE|7419,7424
BLOOD|7426,7431
-|7431,7432
NEG|7432,7435
NITRITE|7436,7443
-|7443,7444
NEG|7444,7447
PROTEIN|7448,7455
-|7455,7456
TR|7456,7458
*|7458,7459
<EOL>|7460,7461
GLUCOSE|7461,7468
-|7468,7469
NEG|7469,7472
KETONE|7473,7479
-|7479,7480
NEG|7480,7483
BILIRUBIN|7484,7493
-|7493,7494
NEG|7494,7497
UROBILNGN|7498,7507
-|7507,7508
NEG|7508,7511
PH|7512,7514
-|7514,7515
7.0|7515,7518
<EOL>|7519,7520
LEUK|7520,7524
-|7524,7525
NEG|7525,7528
<EOL>|7528,7529
_|7529,7530
_|7530,7531
_|7531,7532
04|7533,7535
:|7535,7536
54PM|7536,7540
URINE|7541,7546
COLOR|7548,7553
-|7553,7554
Straw|7554,7559
APPEAR|7560,7566
-|7566,7567
Clear|7567,7572
SP|7573,7575
_|7576,7577
_|7577,7578
_|7578,7579
<EOL>|7579,7580
_|7580,7581
_|7581,7582
_|7582,7583
07|7584,7586
:|7586,7587
53AM|7587,7591
BLOOD|7592,7597
WBC|7598,7601
-|7601,7602
6.5|7602,7605
RBC|7606,7609
-|7609,7610
2|7610,7611
.|7611,7612
70|7612,7614
*|7614,7615
Hgb|7616,7619
-|7619,7620
8|7620,7621
.|7621,7622
2|7622,7623
*|7623,7624
Hct|7625,7628
-|7628,7629
26|7629,7631
.|7631,7632
5|7632,7633
*|7633,7634
<EOL>|7635,7636
MCV|7636,7639
-|7639,7640
98|7640,7642
MCH|7643,7646
-|7646,7647
30.4|7647,7651
MCHC|7652,7656
-|7656,7657
30|7657,7659
.|7659,7660
9|7660,7661
*|7661,7662
RDW|7663,7666
-|7666,7667
16|7667,7669
.|7669,7670
0|7670,7671
*|7671,7672
RDWSD|7673,7678
-|7678,7679
56|7679,7681
.|7681,7682
3|7682,7683
*|7683,7684
Plt|7685,7688
_|7689,7690
_|7690,7691
_|7691,7692
<EOL>|7692,7693
_|7693,7694
_|7694,7695
_|7695,7696
07|7697,7699
:|7699,7700
53AM|7700,7704
BLOOD|7705,7710
Plt|7711,7714
_|7715,7716
_|7716,7717
_|7717,7718
<EOL>|7718,7719
_|7719,7720
_|7720,7721
_|7721,7722
07|7723,7725
:|7725,7726
53AM|7726,7730
BLOOD|7731,7736
Glucose|7737,7744
-|7744,7745
105|7745,7748
*|7748,7749
UreaN|7750,7755
-|7755,7756
43|7756,7758
*|7758,7759
Creat|7760,7765
-|7765,7766
2|7766,7767
.|7767,7768
2|7768,7769
*|7769,7770
Na|7771,7773
-|7773,7774
140|7774,7777
<EOL>|7778,7779
K|7779,7780
-|7780,7781
4.2|7781,7784
Cl|7785,7787
-|7787,7788
102|7788,7791
HCO3|7792,7796
-|7796,7797
27|7797,7799
AnGap|7800,7805
-|7805,7806
11|7806,7808
<EOL>|7808,7809
_|7809,7810
_|7810,7811
_|7811,7812
:|7812,7813
04AM|7813,7817
BLOOD|7818,7823
ALT|7824,7827
-|7827,7828
45|7828,7830
*|7830,7831
AST|7832,7835
-|7835,7836
42|7836,7838
*|7838,7839
AlkPhos|7840,7847
-|7847,7848
113|7848,7851
TotBili|7852,7859
-|7859,7860
0.6|7860,7863
<EOL>|7863,7864
_|7864,7865
_|7865,7866
_|7866,7867
07|7868,7870
:|7870,7871
53AM|7871,7875
BLOOD|7876,7881
Calcium|7882,7889
-|7889,7890
8.6|7890,7893
Phos|7894,7898
-|7898,7899
3.5|7899,7902
Mg|7903,7905
-|7905,7906
2.4|7906,7909
<EOL>|7909,7910
_|7910,7911
_|7911,7912
_|7912,7913
01|7914,7916
:|7916,7917
00PM|7917,7921
BLOOD|7922,7927
calTIBC|7928,7935
-|7935,7936
352|7936,7939
Ferritn|7940,7947
-|7947,7948
111|7948,7951
TRF|7952,7955
-|7955,7956
271|7956,7959
<EOL>|7959,7960
<EOL>|7961,7962
Brief|7962,7967
Hospital|7968,7976
Course|7977,7983
:|7983,7984
<EOL>|7984,7985
TRANSITIONAL|7985,7997
ISSUES|7998,8004
<EOL>|8005,8006
=|8006,8007
=|8007,8008
=|8008,8009
=|8009,8010
=|8010,8011
=|8011,8012
=|8012,8013
=|8013,8014
=|8014,8015
=|8015,8016
=|8016,8017
=|8017,8018
=|8018,8019
=|8019,8020
=|8020,8021
=|8021,8022
=|8022,8023
=|8023,8024
=|8024,8025
=|8025,8026
<EOL>|8027,8028
DISCHARGE|8028,8037
WEIGHT|8038,8044
:|8044,8045
55.6|8046,8050
kg|8051,8053
(|8054,8055
122.57|8055,8061
lb|8062,8064
)|8064,8065
<EOL>|8066,8067
DISCHARGE|8067,8076
Cr|8077,8079
/|8079,8080
BUN|8080,8083
:|8083,8084
Cr|8085,8087
2.2|8088,8091
,|8091,8092
BUN|8093,8096
43|8097,8099
<EOL>|8099,8100
DISCHARGE|8100,8109
DIURETIC|8110,8118
:|8118,8119
40|8120,8122
Torsemide|8123,8132
daily|8133,8138
<EOL>|8138,8139
MEDICATION|8139,8149
CHANGES|8150,8157
:|8157,8158
Decreased|8159,8168
daily|8169,8174
potassium|8175,8184
to|8185,8187
40|8188,8190
mEq|8191,8194
daily|8195,8200
<EOL>|8201,8202
(|8202,8203
from|8203,8207
30|8208,8210
mEq|8211,8214
twice|8215,8220
dailye|8221,8227
)|8227,8228
<EOL>|8228,8229
<EOL>|8229,8230
[|8230,8231
]|8231,8232
Please|8233,8239
obtain|8240,8246
repeat|8247,8253
Chem10|8254,8260
within|8261,8267
2|8268,8269
weeks|8270,8275
and|8276,8279
after|8280,8285
4|8286,8287
weeks|8288,8293
.|8293,8294
<EOL>|8295,8296
Adjust|8296,8302
electrolyte|8303,8314
repletion|8315,8324
accordingly|8325,8336
.|8336,8337
<EOL>|8337,8338
[|8338,8339
]|8339,8340
Please|8341,8347
follow|8348,8354
up|8355,8357
weight|8358,8364
and|8365,8368
volume|8369,8375
status|8376,8382
and|8383,8386
adjust|8387,8393
<EOL>|8394,8395
torsemide|8395,8404
accordingly|8405,8416
.|8416,8417
<EOL>|8418,8419
<EOL>|8419,8420
#|8420,8421
CODE|8421,8425
STATUS|8426,8432
:|8432,8433
Presumed|8434,8442
full|8443,8447
<EOL>|8447,8448
Health|8448,8454
care|8455,8459
proxy|8460,8465
chosen|8466,8472
:|8472,8473
Yes|8474,8477
<EOL>|8478,8479
Name|8479,8483
of|8484,8486
health|8487,8493
care|8494,8498
proxy|8499,8504
:|8504,8505
_|8506,8507
_|8507,8508
_|8508,8509
<EOL>|8510,8511
_|8511,8512
_|8512,8513
_|8513,8514
:|8514,8515
son|8516,8519
<EOL>|8520,8521
Phone|8521,8526
number|8527,8533
:|8533,8534
_|8535,8536
_|8536,8537
_|8537,8538
<EOL>|8539,8540
<EOL>|8540,8541
=|8541,8542
=|8542,8543
=|8543,8544
=|8544,8545
=|8545,8546
=|8546,8547
=|8547,8548
=|8548,8549
=|8549,8550
=|8550,8551
=|8551,8552
=|8552,8553
=|8553,8554
=|8554,8555
=|8555,8556
=|8556,8557
=|8557,8558
=|8558,8559
=|8559,8560
=|8560,8561
<EOL>|8562,8563
PATIENT|8563,8570
SUMMARY|8571,8578
:|8578,8579
<EOL>|8580,8581
=|8581,8582
=|8582,8583
=|8583,8584
=|8584,8585
=|8585,8586
=|8586,8587
=|8587,8588
=|8588,8589
=|8589,8590
=|8590,8591
=|8591,8592
=|8592,8593
=|8593,8594
=|8594,8595
=|8595,8596
=|8596,8597
=|8597,8598
=|8598,8599
=|8599,8600
=|8600,8601
<EOL>|8602,8603
Mr.|8603,8606
_|8607,8608
_|8608,8609
_|8609,8610
is|8611,8613
a|8614,8615
_|8616,8617
_|8617,8618
_|8618,8619
gentleman|8620,8629
with|8630,8634
PMHx|8635,8639
of|8640,8642
CAD|8643,8646
s|8647,8648
/|8648,8649
p|8649,8650
<EOL>|8651,8652
CABG|8652,8656
<EOL>|8656,8657
and|8657,8660
subsequent|8661,8671
PCI|8672,8675
,|8675,8676
HFrEF|8677,8682
(|8683,8684
35|8684,8686
%|8686,8687
_|8688,8689
_|8689,8690
_|8690,8691
,|8691,8692
moderate|8693,8701
tricuspid|8702,8711
<EOL>|8711,8712
regurgitation|8712,8725
,|8725,8726
right|8727,8732
ventricular|8733,8744
dysfunction|8745,8756
,|8756,8757
moderate|8758,8766
pulmonary|8767,8776
<EOL>|8776,8777
hypertension|8777,8789
,|8789,8790
and|8791,8794
paroxysmal|8795,8805
atrial|8806,8812
fibrillation|8813,8825
on|8826,8828
apixaban|8829,8837
,|8837,8838
<EOL>|8838,8839
stage|8839,8844
III|8845,8848
chronic|8849,8856
kidney|8857,8863
disease|8864,8871
(|8872,8873
Baseline|8873,8881
Cr|8882,8884
2.0|8885,8888
-|8888,8889
2.1|8889,8892
)|8892,8893
,|8893,8894
<EOL>|8894,8895
cerebrovascular|8895,8910
disease|8911,8918
,|8918,8919
and|8920,8923
metastatic|8924,8934
melanoma|8935,8943
of|8944,8946
unknown|8947,8954
<EOL>|8954,8955
primary|8955,8962
on|8963,8965
checkpoint|8966,8976
inhibitor|8977,8986
pembrolizumab|8987,9000
who|9001,9004
was|9005,9008
found|9009,9014
<EOL>|9014,9015
volume|9015,9021
overloaded|9022,9032
with|9033,9037
increased|9038,9047
DOE|9048,9051
,|9051,9052
admitted|9053,9061
to|9062,9064
acute|9065,9070
_|9071,9072
_|9072,9073
_|9073,9074
<EOL>|9075,9076
failure|9076,9083
for|9084,9087
IV|9088,9090
diuresis|9091,9099
,|9099,9100
now|9101,9104
transitioned|9105,9117
to|9118,9120
oral|9121,9125
duiretics|9126,9135
.|9135,9136
<EOL>|9137,9138
<EOL>|9138,9139
#|9139,9140
CORONARIES|9141,9151
:|9151,9152
Left|9153,9157
Main|9158,9162
and|9163,9166
two|9167,9170
vessel|9171,9177
coronary|9178,9186
disease|9187,9194
(|9195,9196
_|9196,9197
_|9197,9198
_|9198,9199
)|9199,9200
.|9200,9201
<EOL>|9201,9202
#|9202,9203
PUMP|9204,9208
:|9208,9209
35|9210,9212
%|9212,9213
_|9214,9215
_|9215,9216
_|9216,9217
<EOL>|9218,9219
#|9219,9220
RHYTHM|9221,9227
:|9227,9228
Ectopic|9229,9236
rhythm|9237,9243
,|9243,9244
PR|9245,9247
prolongation|9248,9260
,|9260,9261
left|9262,9266
axis|9267,9271
deviation|9272,9281
,|9281,9282
<EOL>|9283,9284
RBBB|9284,9288
<EOL>|9288,9289
<EOL>|9289,9290
ACTIVE|9290,9296
ISSUES|9297,9303
:|9303,9304
<EOL>|9305,9306
=|9306,9307
=|9307,9308
=|9308,9309
=|9309,9310
=|9310,9311
=|9311,9312
=|9312,9313
=|9313,9314
=|9314,9315
=|9315,9316
=|9316,9317
=|9317,9318
=|9318,9319
=|9319,9320
<EOL>|9321,9322
#|9322,9323
_|9324,9325
_|9325,9326
_|9326,9327
Failure|9328,9335
with|9336,9340
reduced|9341,9348
ejection|9349,9357
fraction|9358,9366
<EOL>|9366,9367
#|9367,9368
Right|9369,9374
ventricular|9375,9386
dysfunction|9387,9398
,|9398,9399
TR|9400,9402
,|9402,9403
pulm|9404,9408
HTN|9409,9412
<EOL>|9412,9413
#|9413,9414
Volume|9415,9421
overload|9422,9430
<EOL>|9430,9431
His|9431,9434
_|9435,9436
_|9436,9437
_|9437,9438
failure|9439,9446
exacerbation|9447,9459
is|9460,9462
likely|9463,9469
secondary|9470,9479
to|9480,9482
his|9483,9486
recent|9487,9493
<EOL>|9493,9494
administration|9494,9508
of|9509,9511
IV|9512,9514
fluids|9515,9521
in|9522,9524
addition|9525,9533
to|9534,9536
his|9537,9540
self|9541,9545
down|9546,9550
<EOL>|9550,9551
titration|9551,9560
of|9561,9563
his|9564,9567
torsemide|9568,9577
over|9578,9582
the|9583,9586
last|9587,9591
week|9592,9596
.|9596,9597
In|9598,9600
addition|9601,9609
,|9609,9610
he|9611,9613
<EOL>|9613,9614
does|9614,9618
not|9619,9622
follow|9623,9629
a|9630,9631
restricted|9632,9642
fluid|9643,9648
intake|9649,9655
and|9656,9659
drinks|9660,9666
_|9667,9668
_|9668,9669
_|9669,9670
glasses|9671,9678
<EOL>|9678,9679
of|9679,9681
water|9682,9687
or|9688,9690
juice|9691,9696
daily|9697,9702
.|9702,9703
Furthermore|9704,9715
,|9715,9716
he|9717,9719
has|9720,9723
not|9724,9727
tolerated|9728,9737
<EOL>|9737,9738
guideline|9738,9747
directed|9748,9756
medical|9757,9764
therapy|9765,9772
due|9773,9776
to|9777,9779
recurrent|9780,9789
issues|9790,9796
with|9797,9801
<EOL>|9801,9802
acute|9802,9807
kidney|9808,9814
injury|9815,9821
and|9822,9825
elevated|9826,9834
transaminitis|9835,9848
while|9849,9854
on|9855,9857
<EOL>|9857,9858
pembrolizumab|9858,9871
therapy|9872,9879
.|9879,9880
He|9881,9883
was|9884,9887
clinically|9888,9898
volume|9899,9905
overloaded|9906,9916
with|9917,9921
<EOL>|9921,9922
elevated|9922,9930
BNP|9931,9934
16020|9935,9940
.|9940,9941
We|9942,9944
initiated|9945,9954
IV|9955,9957
lasix|9958,9963
160|9964,9967
bolus|9968,9973
and|9974,9977
put|9978,9981
him|9982,9985
<EOL>|9986,9987
on|9987,9989
a|9990,9991
lasix|9992,9997
gtt|9998,10001
with|10002,10006
good|10007,10011
response|10012,10020
,|10020,10021
however|10022,10029
he|10030,10032
his|10033,10036
Cr|10037,10039
increased|10040,10049
<EOL>|10050,10051
from|10051,10055
2.1|10056,10059
-|10059,10060
-|10060,10061
>|10061,10062
2.7|10062,10065
.|10065,10066
His|10067,10070
Cr.|10071,10074
improved|10075,10083
with|10084,10088
transition|10089,10099
to|10100,10102
PO|10103,10105
Torsemide|10106,10115
<EOL>|10116,10117
40|10117,10119
mg|10120,10122
daily|10123,10128
.|10128,10129
We|10130,10132
monitored|10133,10142
and|10143,10146
aggressively|10147,10159
repleted|10160,10168
his|10169,10172
<EOL>|10173,10174
potassium|10174,10183
.|10183,10184
No|10185,10187
afterload|10188,10197
reduction|10198,10207
or|10208,10210
neural|10211,10217
hormonal|10218,10226
blockade|10227,10235
<EOL>|10236,10237
was|10237,10240
added|10241,10246
.|10246,10247
<EOL>|10247,10248
<EOL>|10248,10249
#|10249,10250
Chronic|10251,10258
Kidney|10259,10265
Disease|10266,10273
:|10273,10274
Baseline|10275,10283
2.1|10284,10287
-|10287,10288
2.3|10288,10291
.|10292,10293
<EOL>|10294,10295
Cr|10295,10297
2.1|10298,10301
on|10302,10304
admission|10305,10314
(|10314,10315
Stable|10315,10321
)|10322,10323
-|10323,10324
Cr|10325,10327
on|10328,10330
discharge|10331,10340
:|10340,10341
2.2|10341,10344
<EOL>|10344,10345
Cr|10345,10347
initially|10348,10357
uptrended|10358,10367
above|10368,10373
baseline|10374,10382
from|10383,10387
2.1|10388,10391
-|10391,10392
-|10392,10393
-|10393,10394
>|10394,10395
2.7|10396,10399
.|10399,10400
Felt|10401,10405
<EOL>|10406,10407
likely|10407,10413
due|10414,10417
to|10418,10420
increased|10421,10430
diuretic|10431,10439
usage|10440,10445
as|10446,10448
it|10449,10451
improved|10452,10460
with|10461,10465
<EOL>|10466,10467
stopping|10467,10475
diuretics|10476,10485
.|10485,10486
Less|10487,10491
likely|10492,10498
cardiorenal|10499,10510
syndrome|10511,10519
.|10519,10520
In|10521,10523
<EOL>|10524,10525
addition|10525,10533
,|10533,10534
patient|10534,10541
was|10542,10545
recently|10546,10554
seen|10555,10559
in|10560,10562
follow|10563,10569
-|10569,10570
up|10570,10572
by|10573,10575
nephrology|10576,10586
.|10586,10587
<EOL>|10588,10589
They|10589,10593
felt|10594,10598
his|10599,10602
CKD|10603,10606
was|10607,10610
less|10611,10615
likely|10616,10622
to|10623,10625
be|10626,10628
related|10629,10636
to|10637,10639
pembrolizumab|10640,10653
<EOL>|10654,10655
and|10655,10658
more|10659,10663
likely|10664,10670
related|10671,10678
to|10679,10681
age|10682,10685
-|10685,10686
related|10686,10693
decline|10694,10701
in|10702,10704
renal|10705,10710
<EOL>|10711,10712
function|10712,10720
.|10720,10721
Creatinine|10722,10732
2.2|10733,10736
on|10737,10739
discharge|10740,10749
(|10750,10751
stable|10751,10757
)|10757,10758
.|10758,10759
<EOL>|10759,10760
<EOL>|10760,10761
#|10761,10762
Metastatic|10763,10773
Melanoma|10774,10782
<EOL>|10783,10784
He|10784,10786
is|10787,10789
followed|10790,10798
by|10799,10801
Dr.|10802,10805
_|10806,10807
_|10807,10808
_|10808,10809
.|10809,10810
He|10811,10813
was|10814,10817
previously|10818,10828
on|10829,10831
<EOL>|10831,10832
Pembrolizumab|10832,10845
which|10846,10851
was|10852,10855
held|10856,10860
due|10861,10864
diarrhea|10865,10873
,|10873,10874
elevated|10875,10883
LFTs|10884,10888
and|10889,10892
<EOL>|10892,10893
worsening|10893,10902
kidney|10903,10909
function|10910,10918
.|10918,10919
Negative|10920,10928
troponin|10929,10937
and|10938,10941
CK|10942,10944
MB|10945,10947
,|10947,10948
no|10949,10951
<EOL>|10952,10953
concern|10953,10960
<EOL>|10960,10961
for|10961,10964
drug|10965,10969
-|10969,10970
induced|10970,10977
myocarditis|10978,10989
at|10990,10992
this|10993,10997
point|10998,11003
.|11003,11004
Followup|11005,11013
in|11014,11016
<EOL>|11017,11018
_|11018,11019
_|11019,11020
_|11020,11021
clinic|11022,11028
in|11029,11031
2weeks|11032,11038
after|11039,11044
discharge|11045,11054
<EOL>|11054,11055
<EOL>|11055,11056
#|11056,11057
Elevated|11058,11066
transaminiatis|11067,11081
<EOL>|11081,11082
Stable|11082,11088
.|11088,11089
Statin|11090,11096
and|11097,11100
_|11101,11102
_|11102,11103
_|11103,11104
had|11105,11108
previously|11109,11119
been|11120,11124
held|11125,11129
.|11129,11130
No|11131,11133
changes|11134,11141
made|11142,11146
<EOL>|11147,11148
during|11148,11154
admission|11155,11164
.|11164,11165
<EOL>|11166,11167
<EOL>|11167,11168
#|11168,11169
Urinary|11170,11177
frequency|11178,11187
<EOL>|11187,11188
Likely|11188,11194
due|11195,11198
to|11199,11201
diuretic|11202,11210
use|11211,11214
.|11214,11215
Afebrile|11216,11224
and|11225,11228
asx|11229,11232
otherwise|11233,11242
<EOL>|11242,11243
-|11243,11244
Continued|11244,11253
home|11254,11258
tamsulosin|11259,11269
<EOL>|11269,11270
<EOL>|11270,11271
#|11271,11272
Coronary|11273,11281
artery|11282,11288
disease|11289,11296
,|11296,11297
s|11298,11299
/|11299,11300
p|11300,11301
CABG|11302,11306
and|11307,11310
LAD|11311,11314
PCI|11315,11318
.|11318,11319
<EOL>|11319,11320
-|11320,11321
Continued|11321,11330
aspirin|11331,11338
81|11339,11341
mg|11342,11344
daily|11345,11350
<EOL>|11350,11351
-|11351,11352
Statin|11352,11358
stopped|11359,11366
prior|11367,11372
to|11373,11375
admission|11376,11385
due|11386,11389
to|11390,11392
elevated|11393,11401
LFTs|11402,11406
.|11406,11407
<EOL>|11408,11409
Continued|11409,11418
holding|11419,11426
.|11426,11427
<EOL>|11428,11429
<EOL>|11429,11430
CHRONIC|11430,11437
ISSUES|11438,11444
:|11444,11445
<EOL>|11446,11447
=|11447,11448
=|11448,11449
=|11449,11450
=|11450,11451
=|11451,11452
=|11452,11453
=|11453,11454
=|11454,11455
=|11455,11456
=|11456,11457
=|11457,11458
=|11458,11459
=|11459,11460
=|11460,11461
<EOL>|11462,11463
<EOL>|11463,11464
#|11464,11465
Paroxysmal|11466,11476
Atrial|11477,11483
fibrillation|11484,11496
<EOL>|11496,11497
Rythym|11497,11503
:|11503,11504
Continue|11505,11513
amiodarone|11514,11524
200mg|11525,11530
for|11531,11534
rhythm|11535,11541
control|11542,11549
strategy|11550,11558
<EOL>|11558,11559
(|11559,11560
monitoring|11560,11570
safety|11571,11577
labs|11578,11582
)|11582,11583
<EOL>|11583,11584
-|11584,11585
Continued|11585,11594
anticoagulation|11595,11610
with|11611,11615
apixaban|11616,11624
2.5|11625,11628
mg|11628,11630
twice|11631,11636
daily|11637,11642
<EOL>|11642,11643
<EOL>|11643,11644
#|11644,11645
Hypertension|11646,11658
:|11658,11659
Stable|11660,11666
.|11666,11667
<EOL>|11668,11669
<EOL>|11670,11671
Medications|11671,11682
on|11683,11685
Admission|11686,11695
:|11695,11696
<EOL>|11696,11697
The|11697,11700
Preadmission|11701,11713
Medication|11714,11724
list|11725,11729
may|11730,11733
be|11734,11736
inaccurate|11737,11747
and|11748,11751
requires|11752,11760
<EOL>|11761,11762
further|11762,11769
investigation|11770,11783
.|11783,11784
<EOL>|11784,11785
1.|11785,11787
Amiodarone|11788,11798
200|11799,11802
mg|11803,11805
PO|11806,11808
DAILY|11809,11814
<EOL>|11815,11816
2.|11816,11818
Aspirin|11819,11826
81|11827,11829
mg|11830,11832
PO|11833,11835
DAILY|11836,11841
<EOL>|11842,11843
3.|11843,11845
Docusate|11846,11854
Sodium|11855,11861
100|11862,11865
mg|11866,11868
PO|11869,11871
BID|11872,11875
<EOL>|11876,11877
4.|11877,11879
Senna|11880,11885
17.2|11886,11890
mg|11891,11893
PO|11894,11896
HS|11897,11899
<EOL>|11900,11901
5.|11901,11903
Vitamin|11904,11911
D|11912,11913
1000|11914,11918
UNIT|11919,11923
PO|11924,11926
DAILY|11927,11932
<EOL>|11933,11934
6.|11934,11936
Align|11937,11942
(|11943,11944
bifidobacterium|11944,11959
infantis|11960,11968
)|11968,11969
4|11970,11971
mg|11972,11974
oral|11975,11979
DAILY|11980,11985
<EOL>|11986,11987
7.|11987,11989
coenzyme|11990,11998
Q10|11999,12002
100|12003,12006
mg|12007,12009
oral|12010,12014
DAILY|12015,12020
<EOL>|12021,12022
8.|12022,12024
Tamsulosin|12025,12035
0.4|12036,12039
mg|12040,12042
PO|12043,12045
QHS|12046,12049
<EOL>|12050,12051
9.|12051,12053
Torsemide|12054,12063
40|12064,12066
mg|12067,12069
PO|12070,12072
DAILY|12073,12078
<EOL>|12079,12080
10.|12080,12083
Ferrous|12084,12091
Sulfate|12092,12099
325|12100,12103
mg|12104,12106
PO|12107,12109
DAILY|12110,12115
<EOL>|12116,12117
11.|12117,12120
Sertraline|12121,12131
50|12132,12134
mg|12135,12137
PO|12138,12140
DAILY|12141,12146
<EOL>|12147,12148
12.|12148,12151
Potassium|12152,12161
Chloride|12162,12170
30|12171,12173
mEq|12174,12177
PO|12178,12180
BID|12181,12184
<EOL>|12185,12186
13.|12186,12189
Apixaban|12190,12198
2.5|12199,12202
mg|12203,12205
PO|12206,12208
BID|12209,12212
<EOL>|12213,12214
14.|12214,12217
Cephalexin|12218,12228
500|12229,12232
mg|12233,12235
PO|12236,12238
Q6H|12239,12242
<EOL>|12243,12244
<EOL>|12244,12245
<EOL>|12246,12247
Discharge|12247,12256
Medications|12257,12268
:|12268,12269
<EOL>|12269,12270
1.|12270,12272
Potassium|12274,12283
Chloride|12284,12292
40|12293,12295
mEq|12296,12299
PO|12300,12302
DAILY|12303,12308
<EOL>|12309,12310
RX|12310,12312
*|12313,12314
potassium|12314,12323
chloride|12324,12332
20|12333,12335
mEq|12336,12339
2|12340,12341
packet|12342,12348
(|12348,12349
s|12349,12350
)|12350,12351
by|12352,12354
mouth|12355,12360
once|12361,12365
a|12366,12367
day|12368,12371
<EOL>|12372,12373
Disp|12373,12377
#|12378,12379
*|12379,12380
60|12380,12382
Tablet|12383,12389
Refills|12390,12397
:|12397,12398
*|12398,12399
0|12399,12400
<EOL>|12401,12402
2.|12402,12404
Align|12406,12411
(|12412,12413
bifidobacterium|12413,12428
infantis|12429,12437
)|12437,12438
4|12439,12440
mg|12441,12443
oral|12444,12448
DAILY|12449,12454
<EOL>|12456,12457
3.|12457,12459
Amiodarone|12461,12471
200|12472,12475
mg|12476,12478
PO|12479,12481
DAILY|12482,12487
<EOL>|12489,12490
4.|12490,12492
Apixaban|12494,12502
2.5|12503,12506
mg|12507,12509
PO|12510,12512
BID|12513,12516
<EOL>|12518,12519
5.|12519,12521
Aspirin|12523,12530
81|12531,12533
mg|12534,12536
PO|12537,12539
DAILY|12540,12545
<EOL>|12547,12548
6.|12548,12550
coenzyme|12552,12560
Q10|12561,12564
100|12565,12568
mg|12569,12571
oral|12572,12576
DAILY|12577,12582
<EOL>|12584,12585
7.|12585,12587
Docusate|12589,12597
Sodium|12598,12604
100|12605,12608
mg|12609,12611
PO|12612,12614
BID|12615,12618
<EOL>|12620,12621
8.|12621,12623
Ferrous|12625,12632
Sulfate|12633,12640
325|12641,12644
mg|12645,12647
PO|12648,12650
DAILY|12651,12656
<EOL>|12658,12659
9.|12659,12661
Senna|12663,12668
17.2|12669,12673
mg|12674,12676
PO|12677,12679
HS|12680,12682
<EOL>|12684,12685
10.|12685,12688
Sertraline|12690,12700
50|12701,12703
mg|12704,12706
PO|12707,12709
DAILY|12710,12715
<EOL>|12717,12718
11.|12718,12721
Tamsulosin|12723,12733
0.4|12734,12737
mg|12738,12740
PO|12741,12743
QHS|12744,12747
<EOL>|12748,12749
RX|12749,12751
*|12752,12753
tamsulosin|12753,12763
0.4|12764,12767
mg|12768,12770
1|12771,12772
capsule|12773,12780
(|12780,12781
s|12781,12782
)|12782,12783
by|12784,12786
mouth|12787,12792
nightly|12793,12800
Disp|12801,12805
#|12806,12807
*|12807,12808
30|12808,12810
<EOL>|12811,12812
Capsule|12812,12819
Refills|12820,12827
:|12827,12828
*|12828,12829
0|12829,12830
<EOL>|12831,12832
12.|12832,12835
Torsemide|12837,12846
40|12847,12849
mg|12850,12852
PO|12853,12855
DAILY|12856,12861
<EOL>|12863,12864
13|12864,12866
.|12866,12867
Vitamin|12869,12876
D|12877,12878
1000|12879,12883
UNIT|12884,12888
PO|12889,12891
DAILY|12892,12897
<EOL>|12899,12900
<EOL>|12900,12901
<EOL>|12902,12903
Discharge|12903,12912
Disposition|12913,12924
:|12924,12925
<EOL>|12925,12926
Home|12926,12930
With|12931,12935
Service|12936,12943
<EOL>|12943,12944
<EOL>|12945,12946
Facility|12946,12954
:|12954,12955
<EOL>|12955,12956
_|12956,12957
_|12957,12958
_|12958,12959
<EOL>|12959,12960
<EOL>|12961,12962
Discharge|12962,12971
Diagnosis|12972,12981
:|12981,12982
<EOL>|12982,12983
Primary|12983,12990
Diagnosis|12991,13000
<EOL>|13000,13001
=|13001,13002
=|13002,13003
=|13003,13004
=|13004,13005
=|13005,13006
=|13006,13007
=|13007,13008
=|13008,13009
=|13009,13010
=|13010,13011
=|13011,13012
=|13012,13013
=|13013,13014
=|13014,13015
=|13015,13016
=|13016,13017
=|13017,13018
<EOL>|13018,13019
HFrEF|13019,13024
excerterbation|13025,13039
<EOL>|13039,13040
<EOL>|13040,13041
Secondary|13041,13050
diagnosis|13051,13060
<EOL>|13060,13061
=|13061,13062
=|13062,13063
=|13063,13064
=|13064,13065
=|13065,13066
=|13066,13067
=|13067,13068
=|13068,13069
=|13069,13070
=|13070,13071
=|13071,13072
=|13072,13073
=|13073,13074
=|13074,13075
=|13075,13076
=|13076,13077
=|13077,13078
=|13078,13079
=|13079,13080
<EOL>|13080,13081
Transaminitis|13081,13094
<EOL>|13094,13095
Metastatic|13095,13105
melanoma|13106,13114
<EOL>|13114,13115
CKD|13115,13118
<EOL>|13118,13119
Coronary|13119,13127
artery|13128,13134
disease|13135,13142
,|13142,13143
s|13144,13145
/|13145,13146
p|13146,13147
CABG|13148,13152
and|13153,13156
LAD|13157,13160
PCI|13161,13164
<EOL>|13164,13165
<EOL>|13165,13166
<EOL>|13167,13168
Discharge|13168,13177
Condition|13178,13187
:|13187,13188
<EOL>|13188,13189
Mental|13189,13195
Status|13196,13202
:|13202,13203
Clear|13204,13209
and|13210,13213
coherent|13214,13222
.|13222,13223
<EOL>|13223,13224
Level|13224,13229
of|13230,13232
Consciousness|13233,13246
:|13246,13247
Alert|13248,13253
and|13254,13257
interactive|13258,13269
.|13269,13270
<EOL>|13270,13271
Activity|13271,13279
Status|13280,13286
:|13286,13287
Ambulatory|13288,13298
-|13299,13300
requires|13301,13309
assistance|13310,13320
or|13321,13323
aid|13324,13327
(|13328,13329
walker|13329,13335
<EOL>|13336,13337
or|13337,13339
cane|13340,13344
)|13344,13345
.|13345,13346
<EOL>|13346,13347
<EOL>|13347,13348
<EOL>|13349,13350
Discharge|13350,13359
Instructions|13360,13372
:|13372,13373
<EOL>|13373,13374
=|13374,13375
=|13375,13376
=|13376,13377
=|13377,13378
=|13378,13379
=|13379,13380
=|13380,13381
=|13381,13382
=|13382,13383
=|13383,13384
=|13384,13385
=|13385,13386
=|13386,13387
=|13387,13388
=|13388,13389
=|13389,13390
=|13390,13391
=|13391,13392
=|13392,13393
=|13393,13394
=|13394,13395
=|13395,13396
=|13396,13397
=|13397,13398
=|13398,13399
<EOL>|13401,13402
DISCHARGE|13402,13411
INSTRUCTIONS|13412,13424
<EOL>|13426,13427
=|13427,13428
=|13428,13429
=|13429,13430
=|13430,13431
=|13431,13432
=|13432,13433
=|13433,13434
=|13434,13435
=|13435,13436
=|13436,13437
=|13437,13438
=|13438,13439
=|13439,13440
=|13440,13441
=|13441,13442
=|13442,13443
=|13443,13444
=|13444,13445
=|13445,13446
=|13446,13447
=|13447,13448
=|13448,13449
=|13449,13450
=|13450,13451
=|13451,13452
=|13452,13453
<EOL>|13455,13456
<EOL>|13456,13457
Dear|13457,13461
Mr.|13462,13465
_|13466,13467
_|13467,13468
_|13468,13469
,|13470,13471
<EOL>|13473,13474
<EOL>|13474,13475
It|13475,13477
was|13478,13481
a|13482,13483
pleasure|13484,13492
taking|13493,13499
care|13500,13504
of|13505,13507
you|13508,13511
at|13512,13514
_|13515,13516
_|13516,13517
_|13517,13518
<EOL>|13519,13520
_|13520,13521
_|13521,13522
_|13522,13523
.|13523,13524
<EOL>|13525,13526
<EOL>|13527,13528
WHY|13528,13531
WAS|13532,13535
I|13536,13537
ADMITTED|13538,13546
TO|13547,13549
THE|13550,13553
HOSPITAL|13554,13562
?|13562,13563
<EOL>|13565,13566
You|13566,13569
were|13570,13574
feeling|13575,13582
short|13583,13588
of|13589,13591
breath|13592,13598
because|13599,13606
you|13607,13610
had|13611,13614
fluid|13615,13620
in|13621,13623
your|13624,13628
<EOL>|13629,13630
lungs|13630,13635
.|13635,13636
This|13637,13641
was|13642,13645
caused|13646,13652
by|13653,13655
a|13656,13657
condition|13658,13667
called|13668,13674
_|13675,13676
_|13676,13677
_|13677,13678
failure|13679,13686
,|13686,13687
<EOL>|13688,13689
where|13689,13694
your|13695,13699
_|13700,13701
_|13701,13702
_|13702,13703
does|13704,13708
not|13709,13712
pump|13713,13717
hard|13718,13722
enough|13723,13729
and|13730,13733
fluid|13734,13739
backs|13740,13745
up|13746,13748
<EOL>|13749,13750
into|13750,13754
your|13755,13759
lungs|13760,13765
.|13765,13766
<EOL>|13768,13769
<EOL>|13769,13770
WHAT|13770,13774
HAPPENED|13775,13783
WHILE|13784,13789
I|13790,13791
WAS|13792,13795
IN|13796,13798
THE|13799,13802
HOSPITAL|13803,13811
?|13811,13812
<EOL>|13814,13815
You|13815,13818
were|13819,13823
given|13824,13829
medications|13830,13841
to|13842,13844
help|13845,13849
get|13850,13853
the|13854,13857
fluid|13858,13863
out|13864,13867
.|13867,13868
Your|13869,13873
<EOL>|13874,13875
breathing|13875,13884
got|13885,13888
better|13889,13895
and|13896,13899
were|13900,13904
ready|13905,13910
to|13911,13913
leave|13914,13919
the|13920,13923
hospital|13924,13932
.|13932,13933
<EOL>|13935,13936
<EOL>|13936,13937
WHAT|13937,13941
DO|13942,13944
YOU|13945,13948
NEED|13949,13953
TO|13954,13956
DO|13957,13959
WHEN|13960,13964
YOU|13965,13968
LEAVE|13969,13974
THE|13975,13978
HOSPITAL|13979,13987
?|13987,13988
<EOL>|13990,13991
-|13991,13992
Take|13993,13997
all|13998,14001
of|14002,14004
your|14005,14009
medications|14010,14021
as|14022,14024
prescribed|14025,14035
(|14036,14037
listed|14037,14043
below|14044,14049
)|14049,14050
<EOL>|14052,14053
-|14053,14054
Follow|14055,14061
up|14062,14064
with|14065,14069
your|14070,14074
doctors|14075,14082
as|14083,14085
listed|14086,14092
below|14093,14098
<EOL>|14100,14101
-|14101,14102
Weigh|14103,14108
yourself|14109,14117
every|14118,14123
morning|14124,14131
.|14131,14132
Your|14133,14137
weight|14138,14144
on|14145,14147
discharge|14148,14157
is|14158,14160
<EOL>|14161,14162
122.57|14162,14168
lbs|14169,14172
.|14172,14173
Call|14174,14178
your|14179,14183
doctor|14184,14190
if|14191,14193
your|14194,14198
weight|14199,14205
goes|14206,14210
up|14211,14213
more|14214,14218
than|14219,14223
3|14224,14225
<EOL>|14226,14227
pounds|14227,14233
.|14233,14234
<EOL>|14234,14235
-|14235,14236
Call|14237,14241
you|14242,14245
doctor|14246,14252
if|14253,14255
you|14256,14259
notice|14260,14266
any|14267,14270
of|14271,14273
the|14274,14277
"|14278,14279
danger|14279,14285
signs|14286,14291
"|14291,14292
below|14293,14298
.|14298,14299
<EOL>|14300,14301
<EOL>|14302,14303
<EOL>|14304,14305
We|14305,14307
wish|14308,14312
you|14313,14316
the|14317,14320
best|14321,14325
!|14325,14326
<EOL>|14328,14329
Your|14329,14333
_|14334,14335
_|14335,14336
_|14336,14337
Care|14338,14342
Team|14343,14347
<EOL>|14349,14350
<EOL>|14350,14351
<EOL>|14352,14353
Followup|14353,14361
Instructions|14362,14374
:|14374,14375
<EOL>|14375,14376
_|14376,14377
_|14377,14378
_|14378,14379
<EOL>|14379,14380

