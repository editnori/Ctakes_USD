CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|localized swelling in left breast|Finding|false|false|C0006141;C0222601|left breast swellingnull|Left breast|Anatomy|false|false|C1552822;C1549543;C0030193;C0496956;C0567499;C0006152;C0013604;C0038999;C0191838;C2127345|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0222601;C0006141|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swelling of breast|Finding|false|false|C0006141;C0222601|breast swellingnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0222601;C0006141|breastnull|Breast problem|Finding|false|false|C0006141;C0222601|breastnull|Procedures on breast|Procedure|false|false|C0006141;C0222601|breastnull|Breast|Anatomy|false|false|C0567499;C1552822;C0496956;C0006152;C2127345;C0013604;C0038999;C0191838|breastnull|Swelling|Finding|false|false|C0006141;C0222601|swelling
null|Edema|Finding|false|false|C0006141;C0222601|swellingnull|Administration Method - Pain|Finding|false|false|C0222601|pain
null|Pain|Finding|false|false|C0222601|painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Evacuation of hematoma|Procedure|false|false||Evacuation of hematomanull|Evacuation procedure|Procedure|false|false||Evacuationnull|Hematoma|Finding|false|false||hematomanull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0191838;C1881349;C1449563;C0496956;C0567499|breastnull|Cardiomyopathy, Familial Idiopathic|Disorder|false|false|C0006141|IDCnull|LMNA wt Allele|Finding|false|false|C0006141|IDCnull|grade 3 education level|Finding|false|false||Grade 3
null|Tumor grade G3|Finding|false|false||Grade 3
null|Grade three rank|Finding|false|false||Grade 3
null|Simpson Grade 3|Finding|false|false||Grade 3null|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Lumpectomy of breast|Procedure|false|false|C0006141|breast lumpectomynull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0496956;C0191838;C0567499;C0851238;C0796693|breastnull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Sentinel Lymph Node Biopsy|Procedure|false|false|C0006141|SLNBnull|localized swelling in left breast|Finding|false|false|C0006141;C0222601|left breast swellingnull|Left breast|Anatomy|false|false|C0191838;C0496956;C1552822;C2127345;C0006152;C0567499;C0013604;C0038999|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0222601|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swelling of breast|Finding|false|false|C0006141;C0222601|breast swellingnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141;C0222601|breastnull|Breast problem|Finding|false|false|C0222601;C0006141|breastnull|Procedures on breast|Procedure|false|false|C0222601;C0006141|breastnull|Breast|Anatomy|false|false|C0006152;C2127345;C0496956;C0191838;C0567499|breastnull|Swelling|Finding|false|false|C0222601|swelling
null|Edema|Finding|false|false|C0222601|swellingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hematoma|Finding|false|false||hematomanull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false|C0042449|varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0398102;C0042345|veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEs
null|PES1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false|C1418467;C0687136;C4551530|PEs
null|Hindfoot of quadruped|Anatomy|false|false|C1418467;C0687136;C4551530|PEs
null|Paw|Anatomy|false|false|C1418467;C0687136;C4551530|PEs
null|Foot|Anatomy|false|false|C1418467;C0687136;C4551530|PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false|C1167408;C3665580|antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false|C1167408;C3665580|antiphospholipid antibodynull|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibodynull|Antibody (immunoassay)|Procedure|false|false|C1690938;C3853547;C0687080;C0016504;C1167408;C3665580|antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false|C0085278;C4019436;C0003241;C0021027;C4551530;C0162595;C0039082|antibody
null|immunoglobulin complex location|Anatomy|false|false|C0085278;C4019436;C0003241;C0021027;C4551530;C0162595;C0039082|antibodynull|Syndrome|Disorder|false|false|C1167408;C3665580|syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false|C0228174;C0006104|A1Cnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0474680|cerebral
null|Brain|Anatomy|false|false|C0474680|cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|true|false|C0009368;C4071907|colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|true|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|true|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|true|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0032584;C0009376|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0032584;C0009376|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|polyps|Disorder|false|false|C0009368;C4071907|polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false|C3890599|CMC
null|Capillary malformation (disorder)|Disorder|false|false|C3890599|CMCnull|MCC protocol|Procedure|false|false|C3890599|CMCnull|Circulating Melanoma Cell|Anatomy|false|false|C0006845;C0340803;C0065772|CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false|C0392905;C1269611;C0022417|joint arthroplastynull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417|jointnull|null|Anatomy|false|false|C0575044;C5887062;C0003893;C0700235;C0003893|joint
null|Joints|Anatomy|false|false|C0575044;C5887062;C0003893;C0700235;C0003893|joint
null|Articular system|Anatomy|false|false|C0575044;C5887062;C0003893;C0700235;C0003893|jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false|C0392905;C1269611;C0022417|arthroplasty
null|Arthroplasty|Procedure|false|false|C0392905;C1269611;C0022417|arthroplasty
null|Reconstruction of joint|Procedure|false|false|C0392905;C1269611;C0022417|arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false|C0085515;C1550244|rotator cuff repairnull|Rotator Cuff|Anatomy|false|false|C0043240;C4319951;C0015252;C0728940;C0374711;C1705181;C0186666;C3668885|rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false|C1550244;C0085515|cuffnull|Cuff - body part|Anatomy|false|false|C3668885;C0186666|cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false|C0085515|repair
null|Wound Healing|Finding|false|false|C0085515|repairnull|Repair - Remedial Action|Procedure|false|false|C0085515|repair
null|Surgical repair|Procedure|false|false|C0085515|repairnull|Excision|Procedure|false|false|C0085515|excision
null|removal technique|Procedure|false|false|C0085515|excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false|C0582802|digitnull|Digit structure|Anatomy|false|false|C4761764;C4283905;C1546709;C2700045;C0577573;C0577559;C1414542|digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false|C0582802|mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false|C0582802|mass
null|null|Finding|false|false|C0582802|mass
null|FBN1 wt Allele|Finding|false|false|C0582802|mass
null|FBN1 gene|Finding|false|false|C0582802|mass
null|Mass of body region|Finding|false|false|C0582802|massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false|C4482304;C0030288;C0030274;C0687028;C1550227|pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic duct
null|Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic ductnull|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreaticnull|Pancreas|Anatomy|false|false|C0153461;C0030292|pancreaticnull|Duct (organ) structure|Anatomy|false|false|C0153461|duct
null|canal [body parts]|Anatomy|false|false|C0153461|ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false|C4482304;C0030288|explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Entity Name Part Type - family|Finding|false|false|C5239664|family
null|Last Name|Finding|false|false|C5239664|family
null|Living Arrangement - Family|Finding|false|false|C5239664|family
null|Family (taxonomic)|Finding|false|false|C5239664|family
null|Family Collection|Finding|false|false|C5239664|familynull|Family|Subject|false|false||familynull|Deep thrombophlebitis|Disorder|true|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|true|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2700055;C1546847;C1704727;C1301584;C1563343;C2926618|DVTnull|null|Attribute|true|false|C5239664|DVTnull|Sister|Subject|false|false||sistersnull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0344434;C2926591;C0232197;C0004238|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Pleasant|Finding|false|false||pleasantnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|scleranull|examination of sclera|Procedure|false|false|C0036410|scleranull|Sclera|Anatomy|false|false|C2228481;C0036412;C0205180|scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|Increased work of breathing|Finding|true|false||increased work of breathingnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Work of Breathing|Finding|true|false||work of breathingnull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Feeling comfortable|Finding|false|false||comfortablenull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|BREASTnull|Breast problem|Finding|false|false|C0006141|BREASTnull|Procedures on breast|Procedure|false|false|C0006141|BREASTnull|Breast|Anatomy|false|false|C0496956;C0191838;C0567499|BREASTnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C3244310;C0567499;C0496956;C3812660;C0013491;C0191838|breastnull|dependent|Finding|false|false|C0006141|dependentnull|Dependent - ability|Modifier|false|false||dependent
null|Conditional|Modifier|false|false||dependentnull|Ecchymosis|Finding|false|false|C0006141|ecchymosis
null|Skin Bruise|Finding|false|false|C0006141|ecchymosisnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0332803;C0184898;C0496956;C0567499;C0191838|breastnull|Surgical wound|Disorder|false|false|C0006141;C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258;C0006141|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Serosanguineous|Modifier|false|false||serosanguineousnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Hernia|Disorder|true|false||hernianull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Focal Neurologic Deficits|Finding|true|false||focal neurologic deficitsnull|Focal|Modifier|false|false||focalnull|Neurologic Deficits|Finding|true|false||neurologic deficitsnull|Neurologic (qualifier value)|Modifier|false|false||neurologicnull|Deficit|Modifier|false|false||deficitsnull|Psychiatric problem|Disorder|false|false||PSYCH
null|Mental disorders|Disorder|false|false||PSYCHnull|Judgment|Finding|false|false||judgmentnull|Insight|Finding|false|false||insightnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Mood (psychological function)|Finding|false|false||mood
null|mood (physical finding)|Finding|false|false||mood
null|Mood (attribute)|Finding|false|false||moodnull|null|Attribute|false|false||moodnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|Cancer/Testis Antigen|Drug|false|false|C1527391;C0817096|CTAnull|PCYT1A wt Allele|Finding|false|false|C1527391;C0817096|CTA
null|CERNA3 gene|Finding|false|false|C1527391;C0817096|CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false|C1527391;C0817096|CTAnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0741025;C3272310;C3540513;C4554671;C3813556|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0741025;C3272310;C3540513;C4554671;C3813556|CHESTnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Comparison|Event|false|false||COMPARISONnull|Chest CT|Procedure|false|false|C1527391;C0817096|Chest CTnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0202823;C0741025|Chest
null|Anterior thoracic region|Anatomy|false|false|C0202823;C0741025|Chestnull|Malignant neoplasm of heart|Disorder|false|false|C3714653;C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C3714653;C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|HEART
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|HEARTnull|Vasculature|Anatomy|false|false|C0153957;C0153500|VASCULATUREnull|Blood supply aspects|Modifier|false|false||VASCULATUREnull|Central brand of multivitamin with minerals|Drug|true|false||central
null|Central brand of multivitamin with minerals|Drug|true|false||centralnull|Central Minus|Procedure|true|false||centralnull|Central|Modifier|false|false||centralnull|Pulmonary Embolism|Finding|true|false|C0024109|pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268;C0034065;C1704212;C0013922|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|true|false|C0024109|embolism
null|Embolus|Finding|true|false|C0024109|embolismnull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false|C0817096|thoracicnull|Chest|Anatomy|false|false|C5779551|thoracicnull|Procedure on aorta|Procedure|false|false|C4037978;C0003483|aortanull|Chest+Abdomen>Aorta|Anatomy|false|false|C0333288;C3887511;C0869784;C0332120|aorta
null|Aorta|Anatomy|false|false|C0333288;C3887511;C0869784;C0332120|aortanull|Diameter (qualifier value)|LabModifier|false|false||calibernull|Evidence of (contextual qualifier)|Finding|true|false|C4037978;C0003483|evidence ofnull|Evidence|Finding|true|false|C4037978;C0003483|evidencenull|Dissecting hemorrhage|Finding|true|false|C4037978;C0003483|dissectionnull|Tissue Dissection|Procedure|true|false||dissectionnull|Internal|Modifier|false|false||intramuralnull|Hematoma|Finding|false|false||hematomanull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787;C0225991|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787;C0225991|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C1424898;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C1424898;C0795691|heartnull|Pericardial sac structure|Anatomy|false|false||pericardiumnull|Structure of great blood vessel (organ)|Anatomy|false|false|C1424898;C0153957;C0153500|great vesselsnull|RXFP2 gene|Finding|false|false|C0225991;C4037974;C0018787;C0005847|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Blood Vessel|Anatomy|false|false|C1424898|vesselsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Pericardial effusion|Disorder|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial effusion body substance|Finding|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardial
null|Pericardial sac structure|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardialnull|Effusion (substance)|Finding|true|false|C0031050;C0442031|effusion
null|null|Finding|true|false|C0031050;C0442031|effusion
null|effusion|Finding|true|false|C0031050;C0442031|effusionnull|Axilla|Anatomy|false|false|C0153956;C0496915|AXILLAnull|Neoplasm of uncertain or unknown behavior of mediastinum|Disorder|false|false|C0004454;C0025066;C4037971|MEDIASTINUM
null|Benign tumor of mediastinum|Disorder|false|false|C0004454;C0025066;C4037971|MEDIASTINUMnull|Chest>Mediastinum|Anatomy|false|false|C0153956;C0496915|MEDIASTINUM
null|Mediastinum|Anatomy|false|false|C0153956;C0496915|MEDIASTINUMnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Left breast|Anatomy|false|false|C0496956;C0567499;C1552822;C0191838|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0006141;C0222601|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0222601;C0006141|breastnull|Breast problem|Finding|false|false|C0006141;C0222601|breastnull|Procedures on breast|Procedure|false|false|C0006141;C0222601|breastnull|Breast|Anatomy|false|false|C1552822;C0567499;C0496956;C0191838|breastnull|density|LabModifier|false|false||densitynull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Hematoma|Finding|false|false||hematomanull|Focal|Modifier|false|false||foci ofnull|Foci|Finding|false|false||focinull|Focal|Modifier|false|false||focinull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|null|Time|false|false||priornull|Respiratory Aspiration|Disorder|false|false||aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Punctate|Modifier|false|false||punctatenull|Axilla|Anatomy|false|false||axillarynull|Mediastinum|Anatomy|false|false|C0497156;C4282165|mediastinalnull|Mediastinal|Modifier|false|false||mediastinalnull|Hilar lymphadenopathy|Disorder|false|false||hilar lymphadenopathynull|Hilar|Modifier|false|false||hilarnull|Lymphadenopathy|Disorder|false|false|C0025066|lymphadenopathynull|Swollen Lymph Node|Finding|false|false|C0025066|lymphadenopathynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Structure of right axillary region|Anatomy|false|false|C1552823|right axillanull|Table Cell Horizontal Align - right|Finding|false|false|C0004454;C0230337|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Axilla|Anatomy|false|false|C1552823|axillanull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Mediastinal mass|Finding|true|false|C0025066|mediastinal massnull|Mediastinum|Anatomy|false|false|C4283905;C1546709;C2700045;C0577573;C0577559;C1414542;C0240318|mediastinalnull|Mediastinal|Modifier|false|false||mediastinalnull|Mass of body structure|Finding|true|false|C0025066|mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false|C0025066|mass
null|null|Finding|true|false|C0025066|mass
null|FBN1 wt Allele|Finding|true|false|C0025066|mass
null|FBN1 gene|Finding|true|false|C0025066|mass
null|Mass of body region|Finding|true|false|C0025066|massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Pleural cavity|Anatomy|false|false|C0032226|PLEURAL SPACESnull|Pleural Diseases|Disorder|false|false|C0032225;C0178802|PLEURALnull|Pleura|Anatomy|false|false|C0032226|PLEURALnull|Pleural|Modifier|false|false||PLEURALnull|Pleural effusion (disorder)|Finding|true|false|C0032225|pleural effusion
null|Pleural effusion fluid|Finding|true|false|C0032225|pleural effusion
null|null|Finding|true|false|C0032225|pleural effusionnull|Pleural Diseases|Disorder|true|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C2073625;C1253943;C0032227;C0032226;C2317432;C1546613;C0013687|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|true|false|C0032225|effusion
null|null|Finding|true|false|C0032225|effusion
null|effusion|Finding|true|false|C0032225|effusionnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Lung|Anatomy|false|false||LUNGSnull|Airway structure|Anatomy|false|false||AIRWAYSnull|Artificial Airways|Device|false|false||AIRWAYSnull|Lung|Anatomy|false|false|C1550016|lungsnull|Remote control command - Clear|Finding|false|false|C0024109|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Areas <Spilosomini>|Entity|false|false||areasnull|Area|Modifier|false|false||areasnull|Opacification|Modifier|false|false||opacificationnull|Airway structure|Anatomy|false|false|C0030650|airwaysnull|Artificial Airways|Device|false|false||airwaysnull|Legal patent|Finding|false|false|C0458827|patentnull|Open|Modifier|false|false||patentnull|Segmental|Modifier|false|false||segmentalnull|Bronchi|Anatomy|false|false||bronchinull|Base of neck|Anatomy|false|false|C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279;C0812434;C0684335|BASE OF NECKnull|nitrogenous base|Drug|false|false|C3686666;C2987514|BASE
null|Base|Drug|false|false|C3686666;C2987514|BASE
null|Dental Base|Drug|false|false|C3686666;C2987514|BASE
null|base - RoleClass|Drug|false|false|C3686666;C2987514|BASEnull|Base - General Qualifier|Finding|false|false|C3686666;C0027530;C3159206;C2987514|BASE
null|BPIFA4P gene|Finding|false|false|C3686666;C0027530;C3159206;C2987514|BASE
null|Base - RX Component Type|Finding|false|false|C3686666;C0027530;C3159206;C2987514|BASEnull|Anatomical base|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C1549548;C1705938;C1843354;C0812434;C0684335|BASEnull|Base - unit of product usage|LabModifier|false|false||BASEnull|Passive joint movement of neck (finding)|Finding|false|false|C3686666;C0027530;C3159206;C2987514|NECK
null|Neck problem|Finding|false|false|C3686666;C0027530;C3159206;C2987514|NECKnull|dendritic spine neck|Anatomy|false|false|C1549548;C1705938;C1843354;C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C1549548;C1705938;C1843354;C0812434;C0684335|NECKnull|Visual|Finding|false|false|C0027530;C3159206;C2987514|Visualizednull|nitrogenous base|Drug|false|false|C2987514;C0027530;C3159206|base
null|Base|Drug|false|false|C2987514;C0027530;C3159206|base
null|Dental Base|Drug|false|false|C2987514;C0027530;C3159206|base
null|base - RoleClass|Drug|false|false|C2987514;C0027530;C3159206|basenull|Base - General Qualifier|Finding|false|false|C0027530;C3159206;C2987514|base
null|BPIFA4P gene|Finding|false|false|C0027530;C3159206;C2987514|base
null|Base - RX Component Type|Finding|false|false|C0027530;C3159206;C2987514|basenull|Anatomical base|Anatomy|false|false|C0234621;C0812434;C0684335;C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C2987514|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C2987514|necknull|dendritic spine neck|Anatomy|false|false|C0234621;C1549548;C1705938;C1843354;C0812434;C0684335;C1704464;C0178499;C1550601;C1880279|neck
null|Neck|Anatomy|false|false|C0234621;C1549548;C1705938;C1843354;C0812434;C0684335;C1704464;C0178499;C1550601;C1880279|necknull|Show|Entity|false|false||shownull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Skeletal bone|Anatomy|false|false||BONES
null|XXX bone|Anatomy|false|false||BONESnull|Suspicious|Modifier|false|false||suspiciousnull|Bone Tissue, Human|Anatomy|false|false|C0000768|osseous
null|Skeletal bone|Anatomy|false|false|C0000768|osseousnull|Congenital Abnormality|Disorder|true|false|C4520924;C0262950|abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Fracture|Disorder|false|false||fracturenull|Left breast|Anatomy|false|false|C0496956;C0191838;C0018944;C0567499;C0342095;C1552822|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0006141;C0222601|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Breast hematoma|Finding|false|false|C0006141;C0222601|breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0222601;C0006141|breastnull|Breast problem|Finding|false|false|C0006141;C0222601|breastnull|Procedures on breast|Procedure|false|false|C0222601;C0006141|breastnull|Breast|Anatomy|false|false|C0342095;C1552822;C0567499;C0496956;C0018944;C0191838|breastnull|Hematoma|Finding|false|false|C0222601;C0006141|hematomanull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|false|false||bleednull|Timing, LOINC Axis 3|Finding|false|false||timingnull|Timing|Time|false|false||timingnull|Suboptimal|Modifier|false|false||suboptimalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Due to|Finding|false|false||due
null|Due|Finding|false|false||duenull|Document Completion - incomplete|Finding|false|false||incompletenull|Incomplete|Modifier|false|false||incompletenull|Partial|LabModifier|false|false||incompletenull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|View|Modifier|false|false||viewnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|density|LabModifier|false|false||densitynull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Series|LabModifier|false|false||seriesnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0851238;C0191838;C1552822;C0496956;C0557854;C0191838;C0496956;C3245478;C0567499;C2140215;C0567499|breastnull|ActInformationPrivacyReason - service|Finding|false|false|C0222601;C0006141;C0006141|servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false|C0006141;C0222601|servicenull|Lumpectomy of left breast|Procedure|false|false|C0222601;C0006141;C0006141|left breast lumpectomynull|Left breast|Anatomy|false|false|C2140215;C1552822;C3245478;C0191838;C0496956;C0851238;C1262070;C0851238;C0567499;C0557854|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0006141;C0222601;C0006141|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lumpectomy of breast|Procedure|false|false|C0006141;C0006141;C0222601|breast lumpectomynull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141;C0222601;C0006141|breastnull|Breast problem|Finding|false|false|C0006141;C0222601;C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141;C0222601;C0006141|breastnull|Breast|Anatomy|false|false|C0851238;C2140215;C1552822;C0567499;C0496956;C0851238;C1262070;C3245478;C0191838|breastnull|Lumpectomy of breast|Procedure|false|false|C0222601;C0006141|lumpectomy
null|Excision of mass (procedure)|Procedure|false|false|C0222601;C0006141|lumpectomynull|Invasive|Modifier|false|false||invasivenull|Carcinoma|Disorder|false|false||carcinomanull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Left breast|Anatomy|false|false|C0018944;C1720922;C1546717;C2243017;C1552822;C0567499;C0496956;C0191838;C0342095|left breastnull|Table Cell Horizontal Align - left|Finding|false|false|C0006141;C0222601|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Breast hematoma|Finding|false|false|C0006141;C0222601|breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141;C0222601|breastnull|Breast problem|Finding|false|false|C0006141;C0222601|breastnull|Procedures on breast|Procedure|false|false|C0006141;C0222601|breastnull|Breast|Anatomy|false|false|C1552822;C0567499;C0191838;C0342095;C0496956;C0018944|breastnull|Hematoma|Finding|false|false|C0222601;C0006141|hematomanull|null|Procedure|false|false|C0222601|needle aspirationnull|Aspiration needles|Device|false|false||needle aspirationnull|null|Finding|false|false|C0222601|needlenull|Needle device|Device|false|false||needlenull|Needle Shape|Modifier|false|false||needlenull|Respiratory Aspiration|Disorder|false|false|C0222601|aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Examination and observation for unspecified reason|Finding|false|false||observation
null|null|Finding|false|false||observation
null|null|Finding|false|false||observation
null|Observation (finding)|Finding|false|false||observationnull|Observation - diagnostic procedure|Procedure|false|false||observation
null|Observation in research|Procedure|false|false||observation
null|Patient observation|Procedure|false|false||observationnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Evacuation procedure|Procedure|false|false||evacuationnull|Hematoma|Finding|false|false||hematomanull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Evacuation procedure|Procedure|false|false||evacuationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hematoma|Finding|false|false||hematomanull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Surgical drains|Device|false|false||surgical drainnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Hospital course|Finding|false|false||Hospital coursenull|null|Attribute|false|false||Hospital coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||coursenull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986;C0221776|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|per protocol|Finding|false|false||per protocol
null|On Protocol Therapy|Finding|false|false||per protocolnull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Perioperative Period|Time|false|false||perioperative periodnull|perioperative|Time|false|false||perioperativenull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Issue (document)|Finding|true|false||issue
null|Problem|Finding|true|false||issuenull|Issue (action)|Event|true|false||issuenull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Heme|Drug|false|false||Heme
null|Heme|Drug|false|false||Hemenull|Daily|Time|false|false||dailynull|Laboratory test finding|Lab|false|false||labsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Boots|Device|false|false||bootsnull|Boots pharmaceutical company|Entity|false|false||bootsnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Ancef|Drug|false|false||ancef
null|Ancef|Drug|false|false||ancefnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Apyrexial|Finding|false|false||afebrilenull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Endocrine System Diseases|Disorder|false|false||Endo
null|Endometriosis|Disorder|false|false||Endonull|MANEA gene|Finding|false|false||Endonull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Metabolic Syndrome X|Disorder|false|false||metabolic syndromenull|Metabolic Process, Cellular|Finding|false|false||metabolic
null|Metabolic|Finding|false|false||metabolicnull|Multisection metabolic|Procedure|false|false||metabolicnull|Syndrome|Disorder|false|false||syndromenull|Prediabetes syndrome|Disorder|false|false||pre-diabetesnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Carbohydrate diet|Procedure|false|false||carbohydrate dietnull|Carbohydrates|Drug|false|false||carbohydratenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919;C4284232;C1549543;C0030193;C0221776|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false|C0226896|pain
null|Pain|Finding|false|false|C0226896|painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false|C0226896|medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Apyrexial|Finding|false|false||afebrilenull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Early|Time|false|false||earlynull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Active medication list|Finding|false|false||Active Medication listnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|prescription document|Finding|false|false||Prescriptionnull|Prescription (procedure)|Procedure|false|false||Prescriptionnull|Prescription (attribute)|Attribute|false|false||Prescriptionnull|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATE
null|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATEnull|albuterol|Drug|false|false||ALBUTEROL
null|albuterol|Drug|false|false||ALBUTEROLnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATE
null|Sulfates, Inorganic|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATEnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|Solution Dosage Form|Drug|false|false||solution
null|Solutions|Drug|false|false||solution
null|Pharmaceutical Solutions|Drug|false|false||solutionnull|Resolution|Finding|false|false||solutionnull|nebulization-mediated drug administration|Procedure|false|false||nebulizationnull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATE
null|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATEnull|albuterol|Drug|false|false||ALBUTEROL
null|albuterol|Drug|false|false||ALBUTEROLnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATE
null|Sulfates, Inorganic|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATEnull|ProAir|Drug|false|false||PROAIR HFA
null|ProAir|Drug|false|false||PROAIR HFAnull|ProAir|Drug|false|false||PROAIR
null|ProAir|Drug|false|false||PROAIR
null|Pro-Air Procaterol|Drug|false|false||PROAIR
null|Pro-Air Procaterol|Drug|false|false||PROAIRnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Aerosol Dose Form|Drug|false|false||aerosolnull|Aerosols|Device|false|false||aerosolnull|Puff Dosing Unit|LabModifier|false|false||puffsnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||ATORVASTATIN
null|atorvastatin|Drug|false|false||ATORVASTATINnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false|C1138603;C1555587|mouth
null|Oral region|Anatomy|false|false|C1138603;C1555587|mouthnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Transaction counts and value totals - provider|Finding|false|false|C0230028;C0226896|Provider
null|Provider|Finding|false|false|C0230028;C0226896|Providernull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Adjustment - classification term|Finding|false|false||adjustment
null|Personal Adjustment|Finding|false|false||adjustment
null|null|Finding|false|false||adjustment
null|Psychological adjustment|Finding|false|false||adjustment
null|Transaction Type - Adjustment|Finding|false|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|enoxaparin|Drug|false|false||ENOXAPARIN
null|enoxaparin|Drug|false|false||ENOXAPARINnull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Kilogram per Cubic Meter|LabModifier|false|false||mg/mLnull|per milliliter|LabModifier|false|false||/mLnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Syringes|Device|false|false||syringenull|Syringe (unit of presentation)|LabModifier|false|false||syringe
null|Syringe Dosing Unit|LabModifier|false|false||syringenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Approximate|Modifier|false|false||approximatelynull|12 hours (qualifier value)|Time|false|false||12 hoursnull|Hour|Time|false|false||hoursnull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Adjustment - classification term|Finding|false|false||adjustment
null|Personal Adjustment|Finding|false|false||adjustment
null|null|Finding|false|false||adjustment
null|Psychological adjustment|Finding|false|false||adjustment
null|Transaction Type - Adjustment|Finding|false|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|erythromycin|Drug|false|false||ERYTHROMYCIN
null|erythromycin|Drug|false|false||ERYTHROMYCINnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|gram|LabModifier|false|false||gramnull|Ophthalmic Ointment|Drug|false|false|C4266572;C0015392;C0700042|eye ointmentnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C0304651|eye
null|Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C0304651|eye
null|Orbital region|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477;C0304651|eyenull|Ointments|Drug|false|false||ointmentnull|Apply (administration method)|Finding|false|false||Apply
null|Apply (instruction)|Finding|false|false||Apply
null|null|Finding|false|false||Apply
null|Apply|Finding|false|false||Applynull|Inch Unit of Length|LabModifier|false|false||inchnull|Carcinoma in situ of eye|Disorder|false|false|C4266572;C0015392;C0700042|eye
null|Disorder of eye|Disorder|false|false|C4266572;C0015392;C0700042|eyenull|Eye - Specimen Source Code|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye problem|Finding|false|false|C4266572;C0015392;C0700042|eye
null|Eye Specimen|Finding|false|false|C4266572;C0015392;C0700042|eyenull|Head>Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477|eye
null|Eye|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477|eye
null|Orbital region|Anatomy|false|false|C0154094;C0015397;C1550636;C1546630;C0262477|eyenull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|furosemide|Drug|false|false||FUROSEMIDE
null|furosemide|Drug|false|false||FUROSEMIDEnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|leg swellingnull|Leg|Anatomy|false|false|C0581394|leg
null|Lower Extremity|Anatomy|false|false|C0581394|legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|hydromorphone|Drug|false|false||HYDROMORPHONE
null|hydromorphone|Drug|false|false||HYDROMORPHONEnull|hydromorphone|Drug|false|false||hydromorphone
null|hydromorphone|Drug|false|false||hydromorphonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Drink (dietary substance)|Drug|false|false||drinknull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Nebulizers|Device|false|false||NEBULIZERnull|Compressor Air Pump Device|Device|false|false||COMPRESSORnull|Portable nebuliser system|Device|false|false||PORTABLE NEBULIZER SYSTEMnull|Portable|Modifier|false|false||PORTABLEnull|Nebulizers|Device|false|false||NEBULIZERnull|System (basic dose form)|Drug|false|false||SYSTEMnull|System, LOINC Axis 4|Finding|false|false||SYSTEM
null|System|Finding|false|false||SYSTEMnull|Device system|Device|false|false||SYSTEM
null|System - kit|Device|false|false||SYSTEMnull|System (unit of presentation)|LabModifier|false|false||SYSTEMnull|Portable|Modifier|false|false||Portablenull|Nebulizers|Device|false|false||Nebulizernull|System (basic dose form)|Drug|false|false||Systemnull|System, LOINC Axis 4|Finding|false|false||System
null|System|Finding|false|false||Systemnull|Device system|Device|false|false||System
null|System - kit|Device|false|false||Systemnull|System (unit of presentation)|LabModifier|false|false||Systemnull|Use - dosing instruction imperative|Finding|false|false||Use
null|utilization qualifier|Finding|false|false||Use
null|Usage|Finding|false|false||Usenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Nebulizers|Device|false|false||nebulizernull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|omeprazole|Drug|false|false||OMEPRAZOLE
null|omeprazole|Drug|false|false||OMEPRAZOLEnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|release
null|Released (action)|Finding|false|false|C0524463;C1325531|releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|CAPSULEnull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|CAPSULE
null|Structure of organ capsule|Anatomy|false|false|C0006935|CAPSULEnull|Capsule Shape|Modifier|false|false||CAPSULEnull|Capsule (unit of presentation)|LabModifier|false|false||CAPSULE
null|Capsule Dosing Unit|LabModifier|false|false||CAPSULEnull|Twice a day|Time|false|false||TWICE DAILYnull|Daily|Time|false|false||DAILYnull|gastroesophageal|Anatomy|false|false||GASTROESOPHAGEALnull|sertraline|Drug|false|false||SERTRALINE
null|sertraline|Drug|false|false||SERTRALINEnull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|tramadol|Drug|false|false||TRAMADOL
null|tramadol|Drug|false|false||TRAMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TRAMADOLnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|trazodone|Drug|false|false||TRAZODONE
null|trazodone|Drug|false|false||TRAZODONEnull|trazodone|Drug|false|false||trazodone
null|trazodone|Drug|false|false||trazodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|warfarin|Drug|false|false||WARFARIN
null|warfarin|Drug|false|false||WARFARIN
null|warfarin|Drug|false|false||WARFARINnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Five times weekly|Time|false|false||5 times a weeknull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false|C0449201|pernull|Per - dosing instruction fragment|Finding|false|false|C0449201|per
null|PER1 gene|Finding|false|false|C0449201|per
null|Follow|Finding|false|false|C0449201|per
null|PER1 wt Allele|Finding|false|false|C0449201|pernull|PER (body structure)|Anatomy|false|false|C3273590;C4281991;C1418464;C1704764;C1861457|pernull|Per (qualifier)|Modifier|false|false||pernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Adjustment - classification term|Finding|false|false||adjustment
null|Personal Adjustment|Finding|false|false||adjustment
null|null|Finding|false|false||adjustment
null|Psychological adjustment|Finding|false|false||adjustment
null|Transaction Type - Adjustment|Finding|false|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|Acetaminophen [EPC]|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHENnull|Acetaminophen measurement|Procedure|false|false||ACETAMINOPHENnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Multiple Epiphyseal Dysplasia|Disorder|false|false||mednull|Master of Education|Finding|false|false||med
null|COMP wt Allele|Finding|false|false||med
null|COL9A3 gene|Finding|false|false||med
null|SCN8A wt Allele|Finding|false|false||med
null|COL9A2 gene|Finding|false|false||med
null|COMP gene|Finding|false|false||med
null|SCN8A gene|Finding|false|false||mednull|ZDHHC2 protein, human|Drug|false|false||rec
null|ZDHHC2 protein, human|Drug|false|false||recnull|RBPJP4 gene|Finding|false|false||rec
null|MCM8 gene|Finding|false|false||recnull|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROLnull|vitamin D3|Drug|false|false||VITAMIN D3
null|vitamin D3|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMINnull|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferolnull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1720092;C1561538;C1561539|mouth
null|Oral region|Anatomy|false|false|C1527415;C1720092;C1561538;C1561539|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false|C0230028;C0226896|oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|polyethylene glycol 3350|Drug|false|false||POLYETHYLENE GLYCOL 3350
null|polyethylene glycol 3350|Drug|false|false||POLYETHYLENE GLYCOL 3350null|polyethylene glycols|Drug|false|false||POLYETHYLENE GLYCOL
null|polyethylene glycols|Drug|false|false||POLYETHYLENE GLYCOLnull|high-density polyethylene|Drug|false|false||POLYETHYLENE
null|high-density polyethylene|Drug|false|false||POLYETHYLENE
null|polyethylenes|Drug|false|false||POLYETHYLENE
null|polyethylenes|Drug|false|false||POLYETHYLENE
null|Polyethylene|Drug|false|false||POLYETHYLENE
null|Polyethylene|Drug|false|false||POLYETHYLENEnull|ethylene glycol|Drug|false|false||GLYCOL
null|Glycol|Drug|false|false||GLYCOL
null|ethylene glycol|Drug|false|false||GLYCOL
null|Glycols|Drug|false|false||GLYCOLnull|Miralax|Drug|false|false||MIRALAX
null|Miralax|Drug|false|false||MIRALAXnull|Miralax|Drug|false|false||Miralax
null|Miralax|Drug|false|false||Miralaxnull|gram|LabModifier|false|false||gramnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|powder physical state|Drug|false|false||powder
null|Powder dose form|Drug|false|false||powdernull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Dose Adjustment|Procedure|false|false||Dose adjustmentnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Adjustment - classification term|Finding|false|false||adjustment
null|Personal Adjustment|Finding|false|false||adjustment
null|null|Finding|false|false||adjustment
null|Psychological adjustment|Finding|false|false||adjustment
null|Transaction Type - Adjustment|Finding|false|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|sennosides, USP|Drug|false|false||SENNOSIDES
null|sennosides, USP|Drug|false|false||SENNOSIDESnull|sennosides, USP|Drug|false|false||SENNA
null|sennosides, USP|Drug|false|false||SENNAnull|Senna alexandrina|Entity|false|false||SENNA
null|Senna Plant|Entity|false|false||SENNAnull|sennosides, USP|Drug|false|false||senna
null|sennosides, USP|Drug|false|false||sennanull|Senna alexandrina|Entity|false|false||senna
null|Senna Plant|Entity|false|false||sennanull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Indication of (contextual qualifier)|Finding|false|false||Reason fornull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Duplicate component (foundation metadata concept)|Finding|false|false||duplicate
null|Double (qualifier value)|Finding|false|false||duplicatenull|Replicate|Event|false|false||duplicatenull|Duplicate|Modifier|false|false||duplicatenull|Override|Finding|false|false||overridenull|Similarity|Modifier|false|false||similarnull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1422467|mouth
null|Oral region|Anatomy|false|false|C1527415;C1422467|mouthnull|CIAO3 gene|Finding|false|false|C0230028;C0226896|prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Breast hematoma|Finding|false|false|C0006141|breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0496956;C0567499;C0018944;C0342095;C0191838|breastnull|Hematoma|Finding|false|false|C0006141|hematomanull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Self-care interventions|Finding|false|false||Personal Carenull|Personal Attribute|Subject|false|false||Personalnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Surgical incisions|Procedure|false|false||incisionsnull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Cleaning (activity)|Event|false|false||cleannull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Gauzes|Device|false|false||gauzenull|Daily|Time|false|false||dailynull|Cleaning (activity)|Event|false|false||Cleannull|Drain - SpecimenType|Drug|false|false|C1515974|drainnull|Drain Specimen Code|Finding|false|false|C1515974|drainnull|Drain device|Device|false|false||drainnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C1546604;C1550628|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Tubing|Device|false|false||tubingnull|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1547961;C0178298;C0496955;C0020311;C1546781;C0444099;C1705308|skin
null|Skin|Anatomy|false|false|C1547961;C0178298;C0496955;C0020311;C1546781;C0444099;C1705308|skinnull|Soap Dosage Form|Drug|false|false|C1123023;C4520765|soapnull|Soap|Device|false|false||soapnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false|C1123023;C4520765|waternull|Hydrotherapy|Procedure|false|false|C1123023;C4520765|waternull|Compliance Package - Strip|Drug|false|false||Strip
null|Strip Dosage Form|Drug|false|false||Stripnull|strip medical device|Device|false|false||Stripnull|Strip - unit of product usage|LabModifier|false|false||Strip
null|Strip (unit of presentation)|LabModifier|false|false||Strip
null|Strip Dosing Unit|LabModifier|false|false||Stripnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Tubing|Device|false|false||tubingnull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|anatomical bulb|Anatomy|false|false||bulb
null|Medulla Oblongata|Anatomy|false|false||bulbnull|plant bulb|Entity|false|false||bulbnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|written - ParticipationMode|Finding|false|false||written
null|Written - Consent Mode|Finding|false|false||writtennull|Record of (contextual qualifier)|Modifier|false|false||record ofnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|Daily|Time|false|false||dailynull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Drain device|Device|false|false||drainsnull|As soon as possible|Time|false|false||as soon as possiblenull|Possible|Finding|false|false||possiblenull|Possibly Related to Intervention|Modifier|false|false||possible
null|Possible diagnosis|Modifier|false|false||possiblenull|Daily|Time|false|false||dailynull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Acceptable (foundation metadata concept)|Modifier|false|false||acceptable
null|Acceptable|Modifier|false|false||acceptablenull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Operative Surgical Procedures|Procedure|false|false|C0006104|surgical
null|Surgical service|Procedure|false|false|C0006104|surgicalnull|Brain|Anatomy|false|false|C0543467;C0587668|branull|Brassiere|Device|false|false||branull|Braj Language|Entity|false|false||branull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Loose|Modifier|false|false||loosenull|Camisole|Device|false|false||camisolenull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|DERMABOND|Drug|false|false|C1123023;C4520765|Dermabond
null|DERMABOND|Drug|false|false|C1123023;C4520765|Dermabondnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1530215;C0178298;C0496955;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C1530215;C0178298;C0496955;C1546781;C0444099|skinnull|Glues|Drug|false|false||gluenull|day|Time|false|false||daysnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Walking (function)|Finding|false|false||Walknull|More than once a day|Time|false|false||several times a daynull|Several|LabModifier|false|false||severalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Pounds|LabModifier|false|false||poundsnull|Strenuous Exercise|Finding|false|false||strenuous activitynull|Strenuous|Modifier|false|false||strenuousnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Regular|Modifier|false|false||regularnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenol
null|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenolnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Mild pain|Finding|false|false||mild pain
null|Neck Pain Score 2|Finding|false|false||mild painnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Packaging Materials|Device|false|false||packaging
null|Drug Packaging|Device|false|false||packagingnull|Packaging|Phenomenon|false|false||packagingnull|Packing (action)|Event|false|false||packagingnull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|Vicodin|Drug|false|false||Vicodin
null|Vicodin|Drug|false|false||Vicodinnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Active ingredient|Drug|false|false||active ingredientnull|Has active ingredient|Modifier|false|false||active ingredientnull|Ingredient|Drug|false|false||ingredientnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Additional|Finding|false|false||additionalnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C5975557;C3844164;C1527415;C4035627|mouth
null|Oral region|Anatomy|false|false|C5975557;C3844164;C1527415;C4035627|mouthnull|2 times per day|Finding|false|false|C0230028;C0226896|2 times per daynull|2 times|Finding|false|false|C0230028;C0226896|2 timesnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false|C0230028;C0226896|timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Different|Modifier|false|false||differentnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Have Constipation|Finding|false|false||have constipationnull|Constipation|Finding|false|false||constipationnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Etc.|Finding|false|false||etcnull|Drinking (function)|Finding|false|false||drinking
null|Alcohol consumption|Finding|false|false||drinkingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Stool Softener|Drug|false|false||stool softenersnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Food|Drug|false|false||foodsnull|Message Waiting Priority - High|Finding|false|false|C1304649|high
null|high - ActExposureLevelCode|Finding|false|false|C1304649|high
null|IPSS Risk Category High|Finding|false|false|C1304649|high
null|IPSS-R Risk Category High|Finding|false|false|C1304649|high
null|High (finding)|Finding|false|false|C1304649|highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fibernull|Tissue fiber|Anatomy|false|false|C3887512;C5200928;C1561958;C4522209;C5202936;C0225326;C1321801|fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Fever with chills|Finding|false|false||fever with chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Physiologic warmth|Finding|false|false|C1515974|warmth
null|Social warmth|Finding|false|false|C1515974|warmthnull|Emotional tenderness|Finding|false|false|C1515974|tenderness
null|Sore to touch|Finding|false|false|C1515974|tendernessnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0543467;C0587668;C0684239;C0234233;C0518610;C0392197;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Unusual|Modifier|false|false||unusualnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false|C2338258|drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0013103;C0332803|incisionnull|Large amount|LabModifier|false|false||large amountnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Amount class - Amount|Finding|false|false|C2338258|amountnull|Quantity|LabModifier|false|false||amountnull|Hemorrhage|Finding|false|false|C2338258|bleedingnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0019080;C0332803;C1561574|incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Severe Extremity Pain|Finding|false|false||Severe pain
null|Severe pain|Finding|false|false||Severe pain
null|Neck Pain Score 6|Finding|false|false||Severe painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false|C2338258|dischargenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0030685;C0332803|incisionnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Else|Finding|false|false||elsenull|Equipment Alert Level - Serious|Finding|false|false||serious
null|Device Alert Level - Serious|Finding|false|false||serious
null|Alert level - Serious|Finding|false|false||seriousnull|Serious|Modifier|false|false||seriousnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Concern|Finding|false|false||concernnull|ANTICOAGULATION (finding)|Finding|false|false||ANTICOAGULATION
null|Anticoagulation function|Finding|false|false||ANTICOAGULATION
null|Decreased Coagulation Activity [PE]|Finding|false|false||ANTICOAGULATIONnull|Anticoagulation Therapy|Procedure|false|false||ANTICOAGULATIONnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|warfarin dose|Procedure|false|false||warfarin dosenull|null|Attribute|false|false||warfarin dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Evening|Time|false|false||eveningnull|Resume - Remote control command|Finding|false|false||resume
null|Curriculum Vitae|Finding|false|false||resume
null|resume - DataOperation|Finding|false|false||resumenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Regular|Modifier|false|false||regularnull|Dosage|LabModifier|false|false||dosesnull|Bridge Therapy|Procedure|false|false||bridge therapynull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Drain - SpecimenType|Drug|false|false||DRAINnull|Drain Specimen Code|Finding|false|false||DRAINnull|Drain device|Device|false|false||DRAINnull|Discharge instructions|Finding|false|false||DISCHARGE INSTRUCTIONSnull|hospital discharge instructions (treatment)|Procedure|false|false||DISCHARGE INSTRUCTIONSnull|null|Attribute|false|false||DISCHARGE INSTRUCTIONSnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Instructions|Finding|false|false||INSTRUCTIONS
null|Instruction [Publication Type]|Finding|false|false||INSTRUCTIONSnull|null|Attribute|false|false||INSTRUCTIONSnull|Drain device|Device|false|false||drainsnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Drain - SpecimenType|Drug|false|false||Drainnull|Drain Specimen Code|Finding|false|false||Drainnull|Drain device|Device|false|false||Drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Cleaning (activity)|Event|false|false||cleannull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Hand|Anatomy|false|false||handsnull|Thoroughly|Finding|false|false||thoroughlynull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Daily|Time|false|false||each daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Does pull|Finding|false|false||Pullnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|null|Device|false|false||bottlenull|Bottle (unit of presentation)|LabModifier|false|false||bottle
null|Bottle Dosing Unit|LabModifier|false|false||bottlenull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Carcinoma of unknown primary|Disorder|false|false||cupnull|Cup (physical object)|Device|false|false||cup
null|Cup Device|Device|false|false||cupnull|Cup (unit of presentation)|LabModifier|false|false||cup
null|Cup Dosing Unit|LabModifier|false|false||cupnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|Suction drain|Device|false|false||drain suctionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Suction drainage|Procedure|false|false||suctionnull|Location Equipment - Suction|Modifier|false|false||suctionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Daily|Time|false|false||dailynull|Event Log|Finding|false|false|C0228228|lognull|lateral occipital gyrus (human only)|Anatomy|false|false|C1708728;C3245468|lognull|Logarithm|LabModifier|false|false||lognull|Individual - insurance coverage level|Finding|false|false|C0228228|individualnull|Individual|Subject|false|false||individual
null|Persons|Subject|false|false||individualnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Appointments|Event|false|false||appointmentnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions