 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|163,172|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|163,172|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|178,181|false|false|false|C0013343|Dyes|Dye
Drug|Biologically Active Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|SIMPLE_SEGMENT|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|SIMPLE_SEGMENT|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|SIMPLE_SEGMENT|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|SIMPLE_SEGMENT|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Organic Chemical|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|244,255|false|false|false|C1569608|varenicline|Varenicline
Finding|Functional Concept|SIMPLE_SEGMENT|258,267|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|276,291|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|282,291|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|282,291|false|false|false|C5441521|Complaint (finding)|Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|293,312|false|false|false|C2707305||Shortness of Breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|293,312|false|false|false|C0013404|Dyspnea|Shortness of Breath
Finding|Body Substance|SIMPLE_SEGMENT|306,312|false|false|false|C0225386|Breath|Breath
Finding|Classification|SIMPLE_SEGMENT|316,321|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|334,352|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|343,352|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|343,352|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|343,352|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|343,352|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,371|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|361,387|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|361,387|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|372,379|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|372,379|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|372,387|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|380,387|false|false|false|C0221423|Illness (finding)|Illness
Finding|Conceptual Entity|SIMPLE_SEGMENT|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|418,428|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|430,434|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|430,434|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|430,434|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|SIMPLE_SEGMENT|438,442|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|438,442|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|438,442|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|447,453|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|447,466|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|447,466|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|447,466|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|454,466|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|470,478|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|470,478|false|false|false|C1831808|apixaban|apixaban
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|480,492|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|495,498|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|495,498|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|495,498|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|495,498|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|504,518|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|504,518|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Attribute|Clinical Attribute|SIMPLE_SEGMENT|537,556|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|537,556|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|550,556|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|559,564|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|559,564|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|559,564|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|570,578|false|false|false|C0043144|Wheezing|wheezing
Finding|Idea or Concept|SIMPLE_SEGMENT|587,590|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|587,590|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|SIMPLE_SEGMENT|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|605,632|false|false|false|C4718286|Reports shortness of breath|reports shortness of breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|613,632|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|613,632|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|626,632|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|644,649|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|644,649|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|644,649|false|false|false|C0010200|Coughing|cough
Finding|Finding|SIMPLE_SEGMENT|669,672|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|669,672|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Body Substance|SIMPLE_SEGMENT|681,687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|681,687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Sign or Symptom|SIMPLE_SEGMENT|693,701|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|748,757|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|748,757|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|789,800|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|789,800|false|false|false|C0027235|ipratropium|ipratropium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|801,805|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|SIMPLE_SEGMENT|834,840|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|834,840|false|false|false|C0723011|Relief brand of phenylephrine|relief
Finding|Finding|SIMPLE_SEGMENT|834,840|false|false|false|C0564405|Feeling relief|relief
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|869,873|false|false|false|C0806140|Flow|flow
Finding|Idea or Concept|SIMPLE_SEGMENT|892,903|false|false|false|C0750502|Significant|significant
Finding|Conceptual Entity|SIMPLE_SEGMENT|904,915|false|false|false|C2986411|Improvement|improvement
Finding|Finding|SIMPLE_SEGMENT|925,941|false|false|false|C3843777|Currently taking|currently taking
Drug|Hormone|SIMPLE_SEGMENT|951,961|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|951,961|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|951,961|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|988,998|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|988,998|false|false|false|C0213771|tiotropium|tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|1004,1016|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1004,1016|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1004,1016|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|1018,1024|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1018,1024|false|false|false|C0965130|Advair|advair
Finding|Finding|SIMPLE_SEGMENT|1028,1035|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1031,1035|false|false|false|C1553498|home health encounter|home
Finding|Sign or Symptom|SIMPLE_SEGMENT|1062,1066|false|false|false|C0221423|Illness (finding)|sick
Procedure|Health Care Activity|SIMPLE_SEGMENT|1068,1076|false|false|false|C4036459|Contacts|contacts
Finding|Idea or Concept|SIMPLE_SEGMENT|1111,1116|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|1111,1116|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|SIMPLE_SEGMENT|1117,1120|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1149,1154|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1149,1154|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1149,1159|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1149,1159|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1155,1159|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1155,1159|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1155,1159|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1251,1256|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1251,1256|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1257,1263|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1265,1274|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1265,1279|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1275,1279|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1275,1279|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1275,1279|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1281,1287|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1281,1287|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1281,1296|true|false|false|C0027498|Nausea and vomiting|nausea/vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|1288,1296|true|false|false|C0042963|Vomiting|vomiting
Finding|Finding|SIMPLE_SEGMENT|1299,1311|false|false|false|C0030252|Palpitations|palpitations
Finding|Finding|SIMPLE_SEGMENT|1317,1328|false|false|false|C0700590|Increased sweating|diaphoresis
Finding|Finding|SIMPLE_SEGMENT|1379,1386|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1379,1386|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1411,1420|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|SIMPLE_SEGMENT|1411,1420|false|false|false|C1522484|metastatic qualifier|secondary
Drug|Organic Chemical|SIMPLE_SEGMENT|1424,1431|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1424,1431|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Health Care Activity|SIMPLE_SEGMENT|1432,1437|false|false|false|C0441640||taper
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1449,1453|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1449,1453|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1449,1453|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|1455,1467|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1475,1484|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1475,1484|false|false|false|C1179435|Protein Component|component
Finding|Conceptual Entity|SIMPLE_SEGMENT|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1488,1495|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|1488,1495|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Intellectual Product|SIMPLE_SEGMENT|1504,1509|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1510,1514|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1510,1514|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|1510,1514|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|1516,1528|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Organic Chemical|SIMPLE_SEGMENT|1551,1559|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1551,1559|false|false|false|C0038317|Steroids|steroids
Drug|Antibiotic|SIMPLE_SEGMENT|1580,1591|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1618,1627|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|1618,1627|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Finding|Idea or Concept|SIMPLE_SEGMENT|1635,1643|true|false|false|C3887511|Evidence|evidence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1648,1657|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|1648,1657|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1671,1680|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1671,1680|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|1671,1680|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Drug|Organic Chemical|SIMPLE_SEGMENT|1727,1733|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1727,1733|false|false|false|C0965130|Advair|Advair
Drug|Organic Chemical|SIMPLE_SEGMENT|1786,1798|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1786,1798|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1786,1798|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|1803,1814|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1803,1814|false|false|false|C0965618|roflumilast|roflumilast
Finding|Functional Concept|SIMPLE_SEGMENT|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Idea or Concept|SIMPLE_SEGMENT|1838,1842|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|1838,1842|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Antibiotic|SIMPLE_SEGMENT|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Finding|Finding|SIMPLE_SEGMENT|1856,1863|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|1856,1863|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1856,1863|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Classification|SIMPLE_SEGMENT|1889,1899|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|1889,1899|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|SIMPLE_SEGMENT|1900,1906|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|1900,1906|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|1900,1909|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|1900,1909|false|false|false|C1522577|follow-up|follow-up
Drug|Organic Chemical|SIMPLE_SEGMENT|1935,1942|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1935,1942|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Hormone|SIMPLE_SEGMENT|1960,1970|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|1960,1970|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1960,1970|false|false|false|C0032952|prednisone|prednisone
Finding|Intellectual Product|SIMPLE_SEGMENT|1989,1993|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|2013,2017|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Classification|SIMPLE_SEGMENT|2030,2040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|2030,2040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|SIMPLE_SEGMENT|2041,2047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|2041,2047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|2041,2050|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|2041,2050|false|false|false|C1522577|follow-up|follow-up
Finding|Idea or Concept|SIMPLE_SEGMENT|2064,2071|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|SIMPLE_SEGMENT|2072,2077|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2072,2083|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2072,2083|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|2078,2083|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2078,2083|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2117,2121|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2117,2121|false|false|false|C0582103|Medical Examination|Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2138,2145|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|SIMPLE_SEGMENT|2138,2145|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2146,2158|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|2150,2158|false|false|false|C0026649|Movement|movement
Finding|Sign or Symptom|SIMPLE_SEGMENT|2164,2172|false|false|false|C0043144|Wheezing|wheezing
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2187,2191|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|SIMPLE_SEGMENT|2209,2212|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2233,2236|false|false|false|C0201617|Primed lymphocyte test|Plt
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2258,2261|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2258,2261|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2258,2261|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|2283,2286|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2283,2286|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Drug|Organic Chemical|SIMPLE_SEGMENT|2292,2299|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2292,2299|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2292,2299|false|false|false|C0202115|Lactic acid measurement|lactate
Finding|Finding|SIMPLE_SEGMENT|2320,2327|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2320,2327|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2333,2336|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|2344,2348|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Pathologic Function|SIMPLE_SEGMENT|2358,2369|false|false|false|C0004144|Atelectasis|atelectasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2393,2406|true|false|false|C0521530|Lung consolidation|consolidation
Finding|Body Substance|SIMPLE_SEGMENT|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|2443,2453|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2443,2453|false|false|false|C0701466|Solu-Medrol|solumedrol
Finding|Functional Concept|SIMPLE_SEGMENT|2481,2489|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|2481,2489|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|2481,2489|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|SIMPLE_SEGMENT|2502,2509|false|false|false|C1706079||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2502,2509|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2517,2522|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2540,2549|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2540,2549|false|false|false|C1160636|respiratory system process|breathing
Finding|Idea or Concept|SIMPLE_SEGMENT|2565,2571|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|2565,2571|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|2565,2574|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2565,2582|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2565,2582|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|2575,2582|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2588,2591|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Finding|Finding|SIMPLE_SEGMENT|2588,2591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|2588,2591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Sign or Symptom|SIMPLE_SEGMENT|2600,2608|true|false|false|C0018681|Headache|headache
Finding|Functional Concept|SIMPLE_SEGMENT|2610,2616|false|false|false|C0234621|Visual|visual
Finding|Finding|SIMPLE_SEGMENT|2610,2624|true|false|false|C0750280|Visual changes|visual changes
Finding|Functional Concept|SIMPLE_SEGMENT|2617,2624|false|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2627,2638|false|false|false|C0031350|Pharyngitis|pharyngitis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2640,2650|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2652,2657|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|2652,2657|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|2652,2657|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|SIMPLE_SEGMENT|2652,2668|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|2658,2668|false|false|false|C0700148|Congestion|congestion
Finding|Sign or Symptom|SIMPLE_SEGMENT|2670,2676|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|2678,2684|false|false|false|C0085593|Chills|chills
Finding|Body Substance|SIMPLE_SEGMENT|2687,2693|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|2687,2693|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2695,2701|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2695,2701|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|2695,2706|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|2695,2706|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|SIMPLE_SEGMENT|2702,2706|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2708,2717|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|2708,2722|false|false|true|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2718,2722|false|false|true|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2718,2722|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2718,2722|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2724,2730|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2724,2730|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2732,2740|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|SIMPLE_SEGMENT|2742,2750|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2742,2750|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2753,2765|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2767,2779|false|false|false|C0018932|Hematochezia|hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2767,2779|false|false|false|C1321898|Blood in stool|hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2781,2788|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2790,2794|false|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|SIMPLE_SEGMENT|2790,2794|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|2790,2794|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2796,2808|false|false|false|C0030554|Paresthesia|paresthesias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2815,2823|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|2827,2847|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|2832,2839|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2832,2839|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2832,2839|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2832,2839|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2832,2847|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2840,2847|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2840,2847|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2840,2847|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2851,2855|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2851,2855|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2851,2855|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2856,2862|false|false|false|C0004096|Asthma|Asthma
Finding|Idea or Concept|SIMPLE_SEGMENT|2866,2870|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2866,2870|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2866,2870|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|2879,2887|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|2879,2898|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2888,2893|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|2888,2893|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2888,2898|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2888,2898|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2894,2898|false|true|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|2894,2898|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2894,2898|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2901,2913|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2916,2930|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|2916,2930|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2951,2957|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2951,2970|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2951,2970|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2951,2970|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2958,2970|false|false|false|C0232197|Fibrillation|Fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|2974,2982|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2974,2982|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2985,2992|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|2985,2992|false|false|false|C0860603|Anxiety symptoms|Anxiety
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2995,3003|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2995,3015|false|false|false|C0263884|Cervical radiculitis|Cervical Radiculitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3004,3015|false|false|false|C0034544|Radiculitis|Radiculitis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3018,3026|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3018,3038|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|Cervical Spondylosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3027,3038|false|false|false|C0038019|Spondylosis|Spondylosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3041,3049|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3041,3056|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3041,3064|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3050,3056|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|SIMPLE_SEGMENT|3050,3056|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3050,3064|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3057,3064|false|false|false|C0012634|Disease|Disease
Finding|Sign or Symptom|SIMPLE_SEGMENT|3067,3075|false|false|false|C0018681|Headache|Headache
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3078,3084|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|Herpes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3078,3091|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Virus|SIMPLE_SEGMENT|3078,3091|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3085,3091|false|false|false|C0019360|Herpes zoster (disorder)|Zoster
Finding|Pathologic Function|SIMPLE_SEGMENT|3094,3105|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|3097,3105|false|false|false|C0019080|Hemorrhage|Bleeding
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3108,3135|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral Vascular Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3119,3127|false|false|false|C0005847|Blood Vessel|Vascular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3119,3135|false|false|false|C0042373|Vascular Diseases|Vascular Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3128,3135|false|false|false|C0012634|Disease|Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3150,3155|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3150,3162|false|false|false|C0850459|iliac stents|iliac stents
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3169,3172|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|3169,3172|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3169,3172|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3169,3184|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Finding|Functional Concept|SIMPLE_SEGMENT|3173,3184|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|3173,3184|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3173,3184|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Functional Concept|SIMPLE_SEGMENT|3187,3193|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3187,3201|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3194,3201|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3194,3201|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3194,3201|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3207,3213|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3207,3213|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3207,3213|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3207,3213|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3207,3221|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3214,3221|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3214,3221|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3214,3221|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|3223,3229|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3235,3241|false|false|false|C0004096|Asthma|asthma
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3246,3258|false|false|false|C0020538|Hypertensive disease|hypertension
Finding|Conceptual Entity|SIMPLE_SEGMENT|3260,3266|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3260,3266|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3272,3277|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3272,3277|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3272,3277|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|3272,3277|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3272,3284|false|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3278,3284|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|3287,3294|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|SIMPLE_SEGMENT|3287,3294|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3300,3308|false|false|false|C0023418|leukemia|leukemia
Finding|Finding|SIMPLE_SEGMENT|3313,3321|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3313,3321|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3313,3321|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3313,3326|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3313,3326|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3322,3326|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3322,3326|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3328,3337|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|SIMPLE_SEGMENT|3338,3346|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3338,3346|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3338,3346|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3338,3351|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3338,3351|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3347,3351|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3347,3351|false|false|false|C0582103|Medical Examination|EXAM
Finding|Gene or Genome|SIMPLE_SEGMENT|3388,3392|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3388,3392|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Classification|SIMPLE_SEGMENT|3442,3449|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3442,3449|false|false|false|C3812897|General medical service|GENERAL
Finding|Intellectual Product|SIMPLE_SEGMENT|3474,3483|false|false|true|C0876929|Sentence|sentences
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3485,3488|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3485,3488|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|3485,3488|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3501,3504|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3501,3504|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3519,3524|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3532,3537|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3545,3551|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3545,3551|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3545,3551|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|SIMPLE_SEGMENT|3552,3561|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3581,3584|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3581,3584|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3586,3596|false|false|false|C0521367|Oropharyngeal|Oropharynx
Finding|Idea or Concept|SIMPLE_SEGMENT|3600,3605|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3607,3611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3607,3611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3607,3611|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|SIMPLE_SEGMENT|3613,3619|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3624,3627|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3624,3627|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3624,3627|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|3629,3632|true|false|false|C0428897|Jugular venous pressure|JVP
Finding|Intellectual Product|SIMPLE_SEGMENT|3655,3662|false|false|false|C0542560|Academic degree|degrees
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3664,3671|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3664,3671|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|SIMPLE_SEGMENT|3703,3707|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3703,3707|false|false|false|C1549480|Amount type - Rate|rate
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3713,3721|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|3713,3728|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|SIMPLE_SEGMENT|3722,3728|false|false|false|C0018808|Heart murmur|murmur
Finding|Finding|SIMPLE_SEGMENT|3747,3751|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3764,3769|false|false|false|C0024109|Lung|LUNGS
Finding|Organism Function|SIMPLE_SEGMENT|3771,3781|false|false|false|C0231800|Expiration, Respiratory|Expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|3771,3789|false|false|false|C0231875|Expiratory wheezing|Expiratory wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3782,3789|false|false|false|C0043144|Wheezing|wheezes
Finding|Intellectual Product|SIMPLE_SEGMENT|3806,3810|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3811,3823|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|3815,3823|false|false|false|C0026649|Movement|movement
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3825,3832|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3825,3832|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3825,3832|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3839,3843|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3874,3885|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Finding|SIMPLE_SEGMENT|3887,3891|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3887,3891|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3896,3900|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3914,3919|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3914,3919|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|3927,3933|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3927,3933|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3927,3933|false|false|false|C0034107|Pulse taking|pulses
Finding|Finding|SIMPLE_SEGMENT|3977,3983|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Idea or Concept|SIMPLE_SEGMENT|3985,3993|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|SIMPLE_SEGMENT|3998,4007|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3998,4007|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3998,4007|false|false|false|C2229507|sensory exam|sensation
Finding|Finding|SIMPLE_SEGMENT|4017,4023|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Body Substance|SIMPLE_SEGMENT|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4038,4047|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|SIMPLE_SEGMENT|4048,4056|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|4048,4056|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4048,4056|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|4048,4061|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4048,4061|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4057,4061|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4057,4061|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|SIMPLE_SEGMENT|4151,4158|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4151,4158|false|false|false|C3812897|General medical service|GENERAL
Finding|Intellectual Product|SIMPLE_SEGMENT|4177,4186|false|false|false|C0876929|Sentence|sentences
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4188,4191|false|false|true|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4188,4191|false|false|true|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|4188,4191|false|false|true|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4204,4207|false|false|true|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|4204,4207|false|false|true|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4222,4229|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|4222,4229|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|SIMPLE_SEGMENT|4243,4247|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4243,4247|false|false|false|C1549480|Amount type - Rate|rate
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4253,4261|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|4253,4268|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|SIMPLE_SEGMENT|4262,4268|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4281,4286|false|false|false|C0024109|Lung|LUNGS
Finding|Intellectual Product|SIMPLE_SEGMENT|4289,4293|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Sign or Symptom|SIMPLE_SEGMENT|4294,4301|false|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4313,4320|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4313,4320|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4313,4320|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4327,4331|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4362,4373|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Finding|SIMPLE_SEGMENT|4375,4379|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4375,4379|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|4384,4388|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4410,4415|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4410,4415|false|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|SIMPLE_SEGMENT|4475,4484|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4485,4489|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4530,4535|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4530,4535|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4536,4539|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4544,4547|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4544,4547|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4544,4547|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4553,4556|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4553,4556|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4553,4556|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4553,4556|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4562,4565|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4562,4565|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4571,4574|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4571,4574|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4579,4582|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4579,4582|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4579,4582|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4579,4582|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4579,4582|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4588,4592|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4621,4624|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4641,4646|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4641,4646|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4659,4665|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4682,4685|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4682,4685|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4786,4791|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4786,4791|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4786,4799|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4792,4799|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4792,4799|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4832,4837|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4832,4837|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Classification|SIMPLE_SEGMENT|4842,4845|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|4842,4845|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4842,4845|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4850,4854|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4850,4854|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4880,4884|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|4880,4884|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|4880,4884|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4902,4907|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4902,4907|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4902,4915|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|4908,4915|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4908,4915|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4908,4915|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4932,4937|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4932,4937|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4938,4944|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|4938,4944|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4961,4966|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4961,4966|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Research Activity|SIMPLE_SEGMENT|4982,4989|false|false|false|C0947630|Scientific Study|STUDIES
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5020,5023|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|5031,5035|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Pathologic Function|SIMPLE_SEGMENT|5036,5055|false|false|false|C4049574|Basilar atelectasis|basilar atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|5044,5055|false|false|false|C0004144|Atelectasis|atelectasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5080,5093|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Intellectual Product|SIMPLE_SEGMENT|5097,5100|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5097,5100|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5102,5107|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5102,5107|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|5102,5107|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5102,5107|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|SIMPLE_SEGMENT|5102,5114|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Finding|Finding|SIMPLE_SEGMENT|5108,5114|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|5108,5114|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Functional Concept|SIMPLE_SEGMENT|5122,5126|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5122,5140|false|false|false|C0459156|Left bundle branch structure|left bundle branch
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5122,5146|false|false|false|C0023211|Left Bundle-Branch Block|left bundle branch block
Finding|Idea or Concept|SIMPLE_SEGMENT|5122,5146|false|false|false|C2828132|Left Bundle Branch Block Artifact|left bundle branch block
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5122,5146|false|false|false|C0344420||left bundle branch block
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5127,5146|false|false|false|C0006384;C1879286|Bundle-Branch Block;Hereditary bundle branch system defect|bundle branch block
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5134,5140|false|false|false|C1881507|Macromolecular Branch|branch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5141,5146|false|false|false|C1706085|Block Dosage Form|block
Finding|Body Substance|SIMPLE_SEGMENT|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|SIMPLE_SEGMENT|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|SIMPLE_SEGMENT|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Intellectual Product|SIMPLE_SEGMENT|5151,5156|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|5164,5170|false|false|false|C0429103|T wave feature|T wave
Finding|Finding|SIMPLE_SEGMENT|5164,5178|false|false|false|C5780423|T wave changes|T wave changes
Finding|Gene or Genome|SIMPLE_SEGMENT|5166,5170|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5166,5170|false|false|false|C0678544||wave
Finding|Functional Concept|SIMPLE_SEGMENT|5171,5178|false|false|false|C0392747|Changing|changes
Finding|Body Substance|SIMPLE_SEGMENT|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5181,5190|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5191,5195|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5236,5241|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5236,5241|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5242,5245|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5253,5256|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5253,5256|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5253,5256|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5262,5265|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5262,5265|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5262,5265|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5262,5265|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5271,5274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5271,5274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5281,5284|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5281,5284|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5281,5284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5281,5284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5288,5291|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5288,5291|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5288,5291|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5288,5291|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5288,5291|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5297,5301|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5330,5333|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5350,5355|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5350,5355|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5350,5363|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5350,5363|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5350,5363|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5356,5363|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5356,5363|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5356,5363|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5356,5363|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5356,5363|false|false|false|C0337438|Glucose measurement|Glucose
Finding|Intellectual Product|SIMPLE_SEGMENT|5440,5445|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5446,5454|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5446,5461|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5446,5461|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Conceptual Entity|SIMPLE_SEGMENT|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5492,5502|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5504,5508|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5504,5508|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|5504,5508|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|SIMPLE_SEGMENT|5512,5516|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5512,5516|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5512,5516|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5521,5527|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5521,5540|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5521,5540|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5521,5540|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5528,5540|false|false|false|C0232197|Fibrillation|fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|5544,5552|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5544,5552|false|false|false|C1831808|apixaban|apixaban
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5554,5566|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5569,5572|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5569,5572|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|5569,5572|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5569,5572|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5578,5592|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|5578,5592|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5611,5630|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|5611,5630|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|5624,5630|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|5633,5638|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5633,5638|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5633,5638|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5644,5652|false|false|false|C0043144|Wheezing|wheezing
Finding|Idea or Concept|SIMPLE_SEGMENT|5661,5664|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5661,5664|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|5688,5696|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|SIMPLE_SEGMENT|5702,5709|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5702,5709|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5726,5730|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|SIMPLE_SEGMENT|5735,5743|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5735,5743|false|false|false|C0038317|Steroids|steroids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5769,5773|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5769,5773|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|5769,5773|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5769,5786|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|SIMPLE_SEGMENT|5774,5786|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5792,5799|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|5792,5799|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5800,5809|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5800,5809|false|false|false|C1179435|Protein Component|component
Finding|Conceptual Entity|SIMPLE_SEGMENT|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|5841,5848|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|5841,5848|false|false|false|C0039869;C4319827|Thought|thought
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5853,5857|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5853,5857|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|5853,5857|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5853,5870|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|SIMPLE_SEGMENT|5858,5870|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5881,5885|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Organic Chemical|SIMPLE_SEGMENT|5888,5896|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5888,5896|false|false|false|C0038317|Steroids|steroids
Drug|Antibiotic|SIMPLE_SEGMENT|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Finding|Sign or Symptom|SIMPLE_SEGMENT|5917,5925|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|5927,5932|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5927,5932|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5927,5932|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5934,5937|false|false|false|C0013404|Dyspnea|SOB
Finding|Finding|SIMPLE_SEGMENT|5938,5946|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|5938,5946|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Procedure|Health Care Activity|SIMPLE_SEGMENT|5962,5971|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|6000,6004|false|false|false|C5575035|Well (answer to question)|well
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6032,6040|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6032,6040|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6079,6088|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6079,6088|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6079,6088|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6089,6094|false|false|false|C0034991|Rehabilitation therapy|rehab
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6150,6169|false|false|false|C2707305||Shortness of Breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|6150,6169|false|false|false|C0013404|Dyspnea|Shortness of Breath
Finding|Body Substance|SIMPLE_SEGMENT|6163,6169|false|false|false|C0225386|Breath|Breath
Finding|Body Substance|SIMPLE_SEGMENT|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Conceptual Entity|SIMPLE_SEGMENT|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6184,6194|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6195,6199|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6195,6199|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|6195,6199|false|false|false|C1412502|ARCN1 gene|COPD
Procedure|Health Care Activity|SIMPLE_SEGMENT|6212,6221|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|6226,6233|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|6226,6233|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Mental Process|SIMPLE_SEGMENT|6241,6248|false|false|false|C0542559|contextual factors|setting
Drug|Organic Chemical|SIMPLE_SEGMENT|6252,6259|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6252,6259|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Health Care Activity|SIMPLE_SEGMENT|6260,6265|false|false|false|C0441640||taper
Finding|Functional Concept|SIMPLE_SEGMENT|6272,6280|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6272,6280|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|SIMPLE_SEGMENT|6284,6296|false|false|false|C0449450|Presentation|presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|6302,6312|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6302,6317|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|SIMPLE_SEGMENT|6318,6324|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|6318,6324|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6325,6329|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6325,6329|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|6325,6329|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|SIMPLE_SEGMENT|6337,6353|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|6345,6353|false|false|false|C0043144|Wheezing|wheezing
Finding|Intellectual Product|SIMPLE_SEGMENT|6358,6362|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6363,6375|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|6367,6375|false|false|false|C0026649|Movement|movement
Finding|Finding|SIMPLE_SEGMENT|6381,6387|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6381,6387|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|SIMPLE_SEGMENT|6396,6408|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Mental Process|SIMPLE_SEGMENT|6416,6423|false|false|false|C0542559|contextual factors|setting
Finding|Finding|SIMPLE_SEGMENT|6429,6437|false|false|false|C0392756|Reduced|decrease
Drug|Organic Chemical|SIMPLE_SEGMENT|6445,6453|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6445,6453|false|false|false|C0038317|Steroids|steroids
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6476,6485|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6476,6485|false|false|false|C1179435|Protein Component|component
Finding|Conceptual Entity|SIMPLE_SEGMENT|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6489,6496|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|6489,6496|false|false|false|C0860603|Anxiety symptoms|anxiety
Procedure|Health Care Activity|SIMPLE_SEGMENT|6521,6530|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Classification|SIMPLE_SEGMENT|6540,6548|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6540,6548|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6540,6548|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|6540,6552|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6553,6563|false|false|false|C0851162|Infection of musculoskeletal system|infections
Finding|Pathologic Function|SIMPLE_SEGMENT|6553,6563|false|false|false|C3714514|Infection|infections
Finding|Idea or Concept|SIMPLE_SEGMENT|6599,6603|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6599,6603|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6599,6603|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6604,6611|false|false|false|C0905678|Spiriva|spiriva
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6604,6611|false|false|false|C0905678|Spiriva|spiriva
Drug|Organic Chemical|SIMPLE_SEGMENT|6613,6625|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6613,6625|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6613,6625|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|6627,6633|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6627,6633|false|false|false|C0965130|Advair|advair
Drug|Organic Chemical|SIMPLE_SEGMENT|6680,6689|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6680,6689|false|false|false|C0001927|albuterol|albuterol
Finding|Gene or Genome|SIMPLE_SEGMENT|6694,6697|false|false|false|C1422467|CIAO3 gene|prn
Drug|Hormone|SIMPLE_SEGMENT|6702,6712|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|6702,6712|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6702,6712|false|false|false|C0032952|prednisone|prednisone
Procedure|Health Care Activity|SIMPLE_SEGMENT|6750,6755|false|false|false|C0441640||taper
Drug|Antibiotic|SIMPLE_SEGMENT|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|6793,6801|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6793,6801|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6804,6807|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6804,6807|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Conceptual Entity|SIMPLE_SEGMENT|6824,6835|false|false|false|C2986411|Improvement|improvement
Finding|Sign or Symptom|SIMPLE_SEGMENT|6844,6852|false|false|false|C0043144|Wheezing|wheezing
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6869,6877|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6869,6877|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Functional Concept|SIMPLE_SEGMENT|6881,6892|false|false|false|C1514873|Requirement|requirement
Finding|Body Substance|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6968,6977|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|6981,6990|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|6981,6990|false|false|false|C1555324|inpatient encounter|inpatient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6991,7000|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6991,7000|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6991,7000|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6991,7015|false|false|false|C0199529|Pulmonary rehabilitation (procedure)|pulmonary rehabilitation
Finding|Finding|SIMPLE_SEGMENT|7001,7015|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Finding|Functional Concept|SIMPLE_SEGMENT|7001,7015|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7001,7015|false|false|false|C0034991|Rehabilitation therapy|rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7001,7023|false|false|false|C0034991|Rehabilitation therapy|rehabilitation program
Drug|Organic Chemical|SIMPLE_SEGMENT|7016,7023|false|false|false|C2728259|Program|program
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7016,7023|false|false|false|C2728259|Program|program
Finding|Conceptual Entity|SIMPLE_SEGMENT|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Functional Concept|SIMPLE_SEGMENT|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Intellectual Product|SIMPLE_SEGMENT|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7039,7044|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Intellectual Product|SIMPLE_SEGMENT|7098,7102|false|false|false|C1561540|Transaction counts and value totals - week|week
Procedure|Health Care Activity|SIMPLE_SEGMENT|7113,7118|false|false|false|C0441640||taper
Finding|Idea or Concept|SIMPLE_SEGMENT|7150,7158|false|false|false|C0750591|consider|consider
Drug|Organic Chemical|SIMPLE_SEGMENT|7168,7175|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7168,7175|false|false|false|C0591139|Bactrim|bactrim
Finding|Gene or Genome|SIMPLE_SEGMENT|7176,7179|false|false|false|C1418850|PPP4C gene|ppx
Finding|Finding|SIMPLE_SEGMENT|7185,7193|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|SIMPLE_SEGMENT|7185,7193|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7194,7202|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Drug|Organic Chemical|SIMPLE_SEGMENT|7206,7214|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7206,7214|false|false|false|C0038317|Steroids|steroids
Finding|Finding|SIMPLE_SEGMENT|7219,7225|false|false|false|C1299582|Unable|unable
Finding|Classification|SIMPLE_SEGMENT|7270,7280|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7270,7280|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|7287,7291|false|false|false|C1315068|Pulmonary ventilator management|pulm
Finding|Intellectual Product|SIMPLE_SEGMENT|7294,7301|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|7294,7301|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7332,7339|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|7332,7339|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7340,7348|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|7340,7348|false|false|false|C0917801|Sleeplessness|Insomnia
Finding|Idea or Concept|SIMPLE_SEGMENT|7360,7364|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7360,7364|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7360,7364|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7365,7374|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7365,7374|false|false|false|C0024002|lorazepam|lorazepam
Finding|Idea or Concept|SIMPLE_SEGMENT|7376,7384|false|false|false|C0750591|consider|Consider
Finding|Classification|SIMPLE_SEGMENT|7406,7416|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7406,7416|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7421,7427|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7421,7440|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7421,7440|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7421,7440|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7428,7440|false|false|false|C0232197|Fibrillation|Fibrillation
Drug|Organic Chemical|SIMPLE_SEGMENT|7452,7456|false|false|false|C1601858|Dilt|dilt
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7452,7456|false|false|false|C1601858|Dilt|dilt
Event|Activity|SIMPLE_SEGMENT|7461,7465|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|SIMPLE_SEGMENT|7461,7465|false|false|false|C1549480|Amount type - Rate|rate
Finding|Functional Concept|SIMPLE_SEGMENT|7461,7473|false|false|false|C0489879|rate control|rate control
Drug|Organic Chemical|SIMPLE_SEGMENT|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|SIMPLE_SEGMENT|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|SIMPLE_SEGMENT|7479,7487|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7479,7487|false|false|false|C1831808|apixaban|apixaban
Finding|Finding|SIMPLE_SEGMENT|7492,7507|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|7492,7507|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7492,7507|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7511,7523|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Idea or Concept|SIMPLE_SEGMENT|7535,7539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7535,7539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7535,7539|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7540,7545|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7540,7545|false|false|false|C0590690|Imdur|imdur
Drug|Organic Chemical|SIMPLE_SEGMENT|7547,7566|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7547,7566|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|7573,7582|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7573,7582|false|false|false|C0012373|diltiazem|diltiazem
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7586,7589|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7586,7589|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|7586,7589|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7586,7589|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7591,7598|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|7591,7598|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7591,7614|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|7591,7614|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7591,7614|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|7591,7614|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7599,7614|false|false|false|C0007430|Catheterization|catheterization
Finding|Idea or Concept|SIMPLE_SEGMENT|7630,7638|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7630,7641|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|SIMPLE_SEGMENT|7643,7654|false|false|false|C0750502|Significant|significant
Finding|Pathologic Function|SIMPLE_SEGMENT|7655,7663|false|false|false|C1261287|Stenosis|stenosis
Procedure|Health Care Activity|SIMPLE_SEGMENT|7679,7683|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7679,7683|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7732,7743|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7737,7743|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|7744,7757|false|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|7744,7757|false|false|false|C0000769|teratologic|abnormalities
Finding|Idea or Concept|SIMPLE_SEGMENT|7770,7774|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7770,7774|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7770,7774|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7775,7782|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7775,7782|false|false|false|C0004057|aspirin|aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|7787,7799|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7787,7799|false|false|false|C0286651|atorvastatin|atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7803,7809|false|false|false|C0002871|Anemia|Anemia
Finding|Idea or Concept|SIMPLE_SEGMENT|7821,7825|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7821,7825|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7821,7825|false|false|false|C1553498|home health encounter|home
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7826,7830|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7826,7842|false|false|false|C0721124|Iron Supplement|iron supplements
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7826,7842|false|false|false|C0721124|Iron Supplement|iron supplements
Finding|Idea or Concept|SIMPLE_SEGMENT|7845,7857|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Idea or Concept|SIMPLE_SEGMENT|7905,7914|false|false|false|C0549178|Continuous|continued
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7915,7919|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7915,7919|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|7915,7919|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Antibiotic|SIMPLE_SEGMENT|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Finding|Finding|SIMPLE_SEGMENT|8015,8023|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|SIMPLE_SEGMENT|8015,8023|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Drug|Hormone|SIMPLE_SEGMENT|8024,8034|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|8024,8034|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8024,8034|false|false|false|C0032952|prednisone|prednisone
Procedure|Health Care Activity|SIMPLE_SEGMENT|8035,8040|false|false|false|C0441640||taper
Drug|Hormone|SIMPLE_SEGMENT|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Finding|Functional Concept|SIMPLE_SEGMENT|8073,8079|false|false|false|C1706059|Finish - dosing instruction imperative|finish
Procedure|Health Care Activity|SIMPLE_SEGMENT|8101,8106|false|false|false|C0441640||taper
Finding|Idea or Concept|SIMPLE_SEGMENT|8147,8150|false|false|false|C1548556|Etc.|etc
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8175,8178|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8175,8178|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8175,8190|false|false|false|C0747314|pcp prophylaxis|PCP prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8179,8190|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Finding|SIMPLE_SEGMENT|8203,8209|false|false|false|C1299582|Unable|unable
Finding|Finding|SIMPLE_SEGMENT|8213,8217|false|false|false|C0043084|Weaning|wean
Drug|Hormone|SIMPLE_SEGMENT|8219,8229|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|8219,8229|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8219,8229|false|false|false|C0032952|prednisone|prednisone
Finding|Sign or Symptom|SIMPLE_SEGMENT|8264,8267|false|false|false|C0013404|Dyspnea|SOB
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8280,8287|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|8280,8287|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8288,8297|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8288,8297|false|false|false|C1179435|Protein Component|component
Finding|Conceptual Entity|SIMPLE_SEGMENT|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8326,8330|false|false|false|C0360105;C2911696|Selective Serotonin Reuptake Inhibitors;Serotonin Reuptake Inhibitor [EPC]|SSRI
Finding|Functional Concept|SIMPLE_SEGMENT|8331,8345|false|false|false|C0332287|In addition to|in addition to
Finding|Functional Concept|SIMPLE_SEGMENT|8334,8342|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Finding|Idea or Concept|SIMPLE_SEGMENT|8346,8350|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8346,8350|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8346,8350|false|false|false|C1553498|home health encounter|home
Event|Activity|SIMPLE_SEGMENT|8380,8387|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8380,8387|false|false|false|C0392367|Physical contact|CONTACT
Event|Occupational Activity|SIMPLE_SEGMENT|8394,8398|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|8394,8398|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Occupational Activity|SIMPLE_SEGMENT|8401,8405|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|8401,8405|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|SIMPLE_SEGMENT|8401,8412|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8406,8412|false|false|false|C5889824||STATUS
Finding|Idea or Concept|SIMPLE_SEGMENT|8406,8412|false|false|false|C1546481|What subject filter - Status|STATUS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8427,8430|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8427,8430|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Procedure|Health Care Activity|SIMPLE_SEGMENT|8445,8454|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8473,8483|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8473,8483|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8473,8488|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|8484,8488|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|8505,8513|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8505,8513|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8518,8531|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8518,8531|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8518,8531|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|8546,8549|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8550,8554|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|8550,8554|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8550,8554|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8559,8567|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8559,8567|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8576,8579|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8576,8579|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8576,8579|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8576,8579|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8584,8591|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8584,8591|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8611,8623|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8611,8623|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8641,8650|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8641,8650|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|8651,8659|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8651,8659|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8660,8667|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|8660,8667|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8660,8667|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8678,8681|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8678,8681|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8678,8681|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8678,8681|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8686,8694|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8686,8694|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|8686,8701|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8686,8701|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8695,8701|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8695,8701|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8712,8715|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8712,8715|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8712,8715|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8712,8715|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8720,8731|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8720,8731|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|8735,8740|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8750,8754|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|8750,8754|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8755,8764|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8760,8764|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8760,8764|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8765,8768|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8765,8768|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8765,8768|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8765,8768|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8773,8780|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8773,8788|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8773,8788|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|8809,8820|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8809,8820|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|8809,8831|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8809,8831|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|8821,8831|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8832,8837|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|8832,8837|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|8832,8837|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Gene or Genome|SIMPLE_SEGMENT|8854,8857|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8858,8867|false|false|false|C1717415||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|8858,8867|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|8873,8892|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8873,8892|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|8913,8923|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8913,8923|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8913,8935|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8913,8935|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|SIMPLE_SEGMENT|8937,8945|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8937,8945|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8946,8953|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|8946,8953|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8946,8953|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|8976,8987|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8976,8987|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|8995,9000|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9010,9014|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|9010,9014|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9015,9024|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9020,9024|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9020,9024|false|false|false|C5848506||EYES
Drug|Organic Chemical|SIMPLE_SEGMENT|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9050,9053|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Hormone|SIMPLE_SEGMENT|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|9099,9109|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9099,9109|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|9131,9143|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9131,9143|false|false|false|C0039771|theophylline|Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9131,9143|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|9131,9146|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9131,9146|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9157,9160|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9157,9160|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9157,9160|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9157,9160|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9166,9176|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9166,9176|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|9166,9184|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9166,9184|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9177,9184|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9177,9184|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|9187,9190|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9187,9190|false|false|false|C0006935|capsule (pharmacologic)|CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|9187,9190|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9187,9190|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|9205,9216|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9205,9216|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|9205,9224|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9205,9224|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9217,9224|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9217,9224|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|9225,9228|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|9225,9228|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|SIMPLE_SEGMENT|9231,9234|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9231,9234|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|9242,9245|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|9246,9254|false|false|false|C0043144|Wheezing|Wheezing
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|SIMPLE_SEGMENT|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|SIMPLE_SEGMENT|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|SIMPLE_SEGMENT|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|SIMPLE_SEGMENT|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|SIMPLE_SEGMENT|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|SIMPLE_SEGMENT|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|SIMPLE_SEGMENT|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|9264,9269|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|9264,9269|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|SIMPLE_SEGMENT|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|SIMPLE_SEGMENT|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9276,9283|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|9276,9283|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9276,9283|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9285,9289|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9285,9289|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9285,9289|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9285,9289|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9290,9293|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9290,9293|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9290,9293|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9290,9293|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9299,9309|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9299,9309|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9310,9319|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|9321,9328|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9321,9328|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|9321,9336|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9321,9336|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9329,9336|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9329,9336|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9329,9336|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9370,9374|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9370,9374|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9370,9374|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9370,9374|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|9386,9395|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9386,9395|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9386,9403|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9386,9403|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|9421,9431|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|9421,9431|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Drug|Organic Chemical|SIMPLE_SEGMENT|9441,9452|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9441,9452|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9441,9463|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9441,9470|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9441,9470|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|9453,9463|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9453,9463|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Finding|Functional Concept|SIMPLE_SEGMENT|9483,9486|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9490,9493|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9490,9493|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9490,9493|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9490,9493|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9499,9508|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9499,9508|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|9523,9526|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9527,9534|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9527,9534|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Organic Chemical|SIMPLE_SEGMENT|9540,9551|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9540,9551|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|SIMPLE_SEGMENT|9566,9569|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|9570,9575|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9570,9575|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|9570,9575|false|false|false|C0010200|Coughing|cough
Finding|Body Substance|SIMPLE_SEGMENT|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9580,9589|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9580,9601|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9590,9601|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9590,9601|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9590,9601|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9606,9619|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9606,9619|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9606,9619|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|9634,9637|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9638,9642|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|9638,9642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9638,9642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9647,9656|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9647,9656|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|9647,9664|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9647,9664|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|9682,9692|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|9682,9692|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Drug|Organic Chemical|SIMPLE_SEGMENT|9701,9709|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9701,9709|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9718,9721|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9718,9721|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9718,9721|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9718,9721|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9726,9733|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9726,9733|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9753,9765|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9753,9765|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9783,9792|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9783,9792|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|SIMPLE_SEGMENT|9793,9801|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9793,9801|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9802,9809|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|9802,9809|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9802,9809|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9820,9823|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9820,9823|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9820,9823|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9820,9823|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9828,9836|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9828,9836|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|9828,9843|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9828,9843|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9837,9843|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9837,9843|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9854,9857|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9854,9857|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9854,9857|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9854,9857|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9862,9873|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9862,9873|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|SIMPLE_SEGMENT|9877,9882|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9892,9896|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|9892,9896|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9897,9906|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9902,9906|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9902,9906|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9907,9910|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9907,9910|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9907,9910|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9907,9910|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9915,9922|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9915,9930|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9915,9930|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Organic Chemical|SIMPLE_SEGMENT|9952,9963|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9952,9963|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9952,9974|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9952,9974|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|9964,9974|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9975,9980|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|SIMPLE_SEGMENT|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|SIMPLE_SEGMENT|9975,9980|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|SIMPLE_SEGMENT|9975,9980|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Gene or Genome|SIMPLE_SEGMENT|9997,10000|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10001,10010|false|false|false|C1717415||allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|10001,10010|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|10016,10027|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10016,10027|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10016,10038|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|10016,10045|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10016,10045|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|SIMPLE_SEGMENT|10028,10038|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10028,10038|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|SIMPLE_SEGMENT|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Finding|Functional Concept|SIMPLE_SEGMENT|10058,10061|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10065,10068|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10065,10068|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10065,10068|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10065,10068|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10074,10085|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10074,10085|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|SIMPLE_SEGMENT|10100,10103|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|10104,10109|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10104,10109|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|10104,10109|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|SIMPLE_SEGMENT|10115,10134|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10115,10134|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|10155,10165|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10155,10165|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|10155,10177|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10155,10177|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|SIMPLE_SEGMENT|10179,10187|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10179,10187|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10188,10195|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10188,10195|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10188,10195|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|10218,10229|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10218,10229|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|SIMPLE_SEGMENT|10237,10242|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10252,10256|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|10252,10256|false|false|false|C1705648|Dropping|DROP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10257,10266|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10262,10266|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10262,10266|false|false|false|C5848506||EYES
Drug|Organic Chemical|SIMPLE_SEGMENT|10276,10285|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10276,10285|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|10300,10303|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10304,10311|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|10304,10311|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Organic Chemical|SIMPLE_SEGMENT|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10333,10336|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|10351,10361|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10351,10361|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|10383,10395|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10383,10395|false|false|false|C0039771|theophylline|Theophylline
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10383,10395|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|SIMPLE_SEGMENT|10383,10398|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10383,10398|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10409,10412|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10409,10412|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10409,10412|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10409,10412|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10418,10428|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10418,10428|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Organic Chemical|SIMPLE_SEGMENT|10418,10436|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10418,10436|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10429,10436|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10429,10436|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|10439,10442|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10439,10442|false|false|false|C0006935|capsule (pharmacologic)|CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|10439,10442|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10439,10442|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|10457,10467|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10457,10467|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10468,10477|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|10479,10486|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10479,10486|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|SIMPLE_SEGMENT|10479,10494|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10479,10494|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10487,10494|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10487,10494|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10487,10494|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|SIMPLE_SEGMENT|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10528,10532|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10528,10532|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|10528,10532|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|10528,10532|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|SIMPLE_SEGMENT|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|SIMPLE_SEGMENT|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|SIMPLE_SEGMENT|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|SIMPLE_SEGMENT|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|SIMPLE_SEGMENT|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|SIMPLE_SEGMENT|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|SIMPLE_SEGMENT|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|10548,10553|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|10548,10553|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|SIMPLE_SEGMENT|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|SIMPLE_SEGMENT|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10560,10567|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10560,10567|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10560,10567|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10569,10573|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10569,10573|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|10569,10573|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|10569,10573|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10574,10577|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10574,10577|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10574,10577|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10574,10577|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10583,10594|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10583,10594|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|10583,10602|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10583,10602|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10595,10602|false|false|false|C0006222|Bromides|Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10595,10602|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|10603,10606|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|10603,10606|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|SIMPLE_SEGMENT|10609,10612|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|10609,10612|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|10620,10623|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|10624,10632|false|false|false|C0043144|Wheezing|Wheezing
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10638,10646|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|10638,10646|false|false|false|C0028040|nicotine|Nicotine
Drug|Clinical Drug|SIMPLE_SEGMENT|10638,10652|false|false|false|C0358855|Nicotine Transdermal Patch|Nicotine Patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10647,10652|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|SIMPLE_SEGMENT|10647,10652|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Antibiotic|SIMPLE_SEGMENT|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10700,10708|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Drug|Hormone|SIMPLE_SEGMENT|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|SIMPLE_SEGMENT|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10768,10776|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Procedure|Health Care Activity|SIMPLE_SEGMENT|10802,10809|false|false|false|C0441640||Tapered
Finding|Body Substance|SIMPLE_SEGMENT|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10826,10835|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10826,10847|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10826,10847|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10836,10847|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10836,10847|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|10849,10862|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|10858,10862|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|10858,10862|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|10858,10862|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|10865,10873|false|false|false|C4695111|ADMIN.FACILITY|Facility
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10885,10894|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10885,10894|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10885,10894|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10885,10894|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10905,10909|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10905,10909|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|10905,10909|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10905,10922|false|false|false|C0740304|COPD exacerbation|COPD Exacerbation
Finding|Finding|SIMPLE_SEGMENT|10910,10922|false|false|false|C4086268|Exacerbation|Exacerbation
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10924,10933|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|SIMPLE_SEGMENT|10924,10933|false|false|false|C1522484|metastatic qualifier|SECONDARY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10935,10939|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10935,10939|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10940,10947|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|10940,10947|false|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10948,10951|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10952,10955|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10952,10955|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|10952,10955|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|10952,10955|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Body Substance|SIMPLE_SEGMENT|10959,10968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10959,10968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10959,10968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10959,10968|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10969,10978|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10969,10978|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10969,10978|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10980,10986|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10980,10993|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10980,10993|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10987,10993|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10987,10993|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10995,11000|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|11005,11013|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11015,11037|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|11015,11037|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|11024,11037|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|11024,11037|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11039,11044|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|11039,11044|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11039,11044|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|11049,11060|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|11062,11070|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11062,11070|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|11062,11070|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11071,11077|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|11071,11077|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|11079,11089|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Social Behavior|SIMPLE_SEGMENT|11101,11111|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11115,11118|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|11115,11118|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|SIMPLE_SEGMENT|11115,11118|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11115,11118|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Body Substance|SIMPLE_SEGMENT|11141,11150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11141,11150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11141,11150|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11141,11150|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11141,11163|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11141,11163|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|11141,11163|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11151,11163|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11151,11163|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|11165,11169|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11226,11245|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|11226,11245|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|11239,11245|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|11250,11258|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|SIMPLE_SEGMENT|11259,11266|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|11262,11266|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11262,11266|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11262,11266|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11292,11301|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11326,11330|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11326,11330|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|11326,11330|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11326,11343|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|SIMPLE_SEGMENT|11331,11343|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Idea or Concept|SIMPLE_SEGMENT|11376,11382|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Finding|SIMPLE_SEGMENT|11388,11396|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|11388,11396|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|11388,11396|false|false|false|C0031809|Physical Examination|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|11455,11465|false|false|false|C1698490|short stay encounter|short stay
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11469,11478|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11469,11478|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|11469,11478|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Idea or Concept|SIMPLE_SEGMENT|11497,11501|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11497,11501|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11497,11501|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11518,11527|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|11518,11527|false|false|false|C1160636|respiratory system process|breathing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11551,11555|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|SIMPLE_SEGMENT|11551,11555|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11559,11564|false|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Classification|SIMPLE_SEGMENT|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|11621,11625|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Intellectual Product|SIMPLE_SEGMENT|11643,11651|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11643,11651|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11659,11663|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|11659,11663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11659,11663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11659,11666|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|SIMPLE_SEGMENT|11689,11697|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11698,11710|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11698,11710|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

