CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Corgard|Drug|false|false||Corgard
null|Corgard|Drug|false|false||Corgardnull|Vasotec|Drug|false|false||Vasotec
null|Vasotec|Drug|false|false||Vasotecnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Dyspnea on exertion|Finding|false|false||Dyspnea on Exertionnull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Exertion|Finding|false|false||Exertionnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Referral category - Outpatient|Finding|false|false||OUTPATIENT
null|Patient Class - Outpatient|Finding|false|false||OUTPATIENTnull|Outpatients|Subject|false|false||OUTPATIENTnull|Cardiologists|Subject|false|false||CARDIOLOGISTnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Congestive heart failure|Disorder|false|false|C0262212|CHFnull|Choroidal fissure|Anatomy|false|false|C0018802|CHFnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Chief complaint (finding)|Finding|false|false||CHIEF COMPLAINTnull|Complaint (finding)|Finding|false|false||COMPLAINTnull|null|Attribute|false|false||COMPLAINTnull|Dyspnea on exertion|Finding|false|false||Dyspnea on Exertionnull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Exertion|Finding|false|false||Exertionnull|Medical History|Finding|false|false||HISTORY OFnull|History of present illness (finding)|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|Medical History|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|Presentation|Finding|true|false||PRESENTINGnull|Illness (finding)|Finding|false|false||ILLNESSnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Tricuspid regurgitation, moderate|Finding|false|false||moderate tricuspid regurgitationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Tricuspid Valve Insufficiency|Disorder|false|false||tricuspid regurgitationnull|Tricuspid|Modifier|false|false||tricuspidnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Ventricular Dysfunction|Finding|false|false|C0018827|ventricular dysfunctionnull|Heart Ventricle|Anatomy|false|false|C3887505;C0031847;C0277785;C3887504;C0242973|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false|C0018827|dysfunction
null|physiopathological|Finding|false|false|C0018827|dysfunction
null|Functional disorder|Finding|false|false|C0018827|dysfunctionnull|Moderate pulmonary hypertension|Finding|false|false|C0024109|moderate pulmonary hypertensionnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Pulmonary Hypertension|Finding|false|false|C0024109|pulmonary hypertensionnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C5395246;C0020542;C4522268;C0020538;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Hypertensive disease|Disorder|false|false|C0024109|hypertensionnull|Paroxysmal atrial fibrillation|Disorder|false|false|C0018792|paroxysmal atrial fibrillationnull|Paroxysmal|Time|false|false||paroxysmalnull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0344434;C0232197;C0004238;C0235480;C2926591|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0022658;C1552824;C0496927;C0496892;C0812426;C4554465;C0869841;C0012634|kidney
null|Both kidneys|Anatomy|false|false|C0022658;C1552824;C0496927;C0496892;C0812426;C4554465;C0869841;C0012634|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|BaseLine dental cement|Drug|false|false||Baselinenull|baseline - TableCellVerticalAlign|Finding|false|false|C0227665;C0022646|Baselinenull|Baseline|LabModifier|false|false||Baselinenull|Cerebrovascular Disorders|Disorder|false|false||cerebrovascular diseasenull|Cerebrovascular|Modifier|false|false||cerebrovascularnull|Disease|Disorder|false|false||diseasenull|Metastatic melanoma|Disorder|false|false||metastatic melanomanull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Melanoma of Unknown Primary|Disorder|false|false||melanoma of unknown primarynull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Cell Cycle Checkpoints|Finding|false|false||checkpointnull|Inhibitor|Drug|false|false||inhibitornull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Dyspnea on exertion|Finding|false|false||DOEnull|Department of Energy|Subject|false|false||DOEnull|Adult female goat|Entity|false|false||DOEnull|Diuresis|Finding|false|false||diuresisnull|Most recent outpatient|Finding|false|false||most recent outpatientnull|Most Recent|Time|false|false||most recentnull|Recent|Time|false|false||recentnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Congestive heart failure|Disorder|false|false|C0262212|CHFnull|Choroidal fissure|Anatomy|false|false|C0018802|CHFnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Drug|false|false|C1166663|carnull|Carney Complex|Disorder|false|false|C1166663|carnull|Car - Mode of Arrival Code|Finding|false|false|C1166663|car
null|Chimeric antigen receptor|Finding|false|false|C1166663|car
null|CASR wt Allele|Finding|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Finding|false|false|C1166663|car
null|CXADR wt Allele|Finding|false|false|C1166663|car
null|CXADR gene|Finding|false|false|C1166663|car
null|PRKAR1A wt Allele|Finding|false|false|C1166663|car
null|CXADRP1 gene|Finding|false|false|C1166663|car
null|NR1I3 gene|Finding|false|false|C1166663|car
null|SPG7 gene|Finding|false|false|C1166663|car
null|TRIM13 wt Allele|Finding|false|false|C1166663|car
null|Caronte Gene|Finding|false|false|C1166663|car
null|SPG7 wt Allele|Finding|false|false|C1166663|car
null|NR1I3 wt Allele|Finding|false|false|C1166663|carnull|actomyosin contractile ring|Anatomy|false|false|C3540475;C1547285;C3273602;C4039583;C1413828;C3811749;C2239319;C1858724;C1417827;C5890847;C1420354;C5960871;C1706434;C5890846;C2024878;C0013404;C0406810;C0231807;C3539542;C4039583;C5890846|carnull|Automobiles|Device|false|false||carnull|Car <Caridae>|Entity|false|false||car
null|Carib language|Entity|false|false||carnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Cardiologists|Subject|false|false||Cardiologistnull|Increased fatigue|Finding|false|false||increased fatiguenull|Fatigue|Finding|false|false||fatiguenull|Dyspnea on exertion|Finding|false|false|C1166663|exertional dyspneanull|exercise induced|Finding|false|false||exertionalnull|null|Finding|false|false|C1166663|dyspnea
null|Dyspnea|Finding|false|false|C1166663|dyspneanull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|null|Time|false|false||priornull|Low-Dose Treatment|Procedure|false|false||low-dosenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Entresto|Drug|false|false||Entresto
null|Entresto|Drug|false|false||Entrestonull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Lightheadedness|Finding|false|false||lightheadednessnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Patient Outcome - Worsening|Finding|false|false|C0022646|worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0042075;C1546960|renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Concern|Finding|false|false||concernnull|Myocarditis|Disorder|false|false||myocarditisnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Cell Cycle Checkpoints|Finding|false|false||checkpointnull|Inhibitor|Drug|false|false||inhibitornull|Neoplasms|Disorder|false|false||Oncologynull|oncology services|Procedure|false|false||Oncologynull|oncology (field)|Title|false|false||Oncologynull|Team|Subject|false|false||teamnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Somewhat|Finding|false|false||somewhatnull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|null|Attribute|false|false|C0018787|Cardiac biomarkers
null|Cardiac biomarkers|Attribute|false|false|C0018787|Cardiac biomarkersnull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C2735101;C2735102;C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Biological Markers|Attribute|false|false||biomarkersnull|pro-brain natriuretic peptide (1-76)|Drug|false|false||NTproBNP
null|pro-brain natriuretic peptide (1-76)|Drug|false|false||NTproBNPnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|Unexpected|Finding|true|false||unexpectednull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Decompensated|Modifier|false|false||decompensatednull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0812426;C4554465;C0869841;C0496927;C0496892;C0022658;C1561643;C0012634|kidney
null|Both kidneys|Anatomy|false|false|C0812426;C4554465;C0869841;C0496927;C0496892;C0022658;C1561643;C0012634|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|Immunotherapy [APC]|Drug|false|false||immunotherapynull|Immunotherapy|Procedure|false|false||immunotherapynull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Improvement|Finding|false|false||improvementnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumabnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Intravenous Route of Administration|Finding|false|false||intravenousnull|Intravenous|Modifier|false|false||intravenousnull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|More|LabModifier|false|false||morenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||dailynull|Daily|Time|false|false||dailynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Daily|Time|false|false||dailynull|Troponin|Drug|false|false||Troponin
null|Troponin|Drug|false|false||Troponinnull|Troponin measurement|Procedure|false|false||Troponinnull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0042075|renalnull|Insufficiency|Finding|false|false||insufficiencynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Hyperkalemia|Finding|false|false||hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||hyperkalemianull|Potassium supplementation (product)|Drug|false|false||potassium supplementationnull|Potassium supplement therapy|Procedure|false|false||potassium supplementationnull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Dietary Supplementation|Procedure|false|false||supplementationnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Encounter Referral Source - emergency room|Finding|false|false||Emergency roomnull|Accident and Emergency department|Device|false|false||Emergency roomnull|Accident and Emergency department|Entity|false|false||Emergency roomnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Scalp laceration|Disorder|false|false|C0036270|scalp lacerationnull|Scalp structure|Anatomy|false|false|C0043246;C0240937|scalpnull|Laceration|Disorder|false|false|C0036270|lacerationnull|CAT scan of head|Procedure|false|false|C0018670;C0152336;C0460004;C0027530;C3159206|CT headnull|null|Attribute|false|false|C0018670;C0152336|CT headnull|Head and neck structure|Anatomy|false|false|C0876917;C0202691;C0812434;C0684335;C0362076|head and necknull|Problems with head|Disorder|false|false|C0027530;C3159206;C0018670;C0152336;C0460004|headnull|Procedure on head|Procedure|false|false|C0460004;C0027530;C3159206;C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0202691;C0881943;C0362076;C0876917|head
null|Head|Anatomy|false|false|C0202691;C0881943;C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Passive joint movement of neck (finding)|Finding|false|false|C0460004;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0460004;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0362076;C0202691;C0812434;C0684335;C0876917|neck
null|Neck|Anatomy|false|false|C0362076;C0202691;C0812434;C0684335;C0876917|necknull|null|Modifier|false|false||unremarkablenull|Morning|Time|false|false||morningnull|Visit|Finding|false|false||visitnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Recent|Time|false|false||recentlynull|Visit User Code - Home|Finding|false|false|C0222045|home
null|Address type - Home|Finding|false|false|C0222045|homenull|home health encounter|Procedure|false|false|C0222045|homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Scale, LOINC Axis 5|Finding|false|false|C0222045|scale
null|Base Number|Finding|false|false|C0222045|scale
null|Scale - rank|Finding|false|false|C0222045|scalenull|Integumentary scale|Anatomy|false|false|C0349674;C2981742;C1522412;C1553498;C1549632;C1548341;C1947916|scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false|C0222045|scalenull|Decrease in appetite|Finding|false|false||decreased appetitenull|Desire for food|Finding|false|false||appetitenull|Different|Modifier|false|false||differentnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Current (present time)|Time|false|false||currentlynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Low sodium diet|Procedure|false|false||low sodium dietnull|Sodium decreased|Finding|false|false||low sodiumnull|Low sodium diet|Procedure|false|false||low sodiumnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Sodium diet|Procedure|false|false||sodium dietnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Much|Finding|false|false||muchnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Eyeglasses|Device|false|false||glassesnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Juice|Drug|false|false||juicenull|Daily|Time|false|false||dailynull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Daily|Time|false|false||dailynull|Daily|Time|false|false||dailynull|Several days|Finding|false|false||several daysnull|Several|LabModifier|false|false||severalnull|day|Time|false|false||daysnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Frequently|Time|false|false||frequentlynull|tamsulosin|Drug|false|false||tamsulosin
null|tamsulosin|Drug|false|false||tamsulosinnull|Several days|Finding|false|false||several daysnull|Several|LabModifier|false|false||severalnull|day|Time|false|false||daysnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|Step (specific stage)|Finding|false|false||stepsnull|STEPS to Enhance Physical Activity|Procedure|false|false||stepsnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Diuresis|Finding|false|false||diuresisnull|Floor (anatomic)|Anatomy|false|false|C0262926;C1705255;C0019665;C0262512;C2004062|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|History of present illness (finding)|Finding|false|false|C3714591|history
null|History of previous events|Finding|false|false|C3714591|history
null|Historical aspects qualifier|Finding|false|false|C3714591|history
null|Medical History|Finding|false|false|C3714591|history
null|Concept History|Finding|false|false|C3714591|historynull|History|Subject|false|false||historynull|Dyspnea|Finding|false|false||SOBnull|Progressive|Finding|false|false||progressivenull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|MOSTLY|Finding|false|false||Mostlynull|null|LabModifier|false|false||Mostlynull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Slow|Modifier|false|false||slowlynull|Anorexia|Disorder|false|false||lack of appetitenull|Loss of appetite (finding)|Finding|false|false||lack of appetitenull|Lacking|Modifier|false|false||lacknull|Desire for food|Finding|false|false||appetitenull|home health encounter|Procedure|false|false||home healthnull|Home health care specialty|Title|false|false||home healthnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Health|Finding|false|false||healthnull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Daily|Time|false|false||everydaynull|Maxillary right lateral incisor mesial prosthesis|Device|false|false||7pmnull|VISCERAL LEIOMYOPATHY, AFRICAN DEGENERATIVE|Disorder|false|false||ADLnull|Activity of daily living (function)|Finding|false|false||ADL
null|SGCA gene|Finding|false|false||ADL
null|SGCA wt Allele|Finding|false|false||ADLnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C0489633;C1314974;C0449913;C1552617;C0282443;C0699752|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Review of systems (procedure)|Procedure|false|false|C0018787|review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false|C0018787|review ofnull|Review (Publication Type)|Finding|false|false|C0018787|review
null|Act Class - review|Finding|false|false|C0018787|reviewnull|System|Finding|false|false|C0018787|systemsnull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||paroxysmal nocturnal dyspneanull|Paroxysmal|Time|false|false||paroxysmalnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Palpitations|Finding|false|false||palpitationsnull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Presyncope|Finding|false|false||presyncopenull|Reactive Oxygen Species|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|Reactive Oxygen Species|Drug|false|false|C0262327|ROSnull|ROS1 wt Allele|Finding|false|false|C0262327|ROS
null|ROS1 gene|Finding|false|false|C0262327|ROSnull|Review of systems (procedure)|Procedure|false|false|C0262327|ROSnull|rostral sulcus|Anatomy|false|false|C0289313;C0162772;C0489633;C2699077;C0205160;C1513916;C0812281;C1709820|ROSnull|Rh Negative Blood Group|Finding|false|false|C0262327|negative
null|Negative|Finding|false|false|C0262327|negative
null|Negative Finding|Finding|false|false|C0262327|negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Bilateral|Modifier|false|false||BILATERALnull|Moderate - Severity of Illness Code|Finding|false|false||MODERATE
null|Moderate|Finding|false|false||MODERATEnull|Moderate (severity modifier)|Modifier|false|false||MODERATE
null|Moderate - Allergy Severity|Modifier|false|false||MODERATE
null|Moderation|Modifier|false|false||MODERATEnull|carotid disease|Disorder|false|false|C0007272|CAROTID DISEASEnull|Carotid Arteries|Anatomy|false|false|C0012634;C0741975|CAROTIDnull|Disease|Disorder|false|false|C0007272|DISEASEnull|Congestive|Modifier|false|false||CONGESTIVEnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Coronary Artery Disease|Disorder|false|false|C0205042;C0226004;C0003842;C0018787|CORONARY ARTERY DISEASE
null|Coronary Arteriosclerosis|Disorder|false|false|C0205042;C0226004;C0003842;C0018787|CORONARY ARTERY DISEASEnull|Coronary artery|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|CORONARY ARTERYnull|Heart|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Arteriopathic disease|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|ARTERY DISEASEnull|Arterial system|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|ARTERY
null|Arteries|Anatomy|false|false|C0852949;C0012634;C1956346;C0010054|ARTERYnull|Disease|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|DISEASEnull|Gastroesophageal reflux disease|Disorder|false|false|C0744316|GASTROESOPHAGEAL REFLUXnull|Infantile Gastroesophageal Reflux|Finding|false|false|C0744316|GASTROESOPHAGEAL REFLUX
null|Acid reflux|Finding|false|false|C0744316|GASTROESOPHAGEAL REFLUXnull|gastroesophageal|Anatomy|false|false|C0017168;C0232483;C3813607;C4317146|GASTROESOPHAGEALnull|Reflux|Finding|false|false|C0744316|REFLUXnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Severe - Severity of Illness Code|Finding|false|false||SEVERE
null|Intensity and Distress 5|Finding|false|false||SEVERE
null|Severe - Triage Code|Finding|false|false||SEVERE
null|Severe (severity modifier)|Finding|false|false||SEVERE
null|Allergy Severity - Severe|Finding|false|false||SEVEREnull|Pulmonary Emphysema|Disorder|false|false||EMPHYSEMAnull|Pathological accumulation of air in tissues|Finding|false|false||EMPHYSEMAnull|Pulmonary Hypertension|Finding|false|false|C0024109|PULMONARY HYPERTENSIONnull|Pulmonary (intended site)|Finding|false|false|C0024109|PULMONARYnull|Lung|Anatomy|false|false|C4522268;C0020542;C2707265;C0020538|PULMONARYnull|null|Attribute|false|false|C0024109|PULMONARYnull|Pulmonary (qualifier value)|Modifier|false|false||PULMONARYnull|Hypertensive disease|Disorder|false|false|C0024109|HYPERTENSIONnull|Right bundle branch block|Disorder|false|false|C0225916|RIGHT BUNDLE BRANCH BLOCKnull|null|Finding|false|false|C0225916|RIGHT BUNDLE BRANCH BLOCKnull|Structure of right branch of atrioventricular bundle|Anatomy|false|false|C1706085;C0028778;C0332206;C1533157;C1879286;C0006384;C1881507;C1552823;C0344421;C0085615|RIGHT BUNDLE BRANCHnull|Table Cell Horizontal Align - right|Finding|false|false|C0225916|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Bundle-Branch Block|Disorder|false|false|C0225916|BUNDLE BRANCH BLOCK
null|Hereditary bundle branch system defect|Disorder|false|false|C0225916|BUNDLE BRANCH BLOCKnull|Macromolecular Branch|Drug|false|false|C0225916|BRANCHnull|Branch of|Modifier|false|false||BRANCHnull|Block Dosage Form|Drug|false|false|C0225916|BLOCKnull|Fixed Block|Finding|false|false|C0225916|BLOCK
null|Obstruction|Finding|false|false|C0225916|BLOCK
null|Blocking|Finding|false|false|C0225916|BLOCKnull|Geographic Block|Entity|false|false||BLOCKnull|Block (unit of presentation)|LabModifier|false|false||BLOCK
null|Block Dosing Unit|LabModifier|false|false||BLOCK
null|Block (unit of measure)|LabModifier|false|false||BLOCKnull|Benign Prostatic Hyperplasia|Finding|false|false|C0033572|BENIGN PROSTATIC HYPERTROPHYnull|Benign|Modifier|false|false||BENIGNnull|Prostatic Hypertrophy|Disorder|false|false|C0033572|PROSTATIC HYPERTROPHYnull|Benign Prostatic Hyperplasia|Finding|false|false|C0033572|PROSTATIC HYPERTROPHY
null|Prostatic Hyperplasia|Finding|false|false|C0033572|PROSTATIC HYPERTROPHYnull|Prostate|Anatomy|false|false|C1704272;C2937421;C1704272;C1739363;C0020564|PROSTATICnull|Prostatic|Modifier|false|false||PROSTATICnull|Hypertrophy|Finding|false|false|C0033572|HYPERTROPHYnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Paroxysmal atrial fibrillation|Disorder|false|false|C0018792|PAROXYSMAL ATRIAL FIBRILLATIONnull|Paroxysmal|Time|false|false||PAROXYSMALnull|Atrial Fibrillation|Disorder|false|false|C0018792|ATRIAL FIBRILLATIONnull|null|Attribute|false|false|C0018792|ATRIAL FIBRILLATIONnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|ATRIAL FIBRILLATIONnull|Heart Atrium|Anatomy|false|false|C2926591;C0232197;C0235480;C0004238;C0344434|ATRIALnull|Fibrillation|Disorder|false|false|C0018792|FIBRILLATIONnull|History of surgery|Finding|false|false||Past Surgical Historynull|history of prior surgery|Finding|false|false||Surgical Historynull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Electric Countershock|Procedure|false|false||CARDIOVERSIONnull|Structure of right lower lobe of lung|Anatomy|false|false|C3539671;C1428707;C2003888;C0023928;C1552823|RIGHT LOWER LOBEnull|Table Cell Horizontal Align - right|Finding|false|false|C1548802;C1261075;C0225758|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Structure of lower lobe of lung|Anatomy|false|false|C0023928;C3539671;C1428707;C1552823;C2003888|LOWER LOBEnull|Body Site Modifier - Lower|Anatomy|false|false|C0023928;C2003888;C3539671;C1428707;C1552823|LOWERnull|Lower (action)|Event|false|false|C1548802;C1261075;C0225758|LOWERnull|Lower - spatial qualifier|Modifier|false|false||LOWERnull|AKT1S1 wt Allele|Finding|false|false|C1261075;C0796494;C0225758;C1548802|LOBE
null|AKT1S1 gene|Finding|false|false|C1261075;C0796494;C0225758;C1548802|LOBEnull|lobe|Anatomy|false|false|C0023928;C3539671;C1428707|LOBEnull|Lobectomy|Procedure|false|false|C1548802;C0796494;C0225758;C1261075|LOBECTOMYnull|Coronary Artery Bypass Surgery|Procedure|false|false|C0018787|CORONARY BYPASS SURGERYnull|Coronary Artery Bypass Surgery|Procedure|false|false|C0018787|CORONARY BYPASSnull|Heart|Anatomy|false|false|C0543467;C0038895;C1457907;C1547138;C1536078;C0010055;C0010055;C0813207|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Bypass surgery|Procedure|false|false|C0018787|BYPASS SURGERYnull|Creation of shunt|Procedure|false|false|C0018787|BYPASSnull|Level of Care - Surgery|Finding|false|false|C0018787|SURGERY
null|Surgical procedure finding|Finding|false|false|C0018787|SURGERY
null|Surgical aspects|Finding|false|false|C0018787|SURGERYnull|Operative Surgical Procedures|Procedure|false|false|C0018787|SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|Last|Modifier|false|false||lastnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scalp laceration|Disorder|false|false|C0036270|Scalp lacerationnull|Scalp structure|Anatomy|false|false|C0240937;C0043246|Scalpnull|Laceration|Disorder|false|false|C0036270|lacerationnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0036412;C2228481;C0022346|Scleranull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Icterus|Finding|false|false|C0036410|ictericnull|Icteric (color)|Modifier|false|false||ictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Conjunctival Diseases|Disorder|false|false|C0229274;C0009758|Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false|C0229274;C0009758|Conjunctiva
null|null|Finding|false|false|C0229274;C0009758|Conjunctivanull|examination of conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false|C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759|Conjunctiva
null|conjunctiva|Anatomy|false|false|C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759|Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false|C0226896|pallornull|Cyanosis|Finding|true|false|C0226896|cyanosisnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C0241137;C0010520;C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false|C0026724|mucosanull|Mucous Membrane|Anatomy|false|false|C1561514|mucosanull|Eyelid Xanthoma|Disorder|true|false||xanthelasma
null|Xanthoma|Disorder|true|false||xanthelasmanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Hepatojugular Reflex|Finding|false|false||hepatojugular reflexnull|Hepatojugular|Modifier|false|false||hepatojugularnull|Reflex motion descriptor|Finding|false|false||reflex
null|Reflex action|Finding|false|false||reflex
null|Observation of reflex|Finding|false|false||reflexnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|false|false|C3890171|murmurnull|APEX1 protein, human|Drug|false|false|C3890171|apex
null|APEX1 protein, human|Drug|false|false|C3890171|apexnull|APEX1 gene|Finding|false|false|C3890171|apexnull|dinoflagellate apex|Anatomy|false|false|C0140145;C1332102;C0018808|apexnull|Highest|Modifier|false|false||apexnull|Pericardial friction rub|Finding|true|false||rubsnull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|false|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Deformity of chest wall|Disorder|true|false|C1527391;C0817096;C0205076;C4266615|chest wall deformitiesnull|Chest wall structure|Anatomy|false|false|C0000768;C0684239;C0234233;C3164427|chest wall
null|Chest>Chest wall|Anatomy|false|false|C0000768;C0684239;C0234233;C3164427|chest wallnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0684239;C0234233;C0000768;C3164427;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0684239;C0234233;C0000768;C3164427;C0741025|chestnull|Walls of a building|Device|false|false||wallnull|Congenital Abnormality|Disorder|true|false|C0205076;C4266615;C1527391;C0817096|deformitiesnull|deformities qualifier|Modifier|false|false||deformitiesnull|Emotional tenderness|Finding|true|false|C0205076;C4266615;C1527391;C0817096|tenderness
null|Sore to touch|Finding|true|false|C0205076;C4266615;C1527391;C0817096|tendernessnull|Cell Respiration|Finding|false|false||Respiration
null|Respiration|Finding|false|false||Respirationnull|respiratory system process|Phenomenon|false|false||Respirationnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false|C4083049;C0026845|accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false|C4083049;C0026845|accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false|C0158784;C1821466;C1947944;C0042153;C0457083|muscle
null|Muscle Tissue|Anatomy|false|false|C0158784;C1821466;C1947944;C0042153;C0457083|musclenull|Use - dosing instruction imperative|Finding|false|false|C4083049;C0026845|use
null|utilization qualifier|Finding|false|false|C4083049;C0026845|use
null|Usage|Finding|false|false|C4083049;C0026845|usenull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Palpation|Procedure|false|false||palpationnull|Organomegaly|Finding|true|false||organomegalynull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|null|Phenomenon|false|false||Coolnull|Specimen Condition - Cool|Modifier|false|false||Coolnull|1+ pitting edema|Finding|false|false|C0030647|1+ pitting edemanull|Pitting edema|Finding|false|false|C0030647;C1963703;C0022742;C4299094;C0022745|pitting edemanull|Pitting|Finding|false|false|C0030647|pittingnull|Edema|Finding|false|false|C1963703;C0022742;C4299094;C0022745;C0030647|edemanull|null|Attribute|false|false||edemanull|Patella|Anatomy|false|false|C1413120;C1413079;C1720243;C0333243;C2316212;C3662487;C0006935;C0205323;C0013604;C0562271|knee capsnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745;C0030647|kneenull|Knee region structure|Anatomy|false|false|C0562271;C0013604;C0333243;C2316212;C3662487;C1413120;C1413079|knee
null|Knee|Anatomy|false|false|C0562271;C0013604;C0333243;C2316212;C3662487;C1413120;C1413079|knee
null|Lower extremity>Knee|Anatomy|false|false|C0562271;C0013604;C0333243;C2316212;C3662487;C1413120;C1413079|knee
null|Knee joint|Anatomy|false|false|C0562271;C0013604;C0333243;C2316212;C3662487;C1413120;C1413079|kneenull|capsule (pharmacologic)|Drug|false|false|C0030647|capsnull|Cryopyrin-Associated Periodic Syndromes|Disorder|false|false|C0030647;C1963703;C0022742;C4299094;C0022745|caps
null|Catastrophic antiphospholipid syndrome|Disorder|false|false|C0030647;C1963703;C0022742;C4299094;C0022745|capsnull|CAPS gene|Finding|false|false|C0030647;C1963703;C0022742;C4299094;C0022745|caps
null|CADPS gene|Finding|false|false|C0030647;C1963703;C0022742;C4299094;C0022745|capsnull|Patient Caps|Device|false|false||capsnull|Bilateral|Modifier|false|false||bilateralnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Dermatitis|Disorder|false|false||dermatitisnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKIN
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKINnull|Structure of left hand|Anatomy|false|false|C0184922;C0220797;C1546569;C3668914;C1548825;C0005558;C0741992;C1552822|left handnull|Table Cell Horizontal Align - left|Finding|false|false|C0230371|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hand problem|Finding|false|false|C4285005;C0018563;C0230371|handnull|Upper extremity>Hand|Anatomy|false|false|C0741992|hand
null|Hand|Anatomy|false|false|C0741992|handnull|Numerous|LabModifier|false|false||Multiplenull|null|Procedure|false|false|C0230371|open biopsynull|Open|Modifier|false|false||opennull|biopsy characteristics|Finding|false|false|C0230371|biopsy
null|null|Finding|false|false|C0230371|biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false|C0230371|biopsy
null|Biopsy|Procedure|false|false|C0230371|biopsy
null|Consent Type - biopsy|Procedure|false|false|C0230371|biopsynull|Excision|Procedure|false|false||excision
null|removal technique|Procedure|false|false||excisionnull|Site|Modifier|false|false||sitesnull|Anterior part of left leg|Anatomy|false|false||left shinnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Shin|Anatomy|false|false||shinnull|Posterior part of right leg|Anatomy|false|false|C1552823|right calfnull|Table Cell Horizontal Align - right|Finding|false|false|C0489801|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Palpable|Modifier|false|false||palpablenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|physical examination (physical finding)|Finding|false|false||Physical examnull|Physical Examination|Procedure|false|false||Physical examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|Last|Modifier|false|false||lastnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Elderly (population group)|Subject|false|false||elderlynull|Old age|Time|false|false||elderlynull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false|C0036270|dressing
null|Ability to dress|Finding|false|false|C0036270|dressingnull|Dressing patient (procedure)|Procedure|false|false|C0036270|dressing
null|Dressing of skin or wound|Procedure|false|false|C0036270|dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Scalp structure|Anatomy|false|false|C0152053;C0278286;C0085639;C1305428;C0518459|scalpnull|Recent|Time|false|false||recentnull|Falls|Finding|false|false|C0036270;C0036270|fallnull|Autumn|Time|false|false||fallnull|Scalp structure|Anatomy|false|false|C0085639|scalpnull|Laceration|Disorder|false|false||lacerationnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0036412;C2228481;C0022346|Scleranull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Icterus|Finding|false|false|C0036410|ictericnull|Icteric (color)|Modifier|false|false||ictericnull|Pupil|Anatomy|false|false||pupilsnull|Round shape|Modifier|false|false||roundnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Jugular venous pressure|Finding|false|false||JVPnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Hepatojugular Reflex|Finding|false|false||hepatojugular reflexnull|Hepatojugular|Modifier|false|false||hepatojugularnull|Reflex motion descriptor|Finding|false|false||reflex
null|Reflex action|Finding|false|false||reflex
null|Observation of reflex|Finding|false|false||reflexnull|Irregular|Modifier|false|false||irregularnull|Structure of precordium|Anatomy|false|false||precordiumnull|Quiet|Modifier|false|false||quietnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||heavenull|Second heart sound split|Finding|false|false||split S2null|Splitting|Finding|false|false||splitnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Heart murmur|Finding|false|false|C3890171|murmurnull|APEX1 protein, human|Drug|false|false|C3890171|apex
null|APEX1 protein, human|Drug|false|false|C3890171|apexnull|APEX1 gene|Finding|false|false|C3890171|apexnull|dinoflagellate apex|Anatomy|false|false|C0018808;C0140145;C1332102|apexnull|Highest|Modifier|false|false||apexnull|Lung|Anatomy|false|false||LUNGSnull|Exertion|Finding|false|false||effortnull|Legal fine|Entity|false|false||Finenull|Fine (qualifier value)|Modifier|false|false||Finenull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|1+ pitting edema|Finding|false|false|C1140621;C0023216|1+ pitting edemanull|Pitting edema|Finding|false|false|C1140621;C0023216|pitting edemanull|Pitting|Finding|false|false|C1140621;C0023216;C1140621;C0023216|pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Leg|Anatomy|false|false|C0205323|leg
null|Lower Extremity|Anatomy|false|false|C0205323|legnull|Leg|Anatomy|false|false|C1720243;C0205323;C0333243|leg
null|Lower Extremity|Anatomy|false|false|C1720243;C0205323;C0333243|legnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Numerous|LabModifier|false|false||Multiplenull|Excision biopsy|Procedure|false|false||excision biopsynull|Excision|Procedure|false|false|C1140621|excision
null|removal technique|Procedure|false|false|C1140621|excisionnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false|C1140621|biopsy
null|Biopsy|Procedure|false|false|C1140621|biopsy
null|Consent Type - biopsy|Procedure|false|false|C1140621|biopsynull|Traumatic Wound|Disorder|false|false|C1140621|woundsnull|Wounds - qualifier|Modifier|false|false||woundsnull|Leg|Anatomy|false|false|C0015252;C0728940;C5781420;C0043250;C3668914;C1548825;C0005558|legsnull|null|Attribute|false|false|C1140621|legsnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Ferritin|Drug|false|false||FERRITIN
null|Ferritin|Drug|false|false||FERRITIN
null|Ferritin|Drug|false|false||FERRITINnull|Ferritin measurement|Procedure|false|false||FERRITINnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|Iron Drug Class|Drug|false|false||IRON
null|iron|Drug|false|false||IRON
null|iron|Drug|false|false||IRON
null|iron|Drug|false|false||IRON
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||IRONnull|Iron measurement|Procedure|false|false||IRONnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C0201899;C0004002;C0242192;C1121182;C4522245;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hyalin Substance|Finding|false|false||HYALINEnull|Hyaline (appearance)|Modifier|false|false||HYALINEnull|null|Lab|false|false|C0014792|URINE  RBC
null|Red blood cells urine positive|Lab|false|false|C0014792|URINE  RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0221752;C2188659;C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Leukocytes|Anatomy|false|false|C1510439|WBCnull|bacteria aspects|Finding|false|false|C0023516|BACTERIAnull|Bacteria <walking sticks>|Entity|false|false||BACTERIA
null|Bacteria|Entity|false|false||BACTERIAnull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPInull|Exocrine pancreatic insufficiency|Disorder|false|false||EPInull|Eysenck personality inventory|Finding|false|false||EPI
null|TFPI wt Allele|Finding|false|false||EPI
null|TFPI gene|Finding|false|false||EPInull|Electronic Portal Imaging|Procedure|false|false||EPI
null|Echo-Planar Imaging|Procedure|false|false||EPInull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C0004002;C0242192;C1121182;C1415181;C1420113;C5960784;C4522245|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|infant weight for previous delivery (history)|Finding|false|false||WEIGHT
null|Weight symptom (finding)|Finding|false|false||WEIGHTnull|Weighing patient|Procedure|false|false||WEIGHTnull|null|Attribute|false|false||WEIGHTnull|Body Weight|Subject|false|false||WEIGHTnull|Importance Weight|Modifier|false|false||WEIGHTnull|Weight|LabModifier|false|false||WEIGHTnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Diuretic [APC]|Drug|false|false||DIURETIC
null|Diuretics|Drug|false|false||DIURETICnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONnull|medication - HL7 publishing domain|Finding|false|false||MEDICATION
null|Medications|Finding|false|false||MEDICATIONnull|Changing|Finding|false|false||CHANGESnull|Changed status|LabModifier|false|false||CHANGESnull|Daily|Time|false|false||dailynull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|mEq|LabModifier|false|false||mEqnull|Daily|Time|false|false||dailynull|mEq|LabModifier|false|false||mEqnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|4 Weeks|Time|false|false||4 weeksnull|week|Time|false|false||weeksnull|Electrolyte [EPC]|Drug|false|false||electrolyte
null|Electrolytes|Drug|false|false||electrolyte
null|Electrolytes|Drug|false|false||electrolytenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|CODE STATUS|Procedure|false|false||CODE STATUSnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|What subject filter - Status|Finding|false|false||STATUSnull|null|Attribute|false|false||STATUSnull|Social status|Modifier|false|false||STATUS
null|Status|Modifier|false|false||STATUSnull|Full|Modifier|false|false||fullnull|Health Care|Procedure|false|false||Health carenull|Health|Finding|false|false||Healthnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Advance Directive - Proxy|Finding|false|false||proxynull|Proxy|Subject|false|false||proxynull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Health Care|Procedure|false|false||health carenull|Health|Finding|false|false||healthnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Advance Directive - Proxy|Finding|false|false||proxynull|Proxy|Subject|false|false||proxynull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Telephone Number|Finding|false|false||Phone numbernull|Authorization Mode - Phone|Finding|false|false||Phone
null|Visit User Code - Phone|Finding|false|false||Phone
null|Telephone Number|Finding|false|false||Phone
null|MDFAttributeType - Phone|Finding|false|false||Phonenull|Telephone|Device|false|false||Phonenull|Person location type - Phone|Modifier|false|false||Phonenull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|Patient summary|Finding|false|false||PATIENT SUMMARYnull|Relationship modifier - Patient|Finding|false|false||PATIENT
null|Specimen Type - Patient|Finding|false|false||PATIENT
null|Mail Claim Party - Patient|Finding|false|false||PATIENT
null|Report source - Patient|Finding|false|false||PATIENT
null|null|Finding|false|false||PATIENT
null|Disabled Person Code - Patient|Finding|false|false||PATIENTnull|Patients|Subject|false|false||PATIENTnull|Veterinary Patient|Entity|false|false||PATIENTnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Tricuspid|Modifier|false|false||tricuspidnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Right Ventricular Dysfunction|Finding|false|false|C0018827|right ventricular dysfunctionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Ventricular Dysfunction|Finding|false|false|C0018827|ventricular dysfunctionnull|Heart Ventricle|Anatomy|false|false|C0242973;C0242707;C3887505;C0031847;C0277785;C3887504|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false|C0018827|dysfunction
null|physiopathological|Finding|false|false|C0018827|dysfunction
null|Functional disorder|Finding|false|false|C0018827|dysfunctionnull|Moderate - Severity of Illness Code|Finding|false|false|C0024109|moderate
null|Moderate|Finding|false|false|C0024109|moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C5201148;C1547226;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Hypertensive disease|Disorder|false|false||hypertensionnull|Paroxysmal atrial fibrillation|Disorder|false|false|C0018792|paroxysmal atrial fibrillationnull|Paroxysmal|Time|false|false||paroxysmalnull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0232197;C0004238;C0235480;C2926591;C0344434|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C4554465;C0869841;C1552824;C0022658;C0812426;C1561643;C0496927;C0496892|kidney
null|Both kidneys|Anatomy|false|false|C4554465;C0869841;C1552824;C0022658;C0812426;C1561643;C0496927;C0496892|kidneynull|Disease|Disorder|false|false||diseasenull|BaseLine dental cement|Drug|false|false||Baselinenull|baseline - TableCellVerticalAlign|Finding|false|false|C0227665;C0022646|Baselinenull|Baseline|LabModifier|false|false||Baselinenull|Cerebrovascular Disorders|Disorder|false|false||cerebrovascular diseasenull|Cerebrovascular|Modifier|false|false||cerebrovascularnull|Disease|Disorder|false|false||diseasenull|Metastatic melanoma|Disorder|false|false||metastatic melanomanull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Cell Cycle Checkpoints|Finding|false|false||checkpointnull|Inhibitor|Drug|false|false||inhibitornull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Dyspnea on exertion|Finding|false|false||DOEnull|Department of Energy|Subject|false|false||DOEnull|Adult female goat|Entity|false|false||DOEnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Diuresis|Finding|false|false||diuresisnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Main|Modifier|false|false||Main
null|Primary|Modifier|false|false||Mainnull|Double coronary vessel disease|Disorder|false|false|C0010075;C0018787|two vessel coronary diseasenull|Coronary Vessels|Anatomy|false|false|C0581375|vessel coronarynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Disease|Disorder|false|false|C0018787|coronary disease
null|Coronary heart disease|Disorder|false|false|C0018787|coronary diseasenull|Heart|Anatomy|false|false|C0012634;C0581375;C1956346;C0010068|coronarynull|Coronary|Modifier|false|false||coronarynull|Disease|Disorder|false|false|C0018787|diseasenull|matrix metalloproteinase 7 activity|Finding|false|false||PUMPnull|null|Device|false|false||PUMPnull|Pump Dosing Unit|LabModifier|false|false||PUMPnull|Rhythm|Finding|false|false||RHYTHM
null|rhythmic process (biological)|Finding|false|false||RHYTHMnull|Ectopic rhythm|Disorder|false|false|C4050503|Ectopic rhythmnull|Ectopic Graft|Anatomy|false|false|C1399226|Ectopicnull|Ectopic|Modifier|false|false||Ectopicnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Prolonged PR interval|Finding|false|false||PR prolongationnull|Left axis deviation|Finding|false|false|C0004457|left axis deviationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|axis deviation|Finding|false|false|C0004457|axis deviationnull|Fracture of second cervical vertebra|Disorder|false|false|C0004457|axisnull|Axis vertebra|Anatomy|false|false|C0232297;C0262387;C0349013|axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|Protocol Deviation|Finding|false|false||deviationnull|Spatial Displacement|Modifier|false|false||deviation
null|Variant|Modifier|false|false||deviationnull|Right bundle branch block|Disorder|false|false||RBBBnull|null|Finding|false|false||RBBBnull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|Reduced left ventricular ejection fraction|Finding|false|false||reduced ejection fractionnull|stress echo measurements ejection fraction|Finding|false|false||ejection fraction
null|Ejection fraction|Finding|false|false||ejection fractionnull|Ejection fraction (procedure)|Procedure|false|false||ejection fractionnull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|MDFAttributeType - Fraction|Finding|false|false||fractionnull|Fraction of|LabModifier|false|false||fractionnull|Right Ventricular Dysfunction|Finding|false|false|C0018827|Right ventricular dysfunctionnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Ventricular Dysfunction|Finding|false|false|C0018827|ventricular dysfunctionnull|Heart Ventricle|Anatomy|false|false|C3887505;C0242973;C0031847;C0277785;C3887504;C0242707|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false|C0018827|dysfunction
null|physiopathological|Finding|false|false|C0018827|dysfunction
null|Functional disorder|Finding|false|false|C0018827|dysfunctionnull|Pulmonary ventilator management|Procedure|false|false||pulmnull|Hypertensive disease|Disorder|false|false||HTNnull|Hypervolemia (finding)|Finding|false|false||Volume overloadnull|Volume (publication)|Finding|false|false||Volumenull|Volume|LabModifier|false|false||Volumenull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exacerbation|Finding|false|false||exacerbationnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Recent|Time|false|false||recentnull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|In addition to|Finding|false|false||in addition tonull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Titration Method|Procedure|false|false||titrationnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Past Week|Time|false|false||last weeknull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Document Confidentiality Status - Restricted|Finding|false|false||restricted
null|Confidentiality - restricted|Finding|false|false||restricted
null|Confidentiality code - Restricted|Finding|false|false||restricted
null|Restricted|Finding|false|false||restrictednull|Fluid intake|LabModifier|false|false||fluid intakenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Eyeglasses|Device|false|false||glassesnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Juice|Drug|false|false||juicenull|Daily|Time|false|false||dailynull|Guideline (Publication Type)|Finding|false|false||guideline
null|Guidelines|Finding|false|false||guidelinenull|disposition medical therapy|Procedure|false|false||medical therapy
null|Medical therapy|Procedure|false|false||medical therapynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Acute kidney injury|Disorder|false|false|C0227665;C0022646|acute kidney injury
null|Kidney Failure, Acute|Disorder|false|false|C0227665;C0022646|acute kidney injurynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Injury of kidney|Disorder|false|false|C0227665;C0022646|kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidney
null|examination of kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C3263723;C3263722;C0022660;C2609414;C0160420;C0496927;C0496892;C4554465;C0869841;C0812426|kidney
null|Both kidneys|Anatomy|false|false|C3263723;C3263722;C0022660;C2609414;C0160420;C0496927;C0496892;C4554465;C0869841;C0812426|kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false|C0227665;C0022646|injury
null|Traumatic injury|Disorder|false|false|C0227665;C0022646|injurynull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Hypertransaminasaemia|Finding|false|false||transaminitisnull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Response Modality - Bolus|Finding|false|false||bolus
null|Bolus of ingested food|Finding|false|false||bolusnull|bolus infusion|Procedure|false|false||bolusnull|Bolus Dosing Unit|LabModifier|false|false||bolusnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Good response|Finding|false|false||good responsenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Transition Mutation|Disorder|false|false||transitionnull|Transition (action)|Event|false|false||transitionnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||dailynull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Reduced|Finding|true|false||reductionnull|Reduction procedure|Procedure|true|false||reduction
null|Surgical reduction|Procedure|true|false||reductionnull|Reduction (chemical)|Phenomenon|true|false||reductionnull|Neural|Finding|false|false||neuralnull|Hormonal|Modifier|false|false||hormonalnull|Blockade|Drug|false|false||blockade
null|Blockade|Drug|false|false||blockadenull|Blocking|Finding|false|false||blockadenull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|Chronic Kidney Diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|Kidney Diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|Kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|Kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|Kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|Kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|Kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C1561643;C0012634;C0022658;C4554465;C0869841;C0812426|Kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C1561643;C0012634;C0022658;C4554465;C0869841;C0812426|Kidneynull|Disease|Disorder|false|false|C0227665;C0022646|Diseasenull|BaseLine dental cement|Drug|false|false||Baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||Baselinenull|Baseline|LabModifier|false|false||Baselinenull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Initially|Time|false|false||initiallynull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|DIURETIC USAGE|Finding|false|false||diuretic usagenull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|Usage|Finding|false|false||usagenull|Diuretics|Drug|false|false||diureticsnull|Smaller|Modifier|false|false||Lessnull|Less Than|LabModifier|false|false||Lessnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Cardio-Renal Syndrome|Disorder|false|false||cardiorenal syndromenull|Syndrome|Disorder|false|false||syndromenull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recent|Time|false|false||recentlynull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|nephrology (field)|Title|false|false||nephrologynull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumab
null|pembrolizumab|Drug|false|false||pembrolizumabnull|More|LabModifier|false|false||morenull|Adverse Event Probably Related to Intervention|Modifier|false|false||likely relatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false|C0022646|related
null|Related (finding)|Finding|false|false|C0022646|relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0445223;C1552599;C0042075|renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Metastatic melanoma|Disorder|false|false||Metastatic Melanomanull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Melanoma vaccine|Drug|false|false||Melanoma
null|Melanoma vaccine|Drug|false|false||Melanomanull|melanoma|Disorder|false|false||Melanomanull|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumab
null|pembrolizumab|Drug|false|false||Pembrolizumabnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Renal function|Finding|false|false|C0227665;C0022646|kidney functionnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0232804;C0496927;C0496892;C4554465;C0869841;C0812426;C0598463;C0542341;C1705273;C0031843|kidney
null|Both kidneys|Anatomy|false|false|C0232804;C0496927;C0496892;C4554465;C0869841;C0812426;C0598463;C0542341;C1705273;C0031843|kidneynull|Function (attribute)|Finding|false|false|C0227665;C0022646|function
null|physiological aspects|Finding|false|false|C0227665;C0022646|function
null|Mathematical Operator|Finding|false|false|C0227665;C0022646|function
null|Functional Status|Finding|false|false|C0227665;C0022646|functionnull|Function Axis|Subject|false|false||functionnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK MBnull|Creatine kinase MB measurement|Procedure|false|false||CK MBnull|Concern|Finding|false|false||concernnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Myocarditis|Disorder|false|false||myocarditisnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|follow-up|Procedure|false|false||Followupnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statinnull|EEF1A2 gene|Finding|false|false||Statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||Statinnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|During admission|Time|false|false||during admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Increased frequency of micturition|Finding|false|false|C0042027|Urinary frequencynull|Urinary tract|Anatomy|false|false|C4321352;C3898838;C0042023|Urinarynull|urinary|Modifier|false|false||Urinarynull|Frequency|Finding|false|false|C0042027|frequency
null|How Often|Finding|false|false|C0042027|frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Apyrexial|Finding|false|false||Afebrilenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|tamsulosin|Drug|false|false||tamsulosin
null|tamsulosin|Drug|false|false||tamsulosinnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0018787;C0205042|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0018787;C0205042|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C5550999;C0398738;C1956346;C0010054;C0012634;C1414063;C1706333;C0852949|Coronary arterynull|Heart|Anatomy|false|false|C1956346;C0010054|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042|artery diseasenull|Arterial system|Anatomy|false|false|C1956346;C0010054;C0852949;C0012634|artery
null|Arteries|Anatomy|false|false|C1956346;C0010054;C0852949;C0012634|arterynull|Disease|Disorder|false|false|C0226004;C0003842;C0205042|diseasenull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0205042;C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0205042;C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0205042;C0226032|LAD
null|DLD gene|Finding|false|false|C0205042;C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1532338;C1514496;C4724254;C4049621;C1418370;C1705930;C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false|C0226032|PCI
null|SERPINA5 wt Allele|Finding|false|false|C0226032|PCI
null|SERPINA5 gene|Finding|false|false|C0226032|PCInull|Percutaneous Coronary Intervention|Procedure|false|false|C0226032|PCI
null|photochemical internalization|Procedure|false|false|C0226032|PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false|C0226032|PCInull|Picocurie|LabModifier|false|false||PCInull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Daily|Time|false|false||dailynull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statinnull|EEF1A2 gene|Finding|false|false||Statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||Statinnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Paroxysmal atrial fibrillation|Disorder|false|false|C0018792|Paroxysmal Atrial fibrillationnull|Paroxysmal|Time|false|false||Paroxysmalnull|Atrial Fibrillation|Disorder|false|false|C0018792|Atrial fibrillationnull|null|Attribute|false|false|C0018792|Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|Atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0235480;C0004238;C0344434;C0232197;C2926591|Atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Strategy|Finding|false|false||strategynull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Safety|Phenomenon|false|false||safetynull|Laboratory test finding|Lab|false|false||labsnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Further|Modifier|false|false||furthernull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Align|Drug|false|false||Align
null|Align|Drug|false|false||Alignnull|herbal medicines bifidobacterium infantis|Drug|false|false||bifidobacterium infantisnull|Bifidobacterium longum subspecies infantis|Entity|false|false||bifidobacterium infantis
null|Bifidobacterium infantis|Entity|false|false||bifidobacterium infantisnull|Bifidobacterium|Entity|false|false||bifidobacteriumnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10null|Coenzymes|Drug|false|false||coenzyme
null|Coenzymes|Drug|false|false||coenzymenull|AGO2 wt Allele|Finding|false|false||Q10
null|AGO2 gene|Finding|false|false||Q10null|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|tamsulosin|Drug|false|false||Tamsulosin
null|tamsulosin|Drug|false|false||Tamsulosinnull|Once a day, at bedtime|Time|false|false||QHSnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|cephalexin|Drug|false|false||Cephalexin
null|cephalexin|Drug|false|false||Cephalexinnull|Every six hours|Time|false|false||Q6Hnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|Daily|Time|false|false||DAILYnull|potassium chloride|Drug|false|false||potassium chloride
null|potassium chloride|Drug|false|false||potassium chloridenull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|chloride ion|Drug|false|false||chloride
null|Chlorides|Drug|false|false||chloridenull|Chloride metabolic function|Finding|false|false||chloridenull|Chloride measurement|Procedure|false|false||chloridenull|mEq|LabModifier|false|false||mEqnull|Packet - container|Device|false|false||packet
null|Packet (device)|Device|false|false||packetnull|Packet Dosing Unit|LabModifier|false|false||packetnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1720092;C1527415|mouth
null|Oral region|Anatomy|false|false|C1720092;C1527415|mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false|C0230028;C0226896|oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Align|Drug|false|false||Align
null|Align|Drug|false|false||Alignnull|herbal medicines bifidobacterium infantis|Drug|false|false||bifidobacterium infantisnull|Bifidobacterium longum subspecies infantis|Entity|false|false||bifidobacterium infantis
null|Bifidobacterium infantis|Entity|false|false||bifidobacterium infantisnull|Bifidobacterium|Entity|false|false||bifidobacteriumnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10null|Coenzymes|Drug|false|false||coenzyme
null|Coenzymes|Drug|false|false||coenzymenull|AGO2 wt Allele|Finding|false|false||Q10
null|AGO2 gene|Finding|false|false||Q10null|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|tamsulosin|Drug|false|false||Tamsulosin
null|tamsulosin|Drug|false|false||Tamsulosinnull|Once a day, at bedtime|Time|false|false||QHSnull|tamsulosin|Drug|false|false||tamsulosin
null|tamsulosin|Drug|false|false||tamsulosinnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0807726;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0807726;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false|C0524463;C1325531|Refillsnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary Diagnosisnull|Principal diagnosis|Modifier|false|false||Primary Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Secondary diagnosis|Finding|false|false||Secondary diagnosisnull|null|Attribute|false|false||Secondary diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Hypertransaminasaemia|Finding|false|false||Transaminitisnull|Metastatic melanoma|Disorder|false|false||Metastatic melanomanull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Melanoma vaccine|Drug|false|false||melanoma
null|Melanoma vaccine|Drug|false|false||melanomanull|melanoma|Disorder|false|false||melanomanull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0018787;C0205042|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0018787;C0205042|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C0012634;C0010055;C1414063;C1706333;C0852949;C1956346;C0010054;C5550999;C0398738|Coronary arterynull|Heart|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|artery diseasenull|Arterial system|Anatomy|false|false|C1956346;C0010054;C0010055;C0852949;C5550999;C0398738;C1414063;C1706333;C0012634|artery
null|Arteries|Anatomy|false|false|C1956346;C0010054;C0010055;C0852949;C5550999;C0398738;C1414063;C1706333;C0012634|arterynull|Disease|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|diseasenull|Coronary Artery Bypass Surgery|Procedure|false|false|C0205042;C0226004;C0003842|CABGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032;C0226004;C0003842;C0205042|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032;C0226004;C0003842;C0205042|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032;C0205042;C0226004;C0003842|LAD
null|DLD gene|Finding|false|false|C0226032;C0205042;C0226004;C0003842|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Discharge instructions|Finding|false|false||DISCHARGE INSTRUCTIONSnull|hospital discharge instructions (treatment)|Procedure|false|false||DISCHARGE INSTRUCTIONSnull|null|Attribute|false|false||DISCHARGE INSTRUCTIONSnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Instructions|Finding|false|false||INSTRUCTIONS
null|Instruction [Publication Type]|Finding|false|false||INSTRUCTIONSnull|null|Attribute|false|false||INSTRUCTIONSnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Dyspnea|Finding|false|false||short of breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Lung|Anatomy|false|false||lungsnull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Hardness|Modifier|false|false||hardnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false|C0004600|fluidnull|Fluid behavior|Modifier|false|false||fluidnull|null|Anatomy|false|false|C1546638|backsnull|Lung|Anatomy|false|false||lungsnull|Occur (action)|Event|false|false||HAPPENEDnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Patient need for (contextual qualifier)|Finding|false|false||NEEDnull|Needs|Modifier|false|false||NEEDnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Follow-up status|Finding|false|false||Follow upnull|follow-up|Procedure|false|false||Follow upnull|Follow - dosing instruction imperative|Finding|false|false||Follow
null|Follow|Finding|false|false||Follownull|Followed by|Time|false|false||Follownull|Physicians|Subject|false|false||doctorsnull|Every morning|Time|false|false||every morningnull|Morning|Time|false|false||morningnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Pounds|LabModifier|false|false||poundsnull|Call - dosing instruction fragment|Finding|false|false||Call
null|Call (Instruction)|Finding|false|false||Call
null|Decision|Finding|false|false||Call
null|CHL1 gene|Finding|false|false||Callnull|ITPRIP gene|Finding|false|false||dangernull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions