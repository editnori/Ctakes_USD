 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Shortness|293,302
of|303,305
breath|306,312
<EOL>|312,313
<EOL>|314,315
Major|315,320
Surgical|321,329
or|330,332
Invasive|333,341
Procedure|342,351
:|351,352
<EOL>|352,353
None|353,357
<EOL>|357,358
<EOL>|359,360
Ms.|388,391
_|392,393
_|393,394
_|394,395
is|396,398
a|399,400
_|401,402
_|402,403
_|403,404
with|405,409
hx|410,412
COPD|413,417
on|418,420
home|421,425
O2|426,428
,|428,429
atrial|430,436
<EOL>|437,438
fibrillation|438,450
on|451,453
apixaban|454,462
,|462,463
hypertension|464,476
,|476,477
CAD|478,481
,|481,482
and|483,486
hyperlipidemia|487,501
<EOL>|502,503
who|503,506
presented|507,516
with|517,521
dyspnea|522,529
.|529,530
<EOL>|532,533
She|533,536
has|537,540
had|541,544
multiple|545,553
prior|554,559
admissions|560,570
for|571,574
dyspnea|575,582
.|582,583
She|584,587
was|588,591
<EOL>|592,593
recently|593,601
discharged|602,612
on|613,615
_|616,617
_|617,618
_|618,619
after|620,625
3|626,627
day|628,631
inpatient|632,641
admission|642,651
for|652,655
<EOL>|656,657
COPD|657,661
exacerbation|662,674
.|674,675
She|676,679
was|680,683
discharged|684,694
on|695,697
extended|698,706
prednisone|707,717
<EOL>|718,719
taper|719,724
with|725,729
plan|730,734
for|735,738
5d|739,741
40mg|742,746
Prednisone|747,757
(|758,759
to|759,761
finish|762,768
_|769,770
_|770,771
_|771,772
followed|773,781
<EOL>|782,783
by|783,785
10mg|786,790
taper|791,796
every|797,802
5|803,804
days|805,809
(|810,811
35mg|811,815
from|816,820
_|821,822
_|822,823
_|823,824
,|824,825
30mg|826,830
_|831,832
_|832,833
_|833,834
,|834,835
<EOL>|836,837
etc|837,840
...|840,843
)|843,844
.|844,845
She|846,849
initially|850,859
went|860,864
to|865,867
rehab|868,873
and|874,877
subsequently|878,890
went|891,895
home|896,900
<EOL>|901,902
2|902,903
days|904,908
prior|909,914
to|915,917
admission|918,927
.|927,928
<EOL>|930,931
Upon|931,935
arrival|936,943
at|944,946
home|947,951
she|952,955
subsequently|956,968
had|969,972
recrudescence|973,986
of|987,989
<EOL>|990,991
fatigue|991,998
,|998,999
wheezing|1000,1008
,|1008,1009
dyspnea|1010,1017
.|1017,1018
She|1019,1022
also|1023,1027
had|1028,1031
increased|1032,1041
O2|1042,1044
<EOL>|1045,1046
requirements|1046,1058
(|1059,1060
up|1060,1062
to|1063,1065
3L|1066,1068
,|1068,1069
using|1070,1075
oxygen|1076,1082
24hr|1083,1087
instead|1088,1095
of|1096,1098
during|1099,1105
day|1106,1109
<EOL>|1110,1111
only|1111,1115
)|1115,1116
.|1116,1117
Also|1118,1122
with|1123,1127
new|1128,1131
cough|1132,1137
,|1137,1138
non-productive|1139,1153
.|1153,1154
Denies|1155,1161
f|1162,1163
/|1163,1164
c|1164,1165
,|1165,1166
CP|1167,1169
.|1169,1170
No|1171,1173
<EOL>|1174,1175
n|1175,1176
/|1176,1177
v|1177,1178
,|1178,1179
no|1180,1182
myalgias|1183,1191
.|1191,1192
Decreased|1193,1202
hearing|1203,1210
in|1211,1213
right|1214,1219
ear|1220,1223
with|1224,1228
fullness|1229,1237
<EOL>|1238,1239
for|1239,1242
past|1243,1247
4|1248,1249
days|1250,1254
.|1254,1255
She|1256,1259
was|1260,1263
seen|1264,1268
by|1269,1271
PCP|1272,1275
_|1276,1277
_|1277,1278
_|1278,1279
noted|1280,1285
to|1286,1288
have|1289,1293
<EOL>|1294,1295
inspiratory|1295,1306
/|1306,1307
expiratory|1307,1317
wheezes|1318,1325
,|1325,1326
as|1327,1329
well|1330,1334
as|1335,1337
decreased|1338,1347
hearing|1348,1355
and|1356,1359
<EOL>|1360,1361
bulging|1361,1368
TM|1369,1371
right|1372,1377
ear|1378,1381
.|1381,1382
She|1383,1386
was|1387,1390
referred|1391,1399
to|1400,1402
the|1403,1406
_|1407,1408
_|1408,1409
_|1409,1410
ED|1411,1413
for|1414,1417
<EOL>|1418,1419
further|1419,1426
management|1427,1437
.|1437,1438
<EOL>|1440,1441
In|1441,1443
the|1444,1447
ED|1448,1450
,|1450,1451
initial|1452,1459
vital|1460,1465
signs|1466,1471
were|1472,1476
:|1476,1477
98.4|1478,1482
74|1483,1485
142|1486,1489
/|1489,1490
69|1490,1492
16|1493,1495
100|1496,1499
%|1499,1500
(|1500,1501
2L|1501,1503
<EOL>|1504,1505
NC|1505,1507
)|1507,1508
<EOL>|1510,1511
-|1511,1512
Labs|1513,1517
were|1518,1522
notable|1523,1530
for|1531,1534
:|1534,1535
<EOL>|1537,1538
136|1539,1542
95|1543,1545
17|1546,1548
140|1549,1552
<EOL>|1554,1555
3.5|1556,1559
29|1560,1562
1.0|1563,1566
<EOL>|1568,1569
BNP|1570,1573
254|1574,1577
<EOL>|1579,1580
CBC|1581,1584
within|1585,1591
normal|1592,1598
limits|1599,1605
,|1605,1606
but|1607,1610
with|1611,1615
neutrophil|1616,1626
predominance|1627,1639
<EOL>|1641,1642
UA|1643,1645
with|1646,1650
30|1651,1653
protein|1654,1661
<EOL>|1663,1664
VBG|1665,1668
:|1668,1669
pH|1670,1672
7.45|1673,1677
,|1677,1678
pCO2|1679,1683
43|1684,1686
,|1686,1687
pO2|1688,1691
59|1692,1694
,|1694,1695
HCO3|1696,1700
31|1701,1703
<EOL>|1705,1706
Flu|1707,1710
PCR|1711,1714
negative|1715,1723
<EOL>|1725,1726
-|1726,1727
Imaging|1728,1735
:|1735,1736
<EOL>|1738,1739
CXR|1740,1743
notable|1744,1751
for|1752,1755
no|1756,1758
acute|1759,1764
cardiopulmonary|1765,1780
process|1781,1788
.|1788,1789
<EOL>|1791,1792
-|1792,1793
The|1794,1797
patient|1798,1805
was|1806,1809
given|1810,1815
:|1815,1816
<EOL>|1818,1819
_|1820,1821
_|1821,1822
_|1822,1823
16|1824,1826
:|1826,1827
03|1827,1829
IH|1830,1832
Albuterol|1833,1842
0.083|1843,1848
%|1848,1849
Neb|1850,1853
Soln|1854,1858
1|1859,1860
NEB|1861,1864
<EOL>|1866,1867
_|1868,1869
_|1869,1870
_|1870,1871
16|1872,1874
:|1874,1875
03|1875,1877
IH|1878,1880
Ipratropium|1881,1892
Bromide|1893,1900
Neb|1901,1904
1|1905,1906
NEB|1907,1910
<EOL>|1912,1913
_|1914,1915
_|1915,1916
_|1916,1917
17|1918,1920
:|1920,1921
12|1921,1923
IH|1924,1926
Albuterol|1927,1936
0.083|1937,1942
%|1942,1943
Neb|1944,1947
Soln|1948,1952
1|1953,1954
NEB|1955,1958
<EOL>|1960,1961
_|1962,1963
_|1963,1964
_|1964,1965
17|1966,1968
:|1968,1969
12|1969,1971
IH|1972,1974
Ipratropium|1975,1986
Bromide|1987,1994
Neb|1995,1998
1|1999,2000
NEB|2001,2004
<EOL>|2006,2007
_|2008,2009
_|2009,2010
_|2010,2011
18|2012,2014
:|2014,2015
12|2015,2017
IH|2018,2020
Albuterol|2021,2030
0.083|2031,2036
%|2036,2037
Neb|2038,2041
Soln|2042,2046
1|2047,2048
NEB|2049,2052
<EOL>|2054,2055
_|2056,2057
_|2057,2058
_|2058,2059
18|2060,2062
:|2062,2063
12|2063,2065
IH|2066,2068
Ipratropium|2069,2080
Bromide|2081,2088
Neb|2089,2092
1|2093,2094
NEB|2095,2098
<EOL>|2100,2101
_|2102,2103
_|2103,2104
_|2104,2105
21|2106,2108
:|2108,2109
05|2109,2111
IH|2112,2114
Albuterol|2115,2124
0.083|2125,2130
%|2130,2131
Neb|2132,2135
Soln|2136,2140
1|2141,2142
NEB|2143,2146
<EOL>|2148,2149
_|2150,2151
_|2151,2152
_|2152,2153
21|2154,2156
:|2156,2157
05|2157,2159
PO|2160,2162
PredniSONE|2163,2173
60|2174,2176
mg|2177,2179
<EOL>|2181,2182
_|2183,2184
_|2184,2185
_|2185,2186
21|2187,2189
:|2189,2190
05|2190,2192
IV|2193,2195
Magnesium|2196,2205
Sulfate|2206,2213
2|2214,2215
gm|2216,2218
<EOL>|2220,2221
_|2222,2223
_|2223,2224
_|2224,2225
21|2226,2228
:|2228,2229
33|2229,2231
IH|2232,2234
Albuterol|2235,2244
0.083|2245,2250
%|2250,2251
Neb|2252,2255
Soln|2256,2260
1|2261,2262
NEB|2263,2266
<EOL>|2268,2269
Vitals|2270,2276
prior|2277,2282
to|2283,2285
transfer|2286,2294
were|2295,2299
:|2299,2300
<EOL>|2302,2303
98.8|2304,2308
87|2309,2311
131|2312,2315
/|2315,2316
83|2316,2318
16|2319,2321
97|2322,2324
%|2324,2325
(|2326,2327
2L|2327,2329
)|2329,2330
<EOL>|2332,2333
Upon|2333,2337
arrival|2338,2345
to|2346,2348
the|2349,2352
floor|2353,2358
,|2358,2359
she|2360,2363
complained|2364,2374
of|2375,2377
wheezing|2378,2386
and|2387,2390
SOB|2391,2394
,|2394,2395
<EOL>|2396,2397
and|2397,2400
persistent|2401,2411
decreased|2412,2421
hearing|2422,2429
with|2430,2434
fullness|2435,2443
in|2444,2446
right|2447,2452
ear|2453,2456
.|2456,2457
<EOL>|2459,2460
<EOL>|2461,2462
REVIEW|2462,2468
OF|2469,2471
SYSTEMS|2472,2479
:|2479,2480
Per|2481,2484
HPI|2485,2488
.|2488,2489
Denies|2490,2496
headache|2497,2505
,|2505,2506
visual|2507,2513
changes|2514,2521
,|2521,2522
<EOL>|2523,2524
pharyngitis|2524,2535
,|2535,2536
rhinorrhea|2537,2547
,|2547,2548
nasal|2549,2554
congestion|2555,2565
,|2565,2566
cough|2567,2572
,|2572,2573
fevers|2574,2580
,|2580,2581
<EOL>|2582,2583
chills|2583,2589
,|2589,2590
sweats|2591,2597
,|2597,2598
weight|2599,2605
loss|2606,2610
,|2610,2611
dyspnea|2612,2619
,|2619,2620
chest|2621,2626
pain|2627,2631
,|2631,2632
abdominal|2633,2642
<EOL>|2643,2644
pain|2644,2648
,|2648,2649
nausea|2650,2656
,|2656,2657
vomiting|2658,2666
,|2666,2667
diarrhea|2668,2676
,|2676,2677
constipation|2678,2690
,|2690,2691
hematochezia|2692,2704
,|2704,2705
<EOL>|2706,2707
dysuria|2707,2714
,|2714,2715
rash|2716,2720
,|2720,2721
paresthesias|2722,2734
,|2734,2735
and|2736,2739
weakness|2740,2748
.|2748,2749
<EOL>|2749,2750
<EOL>|2751,2752
-|2774,2775
COPD|2776,2780
/|2780,2781
Asthma|2781,2787
on|2788,2790
home|2791,2795
2L|2796,2798
O2|2799,2801
<EOL>|2801,2802
-|2802,2803
Atypical|2804,2812
Chest|2813,2818
Pain|2819,2823
<EOL>|2823,2824
-|2824,2825
Hypertension|2826,2838
<EOL>|2838,2839
-|2839,2840
Hyperlipidemia|2841,2855
<EOL>|2855,2856
-|2856,2857
Osteroarthritis|2858,2873
<EOL>|2873,2874
-|2874,2875
Atrial|2876,2882
Fibrillation|2883,2895
on|2896,2898
Apixaban|2899,2907
<EOL>|2907,2908
-|2908,2909
Anxiety|2910,2917
<EOL>|2917,2918
-|2918,2919
Cervical|2920,2928
Radiculitis|2929,2940
<EOL>|2940,2941
-|2941,2942
Cervical|2943,2951
Spondylosis|2952,2963
<EOL>|2963,2964
-|2964,2965
Coronary|2966,2974
Artery|2975,2981
Disease|2982,2989
<EOL>|2989,2990
-|2990,2991
Headache|2992,3000
<EOL>|3000,3001
-|3001,3002
Herpes|3003,3009
Zoster|3010,3016
<EOL>|3016,3017
-|3017,3018
GI|3019,3021
Bleeding|3022,3030
<EOL>|3030,3031
-|3031,3032
Peripheral|3033,3043
Vascular|3044,3052
Disease|3053,3060
s|3061,3062
/|3062,3063
p|3063,3064
bilateral|3065,3074
iliac|3075,3080
stents|3081,3087
<EOL>|3087,3088
-|3088,3089
s|3090,3091
/|3091,3092
p|3092,3093
hip|3094,3097
replacement|3098,3109
<EOL>|3109,3110
<EOL>|3111,3112
:|3126,3127
<EOL>|3127,3128
_|3128,3129
_|3129,3130
_|3130,3131
<EOL>|3131,3132
:|3146,3147
<EOL>|3147,3148
Mother|3148,3154
with|3155,3159
asthma|3160,3166
and|3167,3170
hypertension|3171,3183
.|3183,3184
Father|3185,3191
with|3192,3196
colon|3197,3202
cancer|3203,3209
.|3209,3210
<EOL>|3211,3212
Brother|3212,3219
with|3220,3224
leukemia|3225,3233
.|3233,3234
<EOL>|3234,3235
<EOL>|3235,3236
<EOL>|3237,3238
PHYSICAL|3253,3261
EXAMINATION|3262,3273
ON|3274,3276
ADMISSION|3277,3286
:|3286,3287
<EOL>|3287,3288
=|3288,3289
=|3289,3290
=|3290,3291
=|3291,3292
=|3292,3293
=|3293,3294
=|3294,3295
=|3295,3296
=|3296,3297
=|3297,3298
=|3298,3299
=|3299,3300
=|3300,3301
=|3301,3302
=|3302,3303
=|3303,3304
=|3304,3305
=|3305,3306
=|3306,3307
=|3307,3308
=|3308,3309
=|3309,3310
=|3310,3311
=|3311,3312
=|3312,3313
=|3313,3314
=|3314,3315
=|3315,3316
=|3316,3317
=|3317,3318
=|3318,3319
=|3319,3320
=|3320,3321
=|3321,3322
<EOL>|3322,3323
VITALS|3323,3329
:|3329,3330
98.1|3331,3335
139|3336,3339
/|3339,3340
79|3340,3342
78|3343,3345
22|3346,3348
98RA|3349,3353
<EOL>|3355,3356
GENERAL|3356,3363
:|3363,3364
Pleasant|3365,3373
,|3373,3374
well|3375,3379
-|3379,3380
appearing|3380,3389
,|3389,3390
in|3391,3393
no|3394,3396
apparent|3397,3405
distress|3406,3414
.|3414,3415
<EOL>|3417,3418
HEENT|3418,3423
-|3424,3425
normocephalic|3426,3439
,|3439,3440
atraumatic|3441,3451
,|3451,3452
no|3453,3455
conjunctival|3456,3468
pallor|3469,3475
or|3476,3478
<EOL>|3479,3480
scleral|3480,3487
icterus|3488,3495
,|3495,3496
PERRLA|3497,3503
,|3503,3504
EOMI|3505,3509
,|3509,3510
OP|3511,3513
clear|3514,3519
.|3519,3520
<EOL>|3522,3523
NECK|3523,3527
:|3527,3528
Supple|3529,3535
,|3535,3536
no|3537,3539
LAD|3540,3543
,|3543,3544
no|3545,3547
thyromegaly|3548,3559
,|3559,3560
JVP|3561,3564
flat|3565,3569
.|3569,3570
<EOL>|3572,3573
CARDIAC|3573,3580
:|3580,3581
Normal|3582,3588
S1|3589,3591
/|3591,3592
S2|3592,3594
,|3594,3595
no|3596,3598
murmurs|3599,3606
rubs|3607,3611
or|3612,3614
gallops|3615,3622
.|3622,3623
<EOL>|3625,3626
PULMONARY|3626,3635
:|3635,3636
Inspiratory|3637,3648
and|3649,3652
expiratory|3653,3663
wheezes|3664,3671
in|3672,3674
all|3675,3678
lung|3679,3683
fields|3684,3690
<EOL>|3691,3692
<EOL>|3693,3694
ABDOMEN|3694,3701
:|3701,3702
Normal|3703,3709
bowel|3710,3715
sounds|3716,3722
,|3722,3723
soft|3724,3728
,|3728,3729
non-tender|3730,3740
,|3740,3741
non-distended|3742,3755
,|3755,3756
<EOL>|3757,3758
no|3758,3760
organomegaly|3761,3773
.|3773,3774
<EOL>|3776,3777
EXTREMITIES|3777,3788
:|3788,3789
Warm|3790,3794
,|3794,3795
well|3796,3800
-|3800,3801
perfused|3801,3809
,|3809,3810
no|3811,3813
cyanosis|3814,3822
,|3822,3823
clubbing|3824,3832
or|3833,3835
<EOL>|3836,3837
edema|3837,3842
.|3842,3843
<EOL>|3845,3846
SKIN|3846,3850
:|3850,3851
Without|3852,3859
rash|3860,3864
.|3864,3865
<EOL>|3867,3868
NEUROLOGIC|3868,3878
:|3878,3879
A|3880,3881
&|3881,3882
Ox3|3882,3885
,|3885,3886
CN|3887,3889
II|3890,3892
-|3892,3893
XII|3893,3896
grossly|3897,3904
normal|3905,3911
,|3911,3912
normal|3913,3919
sensation|3920,3929
,|3929,3930
<EOL>|3931,3932
with|3932,3936
strength|3937,3945
_|3946,3947
_|3947,3948
_|3948,3949
throughout|3950,3960
.|3960,3961
<EOL>|3963,3964
<EOL>|3964,3965
PHYSICAL|3965,3973
EXAMINATION|3974,3985
ON|3986,3988
DISCHARGE|3989,3998
:|3998,3999
<EOL>|3999,4000
=|4000,4001
=|4001,4002
=|4002,4003
=|4003,4004
=|4004,4005
=|4005,4006
=|4006,4007
=|4007,4008
=|4008,4009
=|4009,4010
=|4010,4011
=|4011,4012
=|4012,4013
=|4013,4014
=|4014,4015
=|4015,4016
=|4016,4017
=|4017,4018
=|4018,4019
=|4019,4020
=|4020,4021
=|4021,4022
=|4022,4023
=|4023,4024
=|4024,4025
=|4025,4026
=|4026,4027
=|4027,4028
=|4028,4029
=|4029,4030
=|4030,4031
=|4031,4032
=|4032,4033
=|4033,4034
<EOL>|4034,4035
VITALS|4035,4041
:|4041,4042
98.2|4043,4047
130|4048,4051
-|4051,4052
140|4052,4055
/|4055,4056
70'S|4056,4060
70|4061,4063
-|4063,4064
80's|4064,4068
20|4069,4071
98RA|4073,4077
<EOL>|4079,4080
GENERAL|4080,4087
:|4087,4088
Pleasant|4089,4097
,|4097,4098
well|4099,4103
-|4103,4104
appearing|4104,4113
,|4113,4114
in|4115,4117
no|4118,4120
apparent|4121,4129
distress|4130,4138
.|4138,4139
<EOL>|4141,4142
HEENT|4142,4147
-|4148,4149
normocephalic|4150,4163
,|4163,4164
atraumatic|4165,4175
,|4175,4176
no|4177,4179
conjunctival|4180,4192
pallor|4193,4199
or|4200,4202
<EOL>|4203,4204
scleral|4204,4211
icterus|4212,4219
,|4219,4220
PERRLA|4221,4227
,|4227,4228
EOMI|4229,4233
,|4233,4234
OP|4235,4237
clear|4238,4243
.|4243,4244
<EOL>|4246,4247
NECK|4247,4251
:|4251,4252
Supple|4253,4259
,|4259,4260
no|4261,4263
LAD|4264,4267
,|4267,4268
no|4269,4271
thyromegaly|4272,4283
,|4283,4284
JVP|4285,4288
flat|4289,4293
.|4293,4294
<EOL>|4296,4297
CARDIAC|4297,4304
:|4304,4305
Normal|4306,4312
S1|4313,4315
/|4315,4316
S2|4316,4318
,|4318,4319
no|4320,4322
murmurs|4323,4330
rubs|4331,4335
or|4336,4338
gallops|4339,4346
.|4346,4347
<EOL>|4349,4350
PULMONARY|4350,4359
:|4359,4360
Decreased|4361,4370
inspiratory|4371,4382
and|4383,4386
expiratory|4387,4397
wheezes|4398,4405
in|4406,4408
all|4409,4412
<EOL>|4413,4414
lung|4414,4418
fields|4419,4425
<EOL>|4427,4428
ABDOMEN|4428,4435
:|4435,4436
Normal|4437,4443
bowel|4444,4449
sounds|4450,4456
,|4456,4457
soft|4458,4462
,|4462,4463
non-tender|4464,4474
,|4474,4475
non-distended|4476,4489
,|4489,4490
<EOL>|4491,4492
no|4492,4494
organomegaly|4495,4507
.|4507,4508
<EOL>|4510,4511
EXTREMITIES|4511,4522
:|4522,4523
Warm|4524,4528
,|4528,4529
well|4530,4534
-|4534,4535
perfused|4535,4543
,|4543,4544
no|4545,4547
cyanosis|4548,4556
,|4556,4557
clubbing|4558,4566
or|4567,4569
<EOL>|4570,4571
edema|4571,4576
.|4576,4577
<EOL>|4579,4580
SKIN|4580,4584
:|4584,4585
Without|4586,4593
rash|4594,4598
.|4598,4599
<EOL>|4601,4602
NEUROLOGIC|4602,4612
:|4612,4613
A|4614,4615
&|4615,4616
Ox3|4616,4619
,|4619,4620
CN|4621,4623
II|4624,4626
-|4626,4627
XII|4627,4630
grossly|4631,4638
normal|4639,4645
,|4645,4646
normal|4647,4653
sensation|4654,4663
,|4663,4664
<EOL>|4665,4666
with|4666,4670
strength|4671,4679
_|4680,4681
_|4681,4682
_|4682,4683
throughout|4684,4694
.|4694,4695
<EOL>|4697,4698
<EOL>|4698,4699
<EOL>|4700,4701
Pertinent|4701,4710
Results|4711,4718
:|4718,4719
<EOL>|4719,4720
LABS|4720,4724
ON|4725,4727
ADMISSION|4728,4737
:|4737,4738
<EOL>|4738,4739
=|4739,4740
=|4740,4741
=|4741,4742
=|4742,4743
=|4743,4744
=|4744,4745
=|4745,4746
=|4746,4747
=|4747,4748
=|4748,4749
=|4749,4750
=|4750,4751
=|4751,4752
=|4752,4753
=|4753,4754
=|4754,4755
=|4755,4756
=|4756,4757
<EOL>|4757,4758
_|4758,4759
_|4759,4760
_|4760,4761
04|4762,4764
:|4764,4765
00PM|4765,4769
BLOOD|4770,4775
Neuts|4776,4781
-|4781,4782
92|4782,4784
.|4784,4785
1|4785,4786
*|4786,4787
Lymphs|4788,4794
-|4794,4795
4|4795,4796
.|4796,4797
5|4797,4798
*|4798,4799
Monos|4800,4805
-|4805,4806
2|4806,4807
.|4807,4808
7|4808,4809
*|4809,4810
<EOL>|4811,4812
Eos|4812,4815
-|4815,4816
0|4816,4817
.|4817,4818
0|4818,4819
*|4819,4820
Baso|4821,4825
-|4825,4826
0.0|4826,4829
Im|4830,4832
_|4833,4834
_|4834,4835
_|4835,4836
AbsNeut|4837,4844
-|4844,4845
5|4845,4846
.|4846,4847
51|4847,4849
AbsLymp|4850,4857
-|4857,4858
0|4858,4859
.|4859,4860
27|4860,4862
*|4862,4863
<EOL>|4864,4865
AbsMono|4865,4872
-|4872,4873
0|4873,4874
.|4874,4875
16|4875,4877
*|4877,4878
AbsEos|4879,4885
-|4885,4886
0|4886,4887
.|4887,4888
00|4888,4890
*|4890,4891
AbsBaso|4892,4899
-|4899,4900
0|4900,4901
.|4901,4902
00|4902,4904
*|4904,4905
<EOL>|4905,4906
_|4906,4907
_|4907,4908
_|4908,4909
04|4910,4912
:|4912,4913
00PM|4913,4917
BLOOD|4918,4923
Plt|4924,4927
_|4928,4929
_|4929,4930
_|4930,4931
<EOL>|4931,4932
_|4932,4933
_|4933,4934
_|4934,4935
04|4936,4938
:|4938,4939
00PM|4939,4943
BLOOD|4944,4949
Glucose|4950,4957
-|4957,4958
140|4958,4961
*|4961,4962
UreaN|4963,4968
-|4968,4969
17|4969,4971
Creat|4972,4977
-|4977,4978
1.0|4978,4981
Na|4982,4984
-|4984,4985
136|4985,4988
<EOL>|4989,4990
K|4990,4991
-|4991,4992
3.5|4992,4995
Cl|4996,4998
-|4998,4999
95|4999,5001
*|5001,5002
HCO3|5003,5007
-|5007,5008
29|5008,5010
AnGap|5011,5016
-|5016,5017
16|5017,5019
<EOL>|5019,5020
_|5020,5021
_|5021,5022
_|5022,5023
04|5024,5026
:|5026,5027
00PM|5027,5031
BLOOD|5032,5037
proBNP|5038,5044
-|5044,5045
254|5045,5048
<EOL>|5048,5049
_|5049,5050
_|5050,5051
_|5051,5052
03|5053,5055
:|5055,5056
58PM|5056,5060
BLOOD|5061,5066
_|5067,5068
_|5068,5069
_|5069,5070
pO2|5071,5074
-|5074,5075
59|5075,5077
*|5077,5078
pCO2|5079,5083
-|5083,5084
43|5084,5086
pH|5087,5089
-|5089,5090
7.45|5090,5094
<EOL>|5095,5096
calTCO2|5096,5103
-|5103,5104
31|5104,5106
*|5106,5107
Base|5108,5112
XS|5113,5115
-|5115,5116
4|5116,5117
<EOL>|5117,5118
<EOL>|5118,5119
LABS|5119,5123
ON|5124,5126
DISCHARGE|5127,5136
:|5136,5137
<EOL>|5137,5138
=|5138,5139
=|5139,5140
=|5140,5141
=|5141,5142
=|5142,5143
=|5143,5144
=|5144,5145
=|5145,5146
=|5146,5147
=|5147,5148
=|5148,5149
=|5149,5150
=|5150,5151
=|5151,5152
=|5152,5153
=|5153,5154
=|5154,5155
=|5155,5156
<EOL>|5156,5157
_|5157,5158
_|5158,5159
_|5159,5160
08|5161,5163
:|5163,5164
00AM|5164,5168
BLOOD|5169,5174
WBC|5175,5178
-|5178,5179
5.8|5179,5182
RBC|5183,5186
-|5186,5187
4|5187,5188
.|5188,5189
37|5189,5191
Hgb|5192,5195
-|5195,5196
11.9|5196,5200
Hct|5201,5204
-|5204,5205
38.2|5205,5209
MCV|5210,5213
-|5213,5214
87|5214,5216
<EOL>|5217,5218
MCH|5218,5221
-|5221,5222
27.2|5222,5226
MCHC|5227,5231
-|5231,5232
31|5232,5234
.|5234,5235
2|5235,5236
*|5236,5237
RDW|5238,5241
-|5241,5242
20|5242,5244
.|5244,5245
4|5245,5246
*|5246,5247
RDWSD|5248,5253
-|5253,5254
65|5254,5256
.|5256,5257
6|5257,5258
*|5258,5259
Plt|5260,5263
_|5264,5265
_|5265,5266
_|5266,5267
<EOL>|5267,5268
_|5268,5269
_|5269,5270
_|5270,5271
08|5272,5274
:|5274,5275
00AM|5275,5279
BLOOD|5280,5285
Plt|5286,5289
_|5290,5291
_|5291,5292
_|5292,5293
<EOL>|5293,5294
_|5294,5295
_|5295,5296
_|5296,5297
08|5298,5300
:|5300,5301
00AM|5301,5305
BLOOD|5306,5311
Glucose|5312,5319
-|5319,5320
156|5320,5323
*|5323,5324
UreaN|5325,5330
-|5330,5331
21|5331,5333
*|5333,5334
Creat|5335,5340
-|5340,5341
0.9|5341,5344
Na|5345,5347
-|5347,5348
134|5348,5351
<EOL>|5352,5353
K|5353,5354
-|5354,5355
3.4|5355,5358
Cl|5359,5361
-|5361,5362
92|5362,5364
*|5364,5365
HCO3|5366,5370
-|5370,5371
30|5371,5373
AnGap|5374,5379
-|5379,5380
15|5380,5382
<EOL>|5382,5383
_|5383,5384
_|5384,5385
_|5385,5386
08|5387,5389
:|5389,5390
00AM|5390,5394
BLOOD|5395,5400
Calcium|5401,5408
-|5408,5409
9.7|5409,5412
Phos|5413,5417
-|5417,5418
3.6|5418,5421
Mg|5422,5424
-|5424,5425
2.0|5425,5428
<EOL>|5428,5429
<EOL>|5429,5430
STUDIES|5430,5437
:|5437,5438
<EOL>|5438,5439
=|5439,5440
=|5440,5441
=|5441,5442
=|5442,5443
=|5443,5444
=|5444,5445
=|5445,5446
=|5446,5447
<EOL>|5447,5448
CXR|5448,5451
_|5452,5453
_|5453,5454
_|5454,5455
:|5455,5456
No|5457,5459
acute|5460,5465
cardiopulmonary|5466,5481
process|5482,5489
<EOL>|5491,5492
EKG|5492,5495
:|5495,5496
NSR|5497,5500
rate|5501,5505
72|5506,5508
,|5508,5509
QTC|5510,5513
469|5514,5517
,|5517,5518
LBBB|5519,5523
<EOL>|5523,5524
<EOL>|5525,5526
_|5549,5550
_|5550,5551
_|5551,5552
yo|5553,5555
F|5556,5557
with|5558,5562
history|5563,5570
of|5571,5573
COPD|5574,5578
on|5579,5581
home|5582,5586
O2|5587,5589
,|5589,5590
atrial|5591,5597
fibrillation|5598,5610
on|5611,5613
<EOL>|5614,5615
apixaban|5615,5623
,|5623,5624
hypertension|5625,5637
,|5637,5638
CAD|5639,5642
,|5642,5643
hyperlipidemia|5644,5658
,|5658,5659
and|5660,5663
recurrent|5664,5673
<EOL>|5674,5675
hospitalization|5675,5690
for|5691,5694
COPD|5695,5699
exacerbation|5700,5712
over|5713,5717
the|5718,5721
last|5722,5726
4|5727,5728
months|5729,5735
,|5735,5736
<EOL>|5737,5738
who|5738,5741
presented|5742,5751
with|5752,5756
dyspnea|5757,5764
consistent|5765,5775
with|5776,5780
COPD|5781,5785
exacerbation|5786,5798
,|5798,5799
<EOL>|5800,5801
possibly|5801,5809
secondary|5810,5819
to|5820,5822
acute|5823,5828
viral|5829,5834
URI|5835,5838
with|5839,5843
concurrent|5844,5854
sinusitis|5855,5864
<EOL>|5865,5866
/|5866,5867
Eustachian|5868,5878
tube|5879,5883
dysfunction|5884,5895
<EOL>|5895,5896
<EOL>|5896,5897
#|5897,5898
COPD|5899,5903
exacerbation|5904,5916
:|5916,5917
<EOL>|5919,5920
Patient|5920,5927
has|5928,5931
been|5932,5936
experiencing|5937,5949
recurrent|5950,5959
COPD|5960,5964
exacerbations|5965,5978
over|5979,5983
<EOL>|5984,5985
the|5985,5988
last|5989,5993
4|5994,5995
months|5996,6002
.|6002,6003
She|6004,6007
presented|6008,6017
with|6018,6022
dyspnea|6023,6030
consistent|6031,6041
with|6042,6046
<EOL>|6047,6048
COPD|6048,6052
exacerbation|6053,6065
,|6065,6066
possibly|6067,6075
secondary|6076,6085
to|6086,6088
acute|6089,6094
viral|6095,6100
URI|6101,6104
with|6105,6109
<EOL>|6110,6111
concurrent|6111,6121
sinusitis|6122,6131
/|6132,6133
Eustachian|6134,6144
tube|6145,6149
dysfunction|6150,6161
.|6161,6162
We|6163,6165
continued|6166,6175
<EOL>|6176,6177
home|6177,6181
spiriva|6182,6189
,|6189,6190
theophylline|6191,6203
,|6203,6204
and|6205,6208
advair|6209,6215
.|6215,6216
We|6217,6219
continued|6220,6229
her|6230,6233
steroid|6234,6241
<EOL>|6242,6243
therapy|6243,6250
at|6251,6253
30mg|6254,6258
prednisone|6259,6269
daily|6270,6275
with|6276,6280
a|6281,6282
slow|6283,6287
taper|6288,6293
(|6294,6295
5mg|6295,6298
every|6299,6304
2|6305,6306
<EOL>|6307,6308
weeks|6308,6313
)|6313,6314
.|6314,6315
We|6316,6318
also|6319,6323
treated|6324,6331
her|6332,6335
with|6336,6340
levofloxacin|6341,6353
(|6354,6355
Day|6355,6358
_|6359,6360
_|6360,6361
_|6361,6362
<EOL>|6363,6364
with|6364,6368
plan|6369,6373
for|6374,6377
5|6378,6379
-|6379,6380
day|6380,6383
course|6384,6390
given|6391,6396
COPD|6397,6401
exacerbation|6402,6414
with|6415,6419
<EOL>|6420,6421
concurrent|6421,6431
concern|6432,6439
for|6440,6443
sinusitis|6444,6453
/|6454,6455
bulging|6456,6463
right|6464,6469
tympanic|6470,6478
<EOL>|6479,6480
membrane|6480,6488
.|6488,6489
<EOL>|6489,6490
<EOL>|6490,6491
CHRONIC|6491,6498
ISSUES|6499,6505
:|6505,6506
<EOL>|6508,6509
=|6509,6510
=|6510,6511
=|6511,6512
=|6512,6513
=|6513,6514
=|6514,6515
=|6515,6516
=|6516,6517
=|6517,6518
=|6518,6519
=|6519,6520
=|6520,6521
=|6521,6522
=|6522,6523
=|6523,6524
=|6524,6525
=|6525,6526
=|6526,6527
<EOL>|6529,6530
#|6530,6531
Anxiety|6532,6539
/|6539,6540
Insomnia|6540,6548
:|6548,6549
We|6550,6552
continued|6553,6562
home|6563,6567
lorazepam|6568,6577
.|6577,6578
<EOL>|6580,6581
<EOL>|6581,6582
#|6582,6583
Atrial|6584,6590
Fibrillation|6591,6603
:|6603,6604
We|6605,6607
continued|6608,6617
diltiazem|6618,6627
for|6628,6631
rate|6632,6636
control|6637,6644
<EOL>|6645,6646
and|6646,6649
apixaban|6650,6658
for|6659,6662
anticoagulation|6663,6678
.|6678,6679
<EOL>|6679,6680
<EOL>|6681,6682
#|6682,6683
Hypertension|6684,6696
:|6696,6697
We|6698,6700
continued|6701,6710
home|6711,6715
imdur|6716,6721
,|6721,6722
hydrochlorothiazide|6723,6742
,|6742,6743
<EOL>|6744,6745
and|6745,6748
diltiazem|6749,6758
.|6758,6759
<EOL>|6761,6762
<EOL>|6763,6764
#|6764,6765
CAD|6766,6769
:|6769,6770
Cardiac|6771,6778
catheterization|6779,6794
in|6795,6797
_|6798,6799
_|6799,6800
_|6800,6801
without|6802,6809
evidence|6810,6818
of|6819,6821
<EOL>|6822,6823
significant|6823,6834
stenosis|6835,6843
of|6844,6846
coronaries|6847,6857
.|6857,6858
ECHO|6859,6863
on|6864,6866
_|6867,6868
_|6868,6869
_|6869,6870
with|6871,6875
EF|6876,6878
>|6879,6880
<EOL>|6881,6882
55|6882,6884
%|6884,6885
and|6886,6889
no|6890,6892
regional|6893,6901
or|6902,6904
global|6905,6911
wall|6912,6916
motion|6917,6923
abnormalities|6924,6937
.|6937,6938
We|6939,6941
<EOL>|6942,6943
continued|6943,6952
home|6953,6957
aspirin|6958,6965
and|6966,6969
atorvastatin|6970,6982
.|6982,6983
<EOL>|6985,6986
<EOL>|6987,6988
#|6988,6989
Anemia|6990,6996
:|6996,6997
We|6998,7000
continued|7001,7010
home|7011,7015
iron|7016,7020
supplements|7021,7032
.|7032,7033
<EOL>|7033,7034
<EOL>|7034,7035
*|7035,7036
*|7036,7037
*|7037,7038
TRANSITIONAL|7038,7050
ISSUES|7051,7057
:|7057,7058
*|7058,7059
*|7059,7060
*|7060,7061
<EOL>|7062,7063
-|7063,7064
Continue|7065,7073
levofloxacin|7074,7086
with|7087,7091
plan|7092,7096
for|7097,7100
5|7101,7102
-|7102,7103
day|7103,7106
course|7107,7113
(|7114,7115
Day|7115,7118
<EOL>|7119,7120
_|7120,7121
_|7121,7122
_|7122,7123
end|7124,7127
_|7128,7129
_|7129,7130
_|7130,7131
<EOL>|7131,7132
-|7132,7133
Patient|7134,7141
was|7142,7145
started|7146,7153
Bactrim|7154,7161
PPX|7162,7165
(|7166,7167
1|7167,7168
tab|7169,7172
SS|7173,7175
daily|7176,7181
)|7181,7182
given|7183,7188
<EOL>|7189,7190
extended|7190,7198
courses|7199,7206
of|7207,7209
steroids|7210,7218
,|7218,7219
stop|7220,7224
after|7225,7230
discontinuation|7231,7246
of|7247,7249
<EOL>|7250,7251
steroids|7251,7259
<EOL>|7259,7260
-|7260,7261
Patient|7262,7269
was|7270,7273
discharged|7274,7284
on|7285,7287
prednisone|7288,7298
30|7299,7301
mg|7302,7304
with|7305,7309
plan|7310,7314
for|7315,7318
taper|7319,7324
<EOL>|7325,7326
by|7326,7328
5mg|7329,7332
every|7333,7338
2|7339,7340
weeks|7341,7346
:|7346,7347
<EOL>|7347,7348
Prednisone|7349,7359
30|7360,7362
mg|7363,7365
for|7366,7369
two|7370,7373
weeks|7374,7379
(|7380,7381
Day|7381,7384
1|7385,7386
=|7386,7387
_|7388,7389
_|7389,7390
_|7390,7391
end|7392,7395
<EOL>|7396,7397
_|7397,7398
_|7398,7399
_|7399,7400
<EOL>|7400,7401
Prednisone|7402,7412
25|7413,7415
mg|7416,7418
for|7419,7422
two|7423,7426
weeks|7427,7432
(|7433,7434
Day|7434,7437
1|7438,7439
=|7439,7440
_|7441,7442
_|7442,7443
_|7443,7444
end|7445,7448
<EOL>|7449,7450
_|7450,7451
_|7451,7452
_|7452,7453
<EOL>|7453,7454
Prednisone|7455,7465
20|7466,7468
mg|7469,7471
for|7472,7475
two|7476,7479
weeks|7480,7485
(|7486,7487
Day|7487,7490
1|7491,7492
=|7492,7493
_|7494,7495
_|7495,7496
_|7496,7497
end|7498,7501
<EOL>|7502,7503
_|7503,7504
_|7504,7505
_|7505,7506
<EOL>|7506,7507
etc|7508,7511
...|7511,7514
<EOL>|7514,7515
#|7515,7516
CONTACT|7517,7524
:|7524,7525
_|7526,7527
_|7527,7528
_|7528,7529
(|7530,7531
husband|7531,7538
/|7538,7539
HCP|7539,7542
)|7542,7543
_|7544,7545
_|7545,7546
_|7546,7547
<EOL>|7548,7549
#|7549,7550
CODE|7551,7555
STATUS|7556,7562
:|7562,7563
Full|7564,7568
confirmed|7569,7578
<EOL>|7579,7580
<EOL>|7581,7582
Medications|7582,7593
on|7594,7596
Admission|7597,7606
:|7606,7607
<EOL>|7607,7608
The|7608,7611
Preadmission|7612,7624
Medication|7625,7635
list|7636,7640
is|7641,7643
accurate|7644,7652
and|7653,7656
complete|7657,7665
.|7665,7666
<EOL>|7666,7667
1.|7667,7669
Acetaminophen|7670,7683
325|7684,7687
mg|7688,7690
PO|7691,7693
Q4H|7694,7697
:|7697,7698
PRN|7698,7701
Pain|7702,7706
<EOL>|7707,7708
2.|7708,7710
albuterol|7711,7720
sulfate|7721,7728
90|7729,7731
mcg|7732,7735
/|7735,7736
actuation|7736,7745
inhalation|7746,7756
Q4H|7757,7760
<EOL>|7761,7762
3.|7762,7764
Apixaban|7765,7773
5|7774,7775
mg|7776,7778
PO|7779,7781
BID|7782,7785
<EOL>|7786,7787
4.|7787,7789
Aspirin|7790,7797
81|7798,7800
mg|7801,7803
PO|7804,7806
DAILY|7807,7812
<EOL>|7813,7814
5.|7814,7816
Atorvastatin|7817,7829
10|7830,7832
mg|7833,7835
PO|7836,7838
QPM|7839,7842
<EOL>|7843,7844
6.|7844,7846
Diltiazem|7847,7856
Extended|7857,7865
-|7865,7866
Release|7866,7873
240|7874,7877
mg|7878,7880
PO|7881,7883
BID|7884,7887
<EOL>|7888,7889
7.|7889,7891
Docusate|7892,7900
Sodium|7901,7907
100|7908,7911
mg|7912,7914
PO|7915,7917
BID|7918,7921
<EOL>|7922,7923
8.|7923,7925
Dorzolamide|7926,7937
2|7938,7939
%|7939,7940
Ophth|7941,7946
.|7946,7947
Soln.|7948,7953
1|7954,7955
DROP|7956,7960
BOTH|7961,7965
EYES|7966,7970
BID|7971,7974
<EOL>|7975,7976
9.|7976,7978
Ferrous|7979,7986
Sulfate|7987,7994
325|7995,7998
mg|7999,8001
PO|8002,8004
DAILY|8005,8010
<EOL>|8011,8012
10.|8012,8015
Fluticasone|8016,8027
Propionate|8028,8038
NASAL|8039,8044
2|8045,8046
SPRY|8047,8051
NU|8052,8054
DAILY|8055,8060
:|8060,8061
PRN|8061,8064
allergies|8065,8074
<EOL>|8075,8076
11|8076,8078
.|8078,8079
Fluticasone|8080,8091
-|8091,8092
Salmeterol|8092,8102
Diskus|8103,8109
(|8110,8111
500|8111,8114
/|8114,8115
50|8115,8117
)|8117,8118
1|8120,8121
INH|8122,8125
IH|8126,8128
BID|8129,8132
<EOL>|8133,8134
12.|8134,8137
Guaifenesin|8138,8149
_|8150,8151
_|8151,8152
_|8152,8153
mL|8154,8156
PO|8157,8159
Q4H|8160,8163
:|8163,8164
PRN|8164,8167
cough|8168,8173
<EOL>|8174,8175
13.|8175,8178
Hydrochlorothiazide|8179,8198
50|8199,8201
mg|8202,8204
PO|8205,8207
DAILY|8208,8213
<EOL>|8214,8215
14.|8215,8218
Isosorbide|8219,8229
Mononitrate|8230,8241
(|8242,8243
Extended|8243,8251
Release|8252,8259
)|8259,8260
240|8261,8264
mg|8265,8267
PO|8268,8270
DAILY|8271,8276
<EOL>|8277,8278
15.|8278,8281
Latanoprost|8282,8293
0.005|8294,8299
%|8299,8300
Ophth|8301,8306
.|8306,8307
Soln.|8308,8313
1|8314,8315
DROP|8316,8320
BOTH|8321,8325
EYES|8326,8330
QHS|8331,8334
<EOL>|8335,8336
16|8336,8338
.|8338,8339
Lorazepam|8340,8349
0.5|8350,8353
mg|8354,8356
PO|8357,8359
Q8H|8360,8363
:|8363,8364
PRN|8364,8367
Insomnia|8368,8376
,|8376,8377
anxiety|8378,8385
,|8385,8386
vertigo|8387,8394
<EOL>|8395,8396
17.|8396,8399
Multivitamins|8400,8413
1|8414,8415
TAB|8416,8419
PO|8420,8422
DAILY|8423,8428
<EOL>|8429,8430
18.|8430,8433
Ranitidine|8434,8444
300|8445,8448
mg|8449,8451
PO|8452,8454
DAILY|8455,8460
<EOL>|8461,8462
19|8462,8464
.|8464,8465
Theophylline|8466,8478
SR|8479,8481
300|8482,8485
mg|8486,8488
PO|8489,8491
BID|8492,8495
<EOL>|8496,8497
20|8497,8499
.|8499,8500
Tiotropium|8501,8511
Bromide|8512,8519
1|8520,8521
CAP|8522,8525
IH|8526,8528
DAILY|8529,8534
<EOL>|8535,8536
21|8536,8538
.|8538,8539
Calcitrate|8540,8550
-|8550,8551
Vitamin|8551,8558
D|8559,8560
(|8561,8562
calcium|8562,8569
citrate|8570,8577
-|8577,8578
vitamin|8578,8585
D3|8586,8588
)|8588,8589
315|8590,8593
mg|8594,8596
-|8597,8598
<EOL>|8599,8600
200|8600,8603
units|8604,8609
oral|8611,8615
DAILY|8616,8621
<EOL>|8622,8623
22.|8623,8626
cod|8627,8630
liver|8631,8636
oil|8637,8640
1|8641,8642
capsule|8643,8650
oral|8652,8656
BID|8657,8660
<EOL>|8661,8662
23|8662,8664
.|8664,8665
Ipratropium|8666,8677
Bromide|8678,8685
Neb|8686,8689
1|8690,8691
NEB|8692,8695
IH|8696,8698
Q6H|8699,8702
:|8702,8703
PRN|8703,8706
Wheezing|8707,8715
<EOL>|8716,8717
24|8717,8719
.|8719,8720
PredniSONE|8721,8731
30|8732,8734
mg|8735,8737
PO|8738,8740
DAILY|8741,8746
<EOL>|8747,8748
Tapered|8748,8755
dose|8756,8760
-|8761,8762
DOWN|8763,8767
<EOL>|8768,8769
<EOL>|8769,8770
<EOL>|8771,8772
Discharge|8772,8781
Medications|8782,8793
:|8793,8794
<EOL>|8794,8795
1.|8795,8797
Acetaminophen|8798,8811
325|8812,8815
mg|8816,8818
PO|8819,8821
Q4H|8822,8825
:|8825,8826
PRN|8826,8829
Pain|8830,8834
<EOL>|8835,8836
2.|8836,8838
albuterol|8839,8848
sulfate|8849,8856
90|8857,8859
mcg|8860,8863
/|8863,8864
actuation|8864,8873
inhalation|8874,8884
Q4H|8885,8888
<EOL>|8889,8890
3.|8890,8892
Apixaban|8893,8901
5|8902,8903
mg|8904,8906
PO|8907,8909
BID|8910,8913
<EOL>|8914,8915
4.|8915,8917
Aspirin|8918,8925
81|8926,8928
mg|8929,8931
PO|8932,8934
DAILY|8935,8940
<EOL>|8941,8942
5.|8942,8944
Atorvastatin|8945,8957
10|8958,8960
mg|8961,8963
PO|8964,8966
QPM|8967,8970
<EOL>|8971,8972
6.|8972,8974
Diltiazem|8975,8984
Extended|8985,8993
-|8993,8994
Release|8994,9001
240|9002,9005
mg|9006,9008
PO|9009,9011
BID|9012,9015
<EOL>|9016,9017
7.|9017,9019
Docusate|9020,9028
Sodium|9029,9035
100|9036,9039
mg|9040,9042
PO|9043,9045
BID|9046,9049
<EOL>|9050,9051
8.|9051,9053
Dorzolamide|9054,9065
2|9066,9067
%|9067,9068
Ophth|9069,9074
.|9074,9075
Soln.|9076,9081
1|9082,9083
DROP|9084,9088
BOTH|9089,9093
EYES|9094,9098
BID|9099,9102
<EOL>|9103,9104
9.|9104,9106
Ferrous|9107,9114
Sulfate|9115,9122
325|9123,9126
mg|9127,9129
PO|9130,9132
DAILY|9133,9138
<EOL>|9139,9140
10.|9140,9143
Fluticasone|9144,9155
Propionate|9156,9166
NASAL|9167,9172
2|9173,9174
SPRY|9175,9179
NU|9180,9182
DAILY|9183,9188
:|9188,9189
PRN|9189,9192
allergies|9193,9202
<EOL>|9203,9204
11|9204,9206
.|9206,9207
Fluticasone|9208,9219
-|9219,9220
Salmeterol|9220,9230
Diskus|9231,9237
(|9238,9239
500|9239,9242
/|9242,9243
50|9243,9245
)|9245,9246
1|9248,9249
INH|9250,9253
IH|9254,9256
BID|9257,9260
<EOL>|9261,9262
12.|9262,9265
Guaifenesin|9266,9277
_|9278,9279
_|9279,9280
_|9280,9281
mL|9282,9284
PO|9285,9287
Q4H|9288,9291
:|9291,9292
PRN|9292,9295
cough|9296,9301
<EOL>|9302,9303
13.|9303,9306
Hydrochlorothiazide|9307,9326
50|9327,9329
mg|9330,9332
PO|9333,9335
DAILY|9336,9341
<EOL>|9342,9343
14.|9343,9346
Isosorbide|9347,9357
Mononitrate|9358,9369
(|9370,9371
Extended|9371,9379
Release|9380,9387
)|9387,9388
240|9389,9392
mg|9393,9395
PO|9396,9398
DAILY|9399,9404
<EOL>|9405,9406
15.|9406,9409
Latanoprost|9410,9421
0.005|9422,9427
%|9427,9428
Ophth|9429,9434
.|9434,9435
Soln.|9436,9441
1|9442,9443
DROP|9444,9448
BOTH|9449,9453
EYES|9454,9458
QHS|9459,9462
<EOL>|9463,9464
16|9464,9466
.|9466,9467
Lorazepam|9468,9477
0.5|9478,9481
mg|9482,9484
PO|9485,9487
Q8H|9488,9491
:|9491,9492
PRN|9492,9495
Insomnia|9496,9504
,|9504,9505
anxiety|9506,9513
,|9513,9514
vertigo|9515,9522
<EOL>|9523,9524
17.|9524,9527
Multivitamins|9528,9541
1|9542,9543
TAB|9544,9547
PO|9548,9550
DAILY|9551,9556
<EOL>|9557,9558
18.|9558,9561
PredniSONE|9562,9572
30|9573,9575
mg|9576,9578
PO|9579,9581
DAILY|9582,9587
<EOL>|9588,9589
Please|9589,9595
decrease|9596,9604
dose|9605,9609
by|9610,9612
5mg|9613,9616
every|9617,9622
2|9623,9624
weeks|9625,9630
<EOL>|9631,9632
Tapered|9632,9639
dose|9640,9644
-|9645,9646
DOWN|9647,9651
<EOL>|9652,9653
RX|9653,9655
*|9656,9657
prednisone|9657,9667
10|9668,9670
mg|9671,9673
3|9674,9675
tablets|9676,9683
(|9683,9684
s|9684,9685
)|9685,9686
by|9687,9689
mouth|9690,9695
once|9696,9700
a|9701,9702
day|9703,9706
Disp|9707,9711
#|9712,9713
*|9713,9714
45|9714,9716
<EOL>|9717,9718
Dose|9718,9722
Pack|9723,9727
Refills|9728,9735
:|9735,9736
*|9736,9737
0|9737,9738
<EOL>|9738,9739
19|9739,9741
.|9741,9742
Ranitidine|9743,9753
300|9754,9757
mg|9758,9760
PO|9761,9763
DAILY|9764,9769
<EOL>|9770,9771
20|9771,9773
.|9773,9774
Theophylline|9775,9787
SR|9788,9790
300|9791,9794
mg|9795,9797
PO|9798,9800
BID|9801,9804
<EOL>|9805,9806
21|9806,9808
.|9808,9809
Tiotropium|9810,9820
Bromide|9821,9828
1|9829,9830
CAP|9831,9834
IH|9835,9837
DAILY|9838,9843
<EOL>|9844,9845
22.|9845,9848
Levofloxacin|9849,9861
750|9862,9865
mg|9866,9868
PO|9869,9871
DAILY|9872,9877
Duration|9878,9886
:|9886,9887
5|9888,9889
Days|9890,9894
<EOL>|9895,9896
RX|9896,9898
*|9899,9900
levofloxacin|9900,9912
750|9913,9916
mg|9917,9919
1|9920,9921
tablet|9922,9928
(|9928,9929
s|9929,9930
)|9930,9931
by|9932,9934
mouth|9935,9940
once|9941,9945
a|9946,9947
day|9948,9951
Disp|9952,9956
#|9957,9958
*|9958,9959
4|9959,9960
<EOL>|9961,9962
Tablet|9962,9968
Refills|9969,9976
:|9976,9977
*|9977,9978
0|9978,9979
<EOL>|9979,9980
23|9980,9982
.|9982,9983
Sulfameth|9984,9993
/|9993,9994
Trimethoprim|9994,10006
SS|10007,10009
1|10010,10011
TAB|10012,10015
PO|10016,10018
DAILY|10019,10024
prophylaxis|10025,10036
for|10037,10040
<EOL>|10041,10042
long|10042,10046
term|10047,10051
steroid|10052,10059
use|10060,10063
<EOL>|10064,10065
RX|10065,10067
*|10068,10069
sulfamethoxazole|10069,10085
-|10085,10086
trimethoprim|10086,10098
400|10099,10102
mg|10103,10105
-|10105,10106
80|10106,10108
mg|10109,10111
1|10112,10113
tablet|10114,10120
(|10120,10121
s|10121,10122
)|10122,10123
by|10124,10126
<EOL>|10127,10128
mouth|10128,10133
once|10134,10138
a|10139,10140
day|10141,10144
Disp|10145,10149
#|10150,10151
*|10151,10152
30|10152,10154
Tablet|10155,10161
Refills|10162,10169
:|10169,10170
*|10170,10171
0|10171,10172
<EOL>|10172,10173
24|10173,10175
.|10175,10176
Calcitrate|10177,10187
-|10187,10188
Vitamin|10188,10195
D|10196,10197
(|10198,10199
calcium|10199,10206
citrate|10207,10214
-|10214,10215
vitamin|10215,10222
D3|10223,10225
)|10225,10226
315|10227,10230
mg|10231,10233
-|10234,10235
<EOL>|10236,10237
200|10237,10240
units|10241,10246
oral|10248,10252
DAILY|10253,10258
<EOL>|10259,10260
25.|10260,10263
cod|10264,10267
liver|10268,10273
oil|10274,10277
1|10278,10279
capsule|10280,10287
oral|10289,10293
BID|10294,10297
<EOL>|10298,10299
26|10299,10301
.|10301,10302
Ipratropium|10303,10314
Bromide|10315,10322
Neb|10323,10326
1|10327,10328
NEB|10329,10332
IH|10333,10335
Q6H|10336,10339
:|10339,10340
PRN|10340,10343
Wheezing|10344,10352
<EOL>|10353,10354
<EOL>|10354,10355
<EOL>|10356,10357
Discharge|10357,10366
Disposition|10367,10378
:|10378,10379
<EOL>|10379,10380
Home|10380,10384
With|10385,10389
Service|10390,10397
<EOL>|10397,10398
<EOL>|10399,10400
Facility|10400,10408
:|10408,10409
<EOL>|10409,10410
_|10410,10411
_|10411,10412
_|10412,10413
<EOL>|10413,10414
<EOL>|10415,10416
Discharge|10416,10425
Diagnosis|10426,10435
:|10435,10436
<EOL>|10436,10437
COPD|10456,10460
exacerbation|10461,10473
<EOL>|10473,10474
<EOL>|10474,10475
SECONDARY|10475,10484
DIAGNOSES|10485,10494
:|10494,10495
<EOL>|10495,10496
CAD|10496,10499
<EOL>|10499,10500
Hypertension|10500,10512
anxiety|10513,10520
<EOL>|10520,10521
<EOL>|10522,10523
Mental|10544,10550
Status|10551,10557
:|10557,10558
Clear|10559,10564
and|10565,10568
coherent|10569,10577
.|10577,10578
<EOL>|10578,10579
Level|10579,10584
of|10585,10587
Consciousness|10588,10601
:|10601,10602
Alert|10603,10608
and|10609,10612
interactive|10613,10624
.|10624,10625
<EOL>|10625,10626
Activity|10626,10634
Status|10635,10641
:|10641,10642
Ambulatory|10643,10653
-|10654,10655
Independent|10656,10667
.|10667,10668
<EOL>|10668,10669
<EOL>|10670,10671
Dear|10695,10699
_|10700,10701
_|10701,10702
_|10702,10703
,|10703,10704
<EOL>|10704,10705
<EOL>|10705,10706
_|10706,10707
_|10707,10708
_|10708,10709
was|10710,10713
a|10714,10715
great|10716,10721
pleasure|10722,10730
taking|10731,10737
care|10738,10742
of|10743,10745
you|10746,10749
at|10750,10752
_|10753,10754
_|10754,10755
_|10755,10756
<EOL>|10757,10758
_|10758,10759
_|10759,10760
_|10760,10761
.|10761,10762
You|10763,10766
came|10767,10771
here|10772,10776
because|10777,10784
you|10785,10788
were|10789,10793
<EOL>|10794,10795
experiencing|10795,10807
worsening|10808,10817
shortness|10818,10827
of|10828,10830
breath|10831,10837
as|10838,10840
well|10841,10845
as|10846,10848
nasal|10849,10854
<EOL>|10855,10856
congestion|10856,10866
and|10867,10870
decreased|10871,10880
hearing|10881,10888
.|10888,10889
Your|10890,10894
symptoms|10895,10903
are|10904,10907
likely|10908,10914
<EOL>|10915,10916
related|10916,10923
to|10924,10926
an|10927,10929
upper|10930,10935
respiratory|10936,10947
tract|10948,10953
infection|10954,10963
and|10964,10967
exacerbation|10968,10980
<EOL>|10981,10982
of|10982,10984
your|10985,10989
COPD|10990,10994
.|10994,10995
We|10996,10998
started|10999,11006
you|11007,11010
on|11011,11013
antibiotics|11014,11025
and|11026,11029
continued|11030,11039
your|11040,11044
<EOL>|11045,11046
prednisone|11046,11056
.|11056,11057
<EOL>|11057,11058
<EOL>|11058,11059
The|11059,11062
dose|11063,11067
of|11068,11070
prednisone|11071,11081
will|11082,11086
be|11087,11089
decreased|11090,11099
by|11100,11102
5|11103,11104
mg|11105,11107
every|11108,11113
two|11114,11117
<EOL>|11118,11119
weeks|11119,11124
;|11124,11125
please|11126,11132
take|11133,11137
your|11138,11142
prednisone|11143,11153
as|11154,11156
follows|11157,11164
:|11164,11165
<EOL>|11165,11166
-|11166,11167
Prednisone|11168,11178
30|11179,11181
mg|11182,11184
for|11185,11188
two|11189,11192
weeks|11193,11198
(|11199,11200
Day|11200,11203
1|11204,11205
=|11205,11206
_|11207,11208
_|11208,11209
_|11209,11210
end|11211,11214
<EOL>|11215,11216
_|11216,11217
_|11217,11218
_|11218,11219
<EOL>|11219,11220
-|11220,11221
Prednisone|11222,11232
25|11233,11235
mg|11236,11238
for|11239,11242
two|11243,11246
weeks|11247,11252
(|11253,11254
Day|11254,11257
1|11258,11259
=|11259,11260
_|11261,11262
_|11262,11263
_|11263,11264
end|11265,11268
<EOL>|11269,11270
_|11270,11271
_|11271,11272
_|11272,11273
<EOL>|11273,11274
-|11274,11275
Prednisone|11276,11286
20|11287,11289
mg|11290,11292
for|11293,11296
two|11297,11300
weeks|11301,11306
(|11307,11308
Day|11308,11311
1|11312,11313
=|11313,11314
_|11315,11316
_|11316,11317
_|11317,11318
end|11319,11322
<EOL>|11323,11324
_|11324,11325
_|11325,11326
_|11326,11327
<EOL>|11327,11328
-|11328,11329
Discuss|11330,11337
with|11338,11342
Dr.|11343,11346
_|11347,11348
_|11348,11349
_|11349,11350
further|11351,11358
taper|11359,11364
at|11365,11367
f|11368,11369
/|11369,11370
u|11370,11371
<EOL>|11372,11373
<EOL>|11373,11374
Please|11374,11380
take|11381,11385
all|11386,11389
your|11390,11394
medications|11395,11406
on|11407,11409
time|11410,11414
and|11415,11418
follow|11419,11425
up|11426,11428
with|11429,11433
your|11434,11438
<EOL>|11439,11440
doctors|11440,11447
as|11448,11450
_|11451,11452
_|11452,11453
_|11453,11454
.|11454,11455
<EOL>|11455,11456
<EOL>|11456,11457
Best|11457,11461
regards|11462,11469
,|11469,11470
<EOL>|11470,11471
Your|11471,11475
_|11476,11477
_|11477,11478
_|11478,11479
team|11480,11484
<EOL>|11484,11485
<EOL>|11486,11487
Followup|11487,11495
Instructions|11496,11508
:|11508,11509
<EOL>|11509,11510
_|11510,11511
_|11511,11512
_|11512,11513
<EOL>|11513,11514

