 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
MEDICINE|158,166
<EOL>|166,167
<EOL>|168,169
Sulfa|181,186
(|187,188
Sulfonamide|188,199
Antibiotics|200,211
)|211,212
/|213,214
Codeine|215,222
/|223,224
Bactrim|225,232
<EOL>|232,233
<EOL>|234,235
Attending|235,244
:|244,245
_|246,247
_|247,248
_|248,249
<EOL>|249,250
<EOL>|251,252
nausea|269,275
,|275,276
vomiting|277,285
,|285,286
cough|287,292
<EOL>|292,293
<EOL>|294,295
Major|295,300
Surgical|301,309
or|310,312
Invasive|313,321
Procedure|322,331
:|331,332
<EOL>|332,333
none|333,337
<EOL>|337,338
<EOL>|338,339
<EOL>|340,341
_|369,370
_|370,371
_|371,372
female|373,379
,|379,380
with|381,385
past|386,390
medical|391,398
history|399,406
significant|407,418
for|419,422
<EOL>|423,424
depression|424,434
,|434,435
hyperlipidemia|436,450
,|450,451
Hysterectomy|452,464
,|464,465
B12|466,469
deficiency|470,480
,|480,481
back|482,486
<EOL>|487,488
pain|488,492
,|492,493
carcinoid|494,503
,|503,504
cervical|505,513
DJD|514,517
,|517,518
depression|519,529
,|529,530
hyperlipidemia|531,545
,|545,546
<EOL>|547,548
osteoarthritis|548,562
,|562,563
and|564,567
history|568,575
of|576,578
Exploratory|579,590
laparotomy|591,601
,|601,602
lysis|603,608
of|609,611
<EOL>|612,613
adhesions|613,622
,|622,623
and|624,627
small|628,633
bowel|634,639
resection|640,649
with|650,654
enteroenterostomy|655,672
for|673,676
<EOL>|677,678
a|678,679
high|680,684
grade|685,690
SBO|691,694
_|695,696
_|696,697
_|697,698
who|699,702
presents|703,711
with|712,716
nausea|717,723
,|723,724
vomiting|725,733
,|733,734
<EOL>|735,736
weakness|736,744
x|745,746
2|747,748
weeks|749,754
.|754,755
She|756,759
has|760,763
been|764,768
uable|769,774
to|775,777
tolerate|778,786
PO|787,789
liquids|790,797
,|797,798
<EOL>|799,800
and|800,803
solids|804,810
.|810,811
Had|812,815
similar|816,823
presentation|824,836
_|837,838
_|838,839
_|839,840
for|841,844
high|845,849
grade|850,855
SBO|856,859
.|859,860
<EOL>|861,862
Denies|862,868
passing|869,876
flatus|877,883
today|884,889
.|889,890
However|891,898
reports|899,906
having|907,913
last|914,918
normal|919,925
<EOL>|926,927
bowel|927,932
movement|933,941
this|942,946
AM|947,949
,|949,950
without|951,958
hematochezia|959,971
,|971,972
melena|973,979
.|979,980
Also|981,985
<EOL>|986,987
reporting|987,996
subjective|997,1007
fever|1008,1013
(|1014,1015
100.0|1015,1020
)|1020,1021
,|1021,1022
non|1023,1026
productive|1027,1037
cough|1038,1043
.|1043,1044
Denies|1045,1051
<EOL>|1052,1053
HA|1053,1055
,|1055,1056
myalgias|1057,1065
.|1065,1066
Takes|1067,1072
NSAIDS|1073,1079
sparingly|1080,1089
.|1089,1090
Denies|1091,1097
alcohol|1098,1105
use.|1106,1110
Denies|1111,1117
<EOL>|1118,1119
sick|1119,1123
contacs|1124,1131
/|1131,1132
travel|1133,1139
or|1140,1142
recent|1143,1149
consumption|1150,1161
of|1162,1164
raw|1165,1168
foods|1169,1174
.|1174,1175
Has|1176,1179
<EOL>|1180,1181
never|1181,1186
had|1187,1190
a|1191,1192
colonoscopy|1193,1204
.|1204,1205
<EOL>|1207,1208
.|1208,1209
<EOL>|1211,1212
In|1212,1214
ED|1215,1217
VS|1218,1220
were|1221,1225
97.8|1226,1230
120|1231,1234
121|1235,1238
/|1238,1239
77|1239,1241
20|1242,1244
98|1245,1247
%|1247,1248
RA|1249,1251
<EOL>|1253,1254
Labs|1254,1258
were|1259,1263
remarkable|1264,1274
for|1275,1278
lactate|1279,1286
2.8|1287,1290
,|1290,1291
alk|1292,1295
phos|1296,1300
293|1301,1304
,|1304,1305
HCT|1306,1309
33|1310,1312
,|1312,1313
WBC|1314,1317
<EOL>|1318,1319
13.9|1319,1323
<EOL>|1325,1326
Imaging|1326,1333
:|1333,1334
CT|1335,1337
abdomen|1338,1345
showed|1346,1352
mult|1353,1357
masses|1358,1364
in|1365,1367
the|1368,1371
liver|1372,1377
,|1377,1378
consistent|1379,1389
<EOL>|1390,1391
with|1391,1395
malignancy|1396,1406
.|1406,1407
CXR|1408,1411
also|1412,1416
showed|1417,1423
multiple|1424,1432
nodules|1433,1440
<EOL>|1442,1443
EKG|1443,1446
:|1446,1447
sinus|1448,1453
,|1453,1454
112|1455,1458
,|1458,1459
NA|1460,1462
,|1462,1463
NI|1464,1466
,|1466,1467
TWI|1468,1471
in|1472,1474
III|1475,1478
,|1478,1479
but|1480,1483
largely|1484,1491
unchanged|1492,1501
from|1502,1506
<EOL>|1507,1508
prior|1508,1513
<EOL>|1515,1516
Interventions|1516,1529
:|1529,1530
zofran|1531,1537
,|1537,1538
tylenol|1539,1546
,|1546,1547
2L|1548,1550
NS|1551,1553
,|1553,1554
GI|1555,1557
was|1558,1561
contacted|1562,1571
and|1572,1575
they|1576,1580
<EOL>|1581,1582
are|1582,1585
planning|1586,1594
on|1595,1597
upper|1598,1603
/|1604,1605
lower|1606,1611
endoscopy|1612,1621
for|1622,1625
cancer|1626,1632
work|1633,1637
-|1637,1638
up|1638,1640
.|1640,1641
<EOL>|1643,1644
.|1644,1645
<EOL>|1647,1648
Vitals|1648,1654
on|1655,1657
transfer|1658,1666
were|1667,1671
99.2|1672,1676
113|1677,1680
119|1681,1684
/|1684,1685
47|1685,1687
26|1688,1690
98|1691,1693
%|1693,1694
<EOL>|1696,1697
<EOL>|1697,1698
<EOL>|1699,1700
<EOL>|1721,1722
#|1728,1729
high|1730,1734
grade|1735,1740
SBO|1741,1744
_|1745,1746
_|1746,1747
_|1747,1748
s|1749,1750
/|1750,1751
p|1751,1752
exploratory|1753,1764
laparotomy|1765,1775
,|1775,1776
lysis|1777,1782
of|1783,1785
<EOL>|1786,1787
adhesions|1787,1796
,|1796,1797
and|1798,1801
small|1802,1807
bowel|1808,1813
resection|1814,1823
with|1824,1828
enteroenterostomy|1829,1846
<EOL>|1847,1848
#|1848,1849
carcinoid|1850,1859
<EOL>|1859,1860
#|1860,1861
hyperlipidemia|1862,1876
<EOL>|1876,1877
#|1877,1878
vitamin|1879,1886
B12|1887,1890
deficiency|1891,1901
<EOL>|1901,1902
#|1902,1903
cervical|1904,1912
DJD|1913,1916
<EOL>|1916,1917
#|1917,1918
osteoarthritis|1919,1933
<EOL>|1934,1935
<EOL>|1935,1936
PSH|1936,1939
:|1939,1940
<EOL>|1941,1942
s|1942,1943
/|1943,1944
p|1944,1945
R|1946,1947
lung|1948,1952
resection|1953,1962
in|1963,1965
_|1966,1967
_|1967,1968
_|1968,1969
at|1970,1972
_|1973,1974
_|1974,1975
_|1975,1976
<EOL>|1976,1977
s|1977,1978
/|1978,1979
p|1979,1980
hysterectomy|1981,1993
in|1994,1996
_|1997,1998
_|1998,1999
_|1999,2000
<EOL>|2000,2001
s|2001,2002
/|2002,2003
p|2003,2004
R|2005,2006
arm|2007,2010
surgery|2011,2018
<EOL>|2018,2019
<EOL>|2019,2020
<EOL>|2021,2022
:|2036,2037
<EOL>|2037,2038
_|2038,2039
_|2039,2040
_|2040,2041
<EOL>|2041,2042
:|2056,2057
<EOL>|2057,2058
non|2058,2061
contributory|2062,2074
<EOL>|2074,2075
<EOL>|2076,2077
On|2092,2094
admission|2095,2104
<EOL>|2104,2105
<EOL>|2105,2106
VS|2106,2108
:|2108,2109
98.9|2110,2114
137|2115,2118
/|2118,2119
95|2119,2121
117|2122,2125
20|2126,2128
100|2129,2132
RA|2133,2135
<EOL>|2137,2138
GENERAL|2138,2145
:|2145,2146
AOx3|2147,2151
,|2151,2152
NAD|2153,2156
<EOL>|2158,2159
HEENT|2159,2164
:|2164,2165
MMM|2166,2169
.|2169,2170
no|2171,2173
JVD|2174,2177
.|2177,2178
neck|2179,2183
supple|2184,2190
.|2190,2191
<EOL>|2193,2194
HEART|2194,2199
:|2199,2200
Regular|2201,2208
tachycardic|2209,2220
,|2220,2221
S1|2222,2224
/|2224,2225
S2|2225,2227
heard|2228,2233
.|2233,2234
no|2235,2237
<EOL>|2238,2239
murmurs|2239,2246
/|2246,2247
gallops|2247,2254
/|2254,2255
rubs|2255,2259
.|2259,2260
<EOL>|2262,2263
LUNGS|2263,2268
:|2268,2269
CTAB|2270,2274
,|2274,2275
non|2276,2279
labored|2280,2287
<EOL>|2289,2290
ABDOMEN|2290,2297
:|2297,2298
soft|2299,2303
,|2303,2304
tender|2305,2311
to|2312,2314
palpation|2315,2324
in|2325,2327
epigastrium|2328,2339
.|2339,2340
<EOL>|2342,2343
EXT|2343,2346
:|2346,2347
wwp|2348,2351
,|2351,2352
no|2353,2355
edema|2356,2361
.|2361,2362
DPs|2363,2366
,|2366,2367
PTs|2368,2371
2|2372,2373
+|2373,2374
.|2374,2375
<EOL>|2377,2378
SKIN|2378,2382
:|2382,2383
dry|2384,2387
,|2387,2388
no|2389,2391
rash|2392,2396
<EOL>|2398,2399
NEURO|2399,2404
/|2404,2405
PSYCH|2405,2410
:|2410,2411
CNs|2412,2415
II|2416,2418
-|2418,2419
XII|2419,2422
intact|2423,2429
.|2429,2430
strength|2431,2439
and|2440,2443
sensation|2444,2453
in|2454,2456
U|2457,2458
/|2458,2459
L|2459,2460
<EOL>|2461,2462
extremities|2462,2473
grossly|2474,2481
intact|2482,2488
.|2488,2489
gait|2490,2494
not|2495,2498
assessed|2499,2507
.|2507,2508
<EOL>|2510,2511
<EOL>|2511,2512
On|2512,2514
Discharge|2515,2524
:|2524,2525
<EOL>|2526,2527
VS|2527,2529
:|2529,2530
98.7|2531,2535
118|2538,2541
/|2541,2542
78|2542,2544
97|2547,2549
20|2551,2553
99RA|2554,2558
<EOL>|2558,2559
GENERAL|2559,2566
:|2566,2567
Patient|2568,2575
is|2576,2578
sitting|2579,2586
in|2587,2589
a|2590,2591
chair|2592,2597
,|2597,2598
appears|2599,2606
comfortable|2607,2618
,|2618,2619
<EOL>|2620,2621
A|2621,2622
+|2622,2623
Ox3|2623,2626
,|2626,2627
cooperative|2628,2639
.|2639,2640
<EOL>|2643,2644
HEENT|2644,2649
:|2649,2650
EOMI|2651,2655
,|2655,2656
PERRLA|2657,2663
,|2663,2664
No|2665,2667
Pallor|2668,2674
or|2675,2677
Jaundice|2678,2686
,|2686,2687
MMM|2688,2691
,|2691,2692
no|2693,2695
JVD|2696,2699
,|2699,2700
neck|2701,2705
<EOL>|2706,2707
supple|2707,2713
.|2713,2714
<EOL>|2716,2717
HEART|2717,2722
:|2722,2723
RRR|2724,2727
,|2727,2728
no|2729,2731
m|2732,2733
/|2733,2734
r|2734,2735
/|2735,2736
g|2736,2737
.|2737,2738
<EOL>|2740,2741
LUNGS|2741,2746
:|2746,2747
CTAB|2748,2752
<EOL>|2754,2755
ABDOMEN|2755,2762
:|2762,2763
obese|2764,2769
,|2769,2770
soft|2771,2775
,|2775,2776
mild|2777,2781
tenderness|2782,2792
on|2793,2795
mid|2796,2799
+|2800,2801
right|2801,2806
epigastrium|2807,2818
<EOL>|2819,2820
w|2820,2821
/|2821,2822
o|2822,2823
peritoneal|2824,2834
signs|2835,2840
,|2840,2841
no|2842,2844
shifting|2845,2853
dullness|2854,2862
,|2862,2863
difficult|2864,2873
to|2874,2876
<EOL>|2877,2878
appreciate|2878,2888
organomegaly|2889,2901
.|2901,2902
<EOL>|2904,2905
EXT|2905,2908
:|2908,2909
wwp|2910,2913
,|2913,2914
no|2915,2917
edema|2918,2923
,|2923,2924
no|2925,2927
signs|2928,2933
of|2934,2936
DVT|2937,2940
<EOL>|2942,2943
SKIN|2943,2947
:|2947,2948
no|2949,2951
rash|2952,2956
,|2956,2957
normal|2958,2964
turgor|2965,2971
<EOL>|2973,2974
NEURO|2974,2979
:|2979,2980
no|2981,2983
gross|2984,2989
deficits|2990,2998
<EOL>|2999,3000
PSYCH|3000,3005
:|3005,3006
appropriate|3007,3018
affect|3019,3025
,|3025,3026
no|3027,3029
preceptual|3030,3040
disturbances|3041,3053
,|3053,3054
no|3055,3057
SI|3058,3060
,|3060,3061
<EOL>|3062,3063
normal|3063,3069
judgment|3070,3078
.|3078,3079
<EOL>|3082,3083
<EOL>|3083,3084
<EOL>|3085,3086
Pertinent|3086,3095
Results|3096,3103
:|3103,3104
<EOL>|3104,3105
_|3105,3106
_|3106,3107
_|3107,3108
03|3109,3111
:|3111,3112
14PM|3112,3116
_|3119,3120
_|3120,3121
_|3121,3122
<EOL>|3122,3123
_|3123,3124
_|3124,3125
_|3125,3126
12|3127,3129
:|3129,3130
50PM|3130,3134
URINE|3135,3140
HOURS|3142,3147
-|3147,3148
RANDOM|3148,3154
<EOL>|3154,3155
_|3155,3156
_|3156,3157
_|3157,3158
12|3159,3161
:|3161,3162
50PM|3162,3166
URINE|3167,3172
UHOLD|3174,3179
-|3179,3180
HOLD|3180,3184
<EOL>|3184,3185
_|3185,3186
_|3186,3187
_|3187,3188
12|3189,3191
:|3191,3192
50PM|3192,3196
URINE|3197,3202
COLOR|3204,3209
-|3209,3210
Straw|3210,3215
APPEAR|3216,3222
-|3222,3223
Clear|3223,3228
SP|3229,3231
_|3232,3233
_|3233,3234
_|3234,3235
<EOL>|3235,3236
_|3236,3237
_|3237,3238
_|3238,3239
12|3240,3242
:|3242,3243
50PM|3243,3247
URINE|3248,3253
BLOOD|3255,3260
-|3260,3261
NEG|3261,3264
NITRITE|3265,3272
-|3272,3273
NEG|3273,3276
PROTEIN|3277,3284
-|3284,3285
NEG|3285,3288
<EOL>|3289,3290
GLUCOSE|3290,3297
-|3297,3298
NEG|3298,3301
KETONE|3302,3308
-|3308,3309
NEG|3309,3312
BILIRUBIN|3313,3322
-|3322,3323
NEG|3323,3326
UROBILNGN|3327,3336
-|3336,3337
NEG|3337,3340
PH|3341,3343
-|3343,3344
5.5|3344,3347
<EOL>|3348,3349
LEUK|3349,3353
-|3353,3354
TR|3354,3356
<EOL>|3356,3357
_|3357,3358
_|3358,3359
_|3359,3360
12|3361,3363
:|3363,3364
50PM|3364,3368
URINE|3369,3374
RBC|3376,3379
-|3379,3380
2|3380,3381
WBC|3382,3385
-|3385,3386
2|3386,3387
BACTERIA|3388,3396
-|3396,3397
NONE|3397,3401
YEAST|3402,3407
-|3407,3408
NONE|3408,3412
<EOL>|3413,3414
EPI|3414,3417
-|3417,3418
2|3418,3419
<EOL>|3419,3420
_|3420,3421
_|3421,3422
_|3422,3423
09|3424,3426
:|3426,3427
54AM|3427,3431
LACTATE|3434,3441
-|3441,3442
2|3442,3443
.|3443,3444
8|3444,3445
*|3445,3446
<EOL>|3446,3447
_|3447,3448
_|3448,3449
_|3449,3450
09|3451,3453
:|3453,3454
45AM|3454,3458
GLUCOSE|3461,3468
-|3468,3469
96|3469,3471
UREA|3472,3476
N|3477,3478
-|3478,3479
7|3479,3480
CREAT|3481,3486
-|3486,3487
0.5|3487,3490
SODIUM|3491,3497
-|3497,3498
138|3498,3501
<EOL>|3502,3503
POTASSIUM|3503,3512
-|3512,3513
3.5|3513,3516
CHLORIDE|3517,3525
-|3525,3526
100|3526,3529
TOTAL|3530,3535
CO2|3536,3539
-|3539,3540
27|3540,3542
ANION|3543,3548
GAP|3549,3552
-|3552,3553
15|3553,3555
<EOL>|3555,3556
_|3556,3557
_|3557,3558
_|3558,3559
09|3560,3562
:|3562,3563
45AM|3563,3567
estGFR|3570,3576
-|3576,3577
Using|3577,3582
this|3583,3587
<EOL>|3587,3588
_|3588,3589
_|3589,3590
_|3590,3591
09|3592,3594
:|3594,3595
45AM|3595,3599
ALT|3602,3605
(|3605,3606
SGPT|3606,3610
)|3610,3611
-|3611,3612
17|3612,3614
AST|3615,3618
(|3618,3619
SGOT|3619,3623
)|3623,3624
-|3624,3625
46|3625,3627
*|3627,3628
ALK|3629,3632
PHOS|3633,3637
-|3637,3638
293|3638,3641
*|3641,3642
TOT|3643,3646
<EOL>|3647,3648
BILI|3648,3652
-|3652,3653
0.5|3653,3656
<EOL>|3656,3657
_|3657,3658
_|3658,3659
_|3659,3660
09|3661,3663
:|3663,3664
45AM|3664,3668
LIPASE|3671,3677
-|3677,3678
14|3678,3680
<EOL>|3680,3681
_|3681,3682
_|3682,3683
_|3683,3684
09|3685,3687
:|3687,3688
45AM|3688,3692
ALBUMIN|3695,3702
-|3702,3703
3|3703,3704
.|3704,3705
0|3705,3706
*|3706,3707
<EOL>|3707,3708
_|3708,3709
_|3709,3710
_|3710,3711
09|3712,3714
:|3714,3715
45AM|3715,3719
_|3722,3723
_|3723,3724
_|3724,3725
AFP|3726,3729
-|3729,3730
1.7|3730,3733
<EOL>|3733,3734
_|3734,3735
_|3735,3736
_|3736,3737
09|3738,3740
:|3740,3741
45AM|3741,3745
WBC|3748,3751
-|3751,3752
13|3752,3754
.|3754,3755
9|3755,3756
*|3756,3757
RBC|3758,3761
-|3761,3762
3|3762,3763
.|3763,3764
94|3764,3766
*|3766,3767
HGB|3768,3771
-|3771,3772
9|3772,3773
.|3773,3774
8|3774,3775
*|3775,3776
HCT|3777,3780
-|3780,3781
33|3781,3783
.|3783,3784
0|3784,3785
*|3785,3786
<EOL>|3787,3788
MCV|3788,3791
-|3791,3792
84|3792,3794
#|3794,3795
MCH|3796,3799
-|3799,3800
25|3800,3802
.|3802,3803
0|3803,3804
*|3804,3805
#|3805,3806
MCHC|3807,3811
-|3811,3812
29|3812,3814
.|3814,3815
9|3815,3816
*|3816,3817
RDW|3818,3821
-|3821,3822
16|3822,3824
.|3824,3825
1|3825,3826
*|3826,3827
<EOL>|3827,3828
_|3828,3829
_|3829,3830
_|3830,3831
09|3832,3834
:|3834,3835
45AM|3835,3839
NEUTS|3842,3847
-|3847,3848
75|3848,3850
.|3850,3851
2|3851,3852
*|3852,3853
LYMPHS|3854,3860
-|3860,3861
17|3861,3863
.|3863,3864
9|3864,3865
*|3865,3866
MONOS|3867,3872
-|3872,3873
5.9|3873,3876
EOS|3877,3880
-|3880,3881
0.7|3881,3884
<EOL>|3885,3886
BASOS|3886,3891
-|3891,3892
0.3|3892,3895
<EOL>|3895,3896
_|3896,3897
_|3897,3898
_|3898,3899
09|3900,3902
:|3902,3903
45AM|3903,3907
PLT|3910,3913
COUNT|3914,3919
-|3919,3920
657|3920,3923
*|3923,3924
#|3924,3925
<EOL>|3925,3926
<EOL>|3926,3927
CT|3927,3929
abdomen|3930,3937
/|3937,3938
pelvis|3938,3944
<EOL>|3944,3945
1.|3945,3947
Innumerable|3948,3959
hepatic|3960,3967
and|3968,3971
pulmonary|3972,3981
metastases|3982,3992
.|3992,3993
No|3995,3997
obvious|3998,4005
<EOL>|4006,4007
primary|4007,4014
<EOL>|4015,4016
malignancy|4016,4026
is|4027,4029
identified|4030,4040
on|4041,4043
this|4044,4048
study|4049,4054
.|4054,4055
<EOL>|4056,4057
<EOL>|4059,4060
2|4060,4061
.|4061,4062
No|4063,4065
evidence|4066,4074
of|4075,4077
small|4078,4083
bowel|4084,4089
obstruction|4090,4101
,|4101,4102
ischemic|4103,4111
colitis|4112,4119
,|4119,4120
<EOL>|4121,4122
fluid|4122,4127
collection|4128,4138
,|4138,4139
<EOL>|4140,4141
or|4141,4143
perforation|4144,4155
.|4155,4156
<EOL>|4157,4158
<EOL>|4158,4159
CXR|4159,4162
:|4162,4163
<EOL>|4164,4165
<EOL>|4166,4167
New|4167,4170
nodular|4171,4178
opacities|4179,4188
within|4189,4195
both|4196,4200
upper|4201,4206
lobes|4207,4212
,|4212,4213
left|4214,4218
greater|4219,4226
than|4227,4231
<EOL>|4232,4233
right|4233,4238
.|4238,4239
<EOL>|4240,4241
are|4250,4253
compatible|4254,4264
with|4265,4269
metastases|4270,4280
,|4280,4281
as|4282,4284
was|4285,4288
noted|4289,4294
in|4295,4297
the|4298,4301
<EOL>|4302,4303
lung|4303,4307
bases|4308,4313
on|4314,4316
the|4317,4320
<EOL>|4321,4322
subsequent|4322,4332
CT|4333,4335
of|4336,4338
the|4339,4342
abdomen|4343,4350
and|4351,4354
pelvis|4355,4361
performed|4362,4371
later|4372,4377
the|4378,4381
same|4382,4386
<EOL>|4387,4388
day|4388,4391
.|4391,4392
<EOL>|4393,4394
<EOL>|4394,4395
<EOL>|4396,4397
_|4420,4421
_|4421,4422
_|4422,4423
Female|4424,4430
with|4431,4435
PMH|4436,4439
significant|4440,4451
for|4452,4455
depression|4456,4466
,|4466,4467
<EOL>|4468,4469
hyperlipidemia|4469,4483
,|4483,4484
Hysterectomy|4485,4497
,|4497,4498
B12|4499,4502
deficiency|4503,4513
,|4513,4514
OA|4515,4517
,|4517,4518
carcinoid|4519,4528
,|4528,4529
<EOL>|4530,4531
cervical|4531,4539
DJD|4540,4543
,|4543,4544
depression|4545,4555
,|4555,4556
SBO|4557,4560
who|4561,4564
presented|4565,4574
with|4575,4579
nausea|4580,4586
,|4586,4587
<EOL>|4588,4589
vomiting|4589,4597
,|4597,4598
weakness|4599,4607
x|4608,4609
2|4610,4611
weeks|4612,4617
and|4618,4621
was|4622,4625
found|4626,4631
to|4632,4634
have|4635,4639
multiple|4640,4648
<EOL>|4649,4650
liver|4650,4655
and|4656,4659
lung|4660,4664
masses|4665,4671
per|4672,4675
CT|4676,4678
consistent|4679,4689
with|4690,4694
metastatic|4695,4705
cancer|4706,4712
<EOL>|4713,4714
of|4714,4716
unknown|4717,4724
primary|4725,4732
.|4732,4733
<EOL>|4734,4735
<EOL>|4735,4736
Patient|4736,4743
was|4744,4747
treated|4748,4755
with|4756,4760
IV|4761,4763
fluids|4764,4770
overnight|4771,4780
for|4781,4784
dehydration|4785,4796
.|4796,4797
<EOL>|4798,4799
She|4799,4802
refused|4803,4810
to|4811,4813
stay|4814,4818
in|4819,4821
the|4822,4825
hospital|4826,4834
for|4835,4838
any|4839,4842
further|4843,4850
work|4851,4855
-|4855,4856
up|4856,4858
or|4859,4861
<EOL>|4862,4863
treatment|4863,4872
and|4873,4876
stated|4877,4883
she|4884,4887
would|4888,4893
rather|4894,4900
go|4901,4903
home|4904,4908
to|4909,4911
to|4912,4914
think|4915,4920
and|4921,4924
<EOL>|4925,4926
see|4926,4929
to|4930,4932
her|4933,4936
affairs|4937,4944
over|4945,4949
the|4950,4953
weekend|4954,4961
and|4962,4965
consider|4966,4974
pursuing|4975,4983
<EOL>|4984,4985
further|4985,4992
work|4993,4997
-|4997,4998
up|4998,5000
as|5001,5003
an|5004,5006
outpatient|5007,5017
.|5017,5018
She|5019,5022
tolerated|5023,5032
oral|5033,5037
fluids|5038,5044
well|5045,5049
<EOL>|5050,5051
w|5051,5052
/|5052,5053
o|5053,5054
vomiting|5055,5063
.|5063,5064
She|5065,5068
remained|5069,5077
hemodynamically|5078,5093
stable|5094,5100
and|5101,5104
afebrile|5105,5113
<EOL>|5114,5115
throughout|5115,5125
her|5126,5129
stay|5130,5134
.|5134,5135
<EOL>|5136,5137
<EOL>|5137,5138
Of|5138,5140
note|5141,5145
patient|5146,5153
has|5154,5157
psychiatric|5158,5169
history|5170,5177
of|5178,5180
depressive|5181,5191
symptoms|5192,5200
<EOL>|5201,5202
and|5202,5205
isolation|5206,5215
tendencies|5216,5226
.|5226,5227
She|5228,5231
denied|5232,5238
any|5239,5242
SI|5243,5245
/|5245,5246
SA|5246,5248
or|5249,5251
any|5252,5255
risk|5256,5260
to|5261,5263
<EOL>|5264,5265
herself|5265,5272
.|5272,5273
She|5275,5278
has|5279,5282
little|5283,5289
social|5290,5296
supports|5297,5305
but|5306,5309
does|5310,5314
have|5315,5319
a|5320,5321
good|5322,5326
<EOL>|5327,5328
relationship|5328,5340
with|5341,5345
her|5346,5349
driver|5350,5356
and|5357,5360
friend|5361,5367
who|5368,5371
came|5372,5376
in|5377,5379
and|5380,5383
was|5384,5387
<EOL>|5388,5389
updated|5389,5396
by|5397,5399
the|5400,5403
medical|5404,5411
team|5412,5416
on|5417,5419
the|5420,5423
morning|5424,5431
of|5432,5434
discharge|5435,5444
and|5445,5448
will|5449,5453
<EOL>|5454,5455
be|5455,5457
taking|5458,5464
her|5465,5468
home|5469,5473
.|5473,5474
She|5475,5478
sees|5479,5483
a|5484,5485
mental|5486,5492
health|5493,5499
provider|5500,5508
at|5509,5511
_|5512,5513
_|5513,5514
_|5514,5515
<EOL>|5516,5517
once|5517,5521
a|5522,5523
month|5524,5529
and|5530,5533
has|5534,5537
a|5538,5539
good|5540,5544
relationship|5545,5557
with|5558,5562
her|5563,5566
primary|5567,5574
care|5575,5579
<EOL>|5580,5581
physician|5581,5590
.|5590,5591
Patient|5592,5599
was|5600,5603
dischaerged|5604,5615
home|5616,5620
at|5621,5623
her|5624,5627
request|5628,5635
.|5635,5636
Home|5637,5641
<EOL>|5642,5643
medications|5643,5654
were|5655,5659
continued|5660,5669
to|5670,5672
which|5673,5678
we|5679,5681
added|5682,5687
some|5688,5692
symptomatic|5693,5704
<EOL>|5705,5706
treatment|5706,5715
for|5716,5719
her|5720,5723
cough|5724,5729
with|5730,5734
benzonatate|5735,5746
and|5747,5750
Guaifenesin|5751,5762
.|5762,5763
We|5764,5766
<EOL>|5767,5768
held|5768,5772
off|5773,5776
on|5777,5779
anti-emetics|5780,5792
for|5793,5796
now|5797,5800
as|5801,5803
she|5804,5807
did|5808,5811
not|5812,5815
want|5816,5820
to|5821,5823
stay|5824,5828
<EOL>|5829,5830
inhouse|5830,5837
to|5838,5840
make|5841,5845
sure|5846,5850
these|5851,5856
would|5857,5862
be|5863,5865
well|5866,5870
tolerated|5871,5880
(|5881,5882
would|5882,5887
need|5888,5892
<EOL>|5893,5894
to|5894,5896
monitor|5897,5904
for|5905,5908
drug|5909,5913
interactions|5914,5926
given|5927,5932
multiple|5933,5941
QTc|5942,5945
prolonging|5946,5956
<EOL>|5957,5958
and|5958,5961
serotonergic|5962,5974
medications|5975,5986
on|5987,5989
her|5990,5993
home|5994,5998
meds|5999,6003
)|6003,6004
.|6004,6005
She|6007,6010
was|6011,6014
<EOL>|6015,6016
instructed|6016,6026
to|6027,6029
maintain|6030,6038
good|6039,6043
hydration|6044,6053
and|6054,6057
try|6058,6061
a|6062,6063
soft|6064,6068
diet|6069,6073
at|6074,6076
<EOL>|6077,6078
home|6078,6082
if|6083,6085
she|6086,6089
can|6090,6093
not|6094,6097
tolerate|6098,6106
regular|6107,6114
diet|6115,6119
.|6119,6120
The|6121,6124
patient|6125,6132
met|6133,6136
with|6137,6141
<EOL>|6142,6143
SW|6143,6145
who|6146,6149
provided|6150,6158
her|6159,6162
with|6163,6167
resources|6168,6177
for|6178,6181
community|6182,6191
councelling|6192,6203
.|6203,6204
<EOL>|6205,6206
Outpatient|6206,6216
appointments|6217,6229
with|6230,6234
oncology|6235,6243
,|6243,6244
GI|6245,6247
and|6248,6251
her|6252,6255
PCP|6256,6259
were|6260,6264
set|6265,6268
<EOL>|6269,6270
up|6270,6272
and|6273,6276
her|6277,6280
PCP|6281,6284
and|6285,6288
mental|6289,6295
health|6296,6302
provider|6303,6311
were|6312,6316
updated|6317,6324
.|6324,6325
Her|6326,6329
PCP|6330,6333
<EOL>|6334,6335
_|6335,6336
_|6336,6337
_|6337,6338
also|6339,6343
_|6344,6345
_|6345,6346
_|6346,6347
with|6348,6352
her|6353,6356
later|6357,6362
today|6363,6368
by|6369,6371
telephone|6372,6381
.|6381,6382
<EOL>|6383,6384
<EOL>|6385,6386
Medications|6386,6397
on|6398,6400
Admission|6401,6410
:|6410,6411
<EOL>|6411,6412
The|6412,6415
Preadmission|6416,6428
Medication|6429,6439
list|6440,6444
is|6445,6447
accurate|6448,6456
and|6457,6460
complete|6461,6469
<EOL>|6469,6470
1.|6470,6472
Albuterol|6473,6482
Inhaler|6483,6490
_|6491,6492
_|6492,6493
_|6493,6494
PUFF|6495,6499
IH|6500,6502
Q6H|6503,6506
:|6506,6507
PRN|6507,6510
wheezing|6511,6519
/|6519,6520
SOB|6520,6523
<EOL>|6524,6525
2.|6525,6527
BuPROPion|6528,6537
150|6538,6541
mg|6542,6544
PO|6545,6547
DAILY|6548,6553
<EOL>|6554,6555
3.|6555,6557
Gabapentin|6558,6568
300|6569,6572
mg|6573,6575
PO|6576,6578
TID|6579,6582
<EOL>|6583,6584
4.|6584,6586
Ibuprofen|6587,6596
800|6597,6600
mg|6601,6603
PO|6604,6606
Q8H|6607,6610
:|6610,6611
PRN|6611,6614
pain|6615,6619
<EOL>|6620,6621
5.|6621,6623
Sertraline|6624,6634
200|6635,6638
mg|6639,6641
PO|6642,6644
DAILY|6645,6650
<EOL>|6651,6652
6.|6652,6654
Simvastatin|6655,6666
40|6667,6669
mg|6670,6672
PO|6673,6675
DAILY|6676,6681
<EOL>|6682,6683
7.|6683,6685
Tizanidine|6686,6696
4|6697,6698
mg|6699,6701
PO|6702,6704
BID|6705,6708
:|6708,6709
PRN|6709,6712
muscle|6713,6719
spasms|6720,6726
/|6726,6727
pain|6727,6731
<EOL>|6732,6733
8.|6733,6735
traZODONE|6736,6745
100|6746,6749
mg|6750,6752
PO|6753,6755
HS|6756,6758
:|6758,6759
PRN|6759,6762
sleep|6763,6768
<EOL>|6769,6770
9.|6770,6772
Triamcinolone|6773,6786
Acetonide|6787,6796
0.1|6797,6800
%|6800,6801
Cream|6802,6807
1|6808,6809
Appl|6810,6814
TP|6815,6817
TID|6818,6821
<EOL>|6822,6823
<EOL>|6823,6824
<EOL>|6825,6826
Discharge|6826,6835
Medications|6836,6847
:|6847,6848
<EOL>|6848,6849
1.|6849,6851
Albuterol|6852,6861
Inhaler|6862,6869
_|6870,6871
_|6871,6872
_|6872,6873
PUFF|6874,6878
IH|6879,6881
Q6H|6882,6885
:|6885,6886
PRN|6886,6889
SOB|6890,6893
<EOL>|6894,6895
2.|6895,6897
BuPROPion|6898,6907
150|6908,6911
mg|6912,6914
PO|6915,6917
DAILY|6918,6923
<EOL>|6924,6925
3.|6925,6927
Gabapentin|6928,6938
300|6939,6942
mg|6943,6945
PO|6946,6948
TID|6949,6952
<EOL>|6953,6954
4.|6954,6956
Sertraline|6957,6967
200|6968,6971
mg|6972,6974
PO|6975,6977
DAILY|6978,6983
<EOL>|6984,6985
5.|6985,6987
Simvastatin|6988,6999
40|7000,7002
mg|7003,7005
PO|7006,7008
DAILY|7009,7014
<EOL>|7015,7016
6.|7016,7018
Tizanidine|7019,7029
4|7030,7031
mg|7032,7034
PO|7035,7037
BID|7038,7041
:|7041,7042
PRN|7042,7045
muscle|7046,7052
spasms|7053,7059
/|7059,7060
pain|7060,7064
<EOL>|7065,7066
7.|7066,7068
traZODONE|7069,7078
100|7079,7082
mg|7083,7085
PO|7086,7088
HS|7089,7091
:|7091,7092
PRN|7092,7095
sleep|7096,7101
<EOL>|7102,7103
8.|7103,7105
Ibuprofen|7106,7115
800|7116,7119
mg|7120,7122
PO|7123,7125
Q8H|7126,7129
:|7129,7130
PRN|7130,7133
pain|7134,7138
<EOL>|7139,7140
9.|7140,7142
Triamcinolone|7143,7156
Acetonide|7157,7166
0.1|7167,7170
%|7170,7171
Cream|7172,7177
1|7178,7179
Appl|7180,7184
TP|7185,7187
TID|7188,7191
<EOL>|7192,7193
10.|7193,7196
Benzonatate|7197,7208
100|7209,7212
mg|7213,7215
PO|7216,7218
TID|7219,7222
:|7222,7223
PRN|7223,7226
cough|7227,7232
<EOL>|7233,7234
RX|7234,7236
*|7237,7238
benzonatate|7238,7249
100|7250,7253
mg|7254,7256
1|7257,7258
capsule|7259,7266
(|7266,7267
s|7267,7268
)|7268,7269
by|7270,7272
mouth|7273,7278
TID|7279,7282
:|7282,7283
PRN|7284,7287
cough|7288,7293
Disp|7294,7298
<EOL>|7299,7300
#|7300,7301
*|7301,7302
60|7302,7304
Capsule|7305,7312
Refills|7313,7320
:|7320,7321
*|7321,7322
0|7322,7323
<EOL>|7323,7324
11.|7324,7327
Guaifenesin|7328,7339
_|7340,7341
_|7341,7342
_|7342,7343
mL|7344,7346
PO|7347,7349
Q6H|7350,7353
:|7353,7354
PRN|7354,7357
cough|7358,7363
<EOL>|7364,7365
RX|7365,7367
*|7368,7369
guaifenesin|7369,7380
100|7381,7384
mg|7385,7387
/|7387,7388
5|7388,7389
mL|7390,7392
_|7393,7394
_|7394,7395
_|7395,7396
ml|7397,7399
by|7400,7402
mouth|7403,7408
Q6H|7409,7412
:|7412,7413
PRN|7413,7416
cough|7417,7422
Disp|7423,7427
<EOL>|7428,7429
#|7429,7430
*|7430,7431
1|7431,7432
Bottle|7433,7439
Refills|7440,7447
:|7447,7448
*|7448,7449
0|7449,7450
<EOL>|7450,7451
<EOL>|7451,7452
<EOL>|7453,7454
Discharge|7454,7463
Disposition|7464,7475
:|7475,7476
<EOL>|7476,7477
Home|7477,7481
<EOL>|7481,7482
<EOL>|7483,7484
Discharge|7484,7493
Diagnosis|7494,7503
:|7503,7504
<EOL>|7504,7505
Liver|7505,7510
and|7511,7514
Lung|7515,7519
Mets|7520,7524
of|7525,7527
unkown|7528,7534
primary|7535,7542
<EOL>|7542,7543
<EOL>|7543,7544
<EOL>|7545,7546
Mental|7567,7573
Status|7574,7580
:|7580,7581
Clear|7582,7587
and|7588,7591
coherent|7592,7600
.|7600,7601
<EOL>|7601,7602
Level|7602,7607
of|7608,7610
Consciousness|7611,7624
:|7624,7625
Alert|7626,7631
and|7632,7635
interactive|7636,7647
.|7647,7648
<EOL>|7648,7649
Activity|7649,7657
Status|7658,7664
:|7664,7665
Ambulatory|7666,7676
-|7677,7678
Independent|7679,7690
.|7690,7691
<EOL>|7691,7692
<EOL>|7692,7693
<EOL>|7694,7695
Dear|7719,7723
_|7724,7725
_|7725,7726
_|7726,7727
,|7727,7728
<EOL>|7729,7730
<EOL>|7730,7731
_|7731,7732
_|7732,7733
_|7733,7734
were|7735,7739
seen|7740,7744
in|7745,7747
the|7748,7751
ED|7752,7754
for|7755,7758
ongoing|7759,7766
cough|7767,7772
,|7772,7773
nausea|7774,7780
and|7781,7784
vomiting|7785,7793
<EOL>|7794,7795
and|7795,7798
had|7799,7802
imaging|7803,7810
studies|7811,7818
which|7819,7824
unfortunately|7825,7838
showed|7839,7845
spots|7846,7851
in|7852,7854
your|7855,7859
<EOL>|7860,7861
liver|7861,7866
and|7867,7870
lungs|7871,7876
which|7877,7882
are|7883,7886
likely|7887,7893
due|7894,7897
to|7898,7900
wide|7901,7905
-|7905,7906
spread|7906,7912
cancer|7913,7919
.|7919,7920
_|7921,7922
_|7922,7923
_|7923,7924
<EOL>|7925,7926
were|7926,7930
admitted|7931,7939
for|7940,7943
further|7944,7951
work|7952,7956
-|7956,7957
up|7957,7959
and|7960,7963
treatment|7964,7973
of|7974,7976
your|7977,7981
<EOL>|7982,7983
symptoms|7983,7991
.|7991,7992
_|7993,7994
_|7994,7995
_|7995,7996
chose|7997,8002
to|8003,8005
not|8006,8009
have|8010,8014
any|8015,8018
more|8019,8023
work|8024,8028
-|8028,8029
up|8029,8031
in|8032,8034
the|8035,8038
hospital|8039,8047
<EOL>|8048,8049
and|8049,8052
wanted|8053,8059
to|8060,8062
be|8063,8065
discharged|8066,8076
home|8077,8081
as|8082,8084
soon|8085,8089
as|8090,8092
possible|8093,8101
.|8101,8102
<EOL>|8103,8104
Please|8104,8110
make|8111,8115
sure|8116,8120
_|8121,8122
_|8122,8123
_|8123,8124
keep|8125,8129
well|8130,8134
hydrated|8135,8143
by|8144,8146
taking|8147,8153
water|8154,8159
sips|8160,8164
<EOL>|8165,8166
throughout|8166,8176
the|8177,8180
day|8181,8184
.|8184,8185
I|8186,8187
also|8188,8192
prescribed|8193,8203
some|8204,8208
symptomatic|8209,8220
treatment|8221,8230
<EOL>|8231,8232
for|8232,8235
your|8236,8240
nausea|8241,8247
and|8248,8251
cough|8252,8257
.|8257,8258
<EOL>|8259,8260
I|8260,8261
updated|8262,8269
your|8270,8274
PCP|8275,8278
and|8279,8282
_|8283,8284
_|8284,8285
_|8285,8286
and|8287,8290
have|8291,8295
set|8296,8299
up|8300,8302
_|8303,8304
_|8304,8305
_|8305,8306
<EOL>|8307,8308
appointments|8308,8320
as|8321,8323
below|8324,8329
.|8329,8330
<EOL>|8332,8333
<EOL>|8334,8335
Followup|8335,8343
Instructions|8344,8356
:|8356,8357
<EOL>|8357,8358
_|8358,8359
_|8359,8360
_|8360,8361
<EOL>|8361,8362

