 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|179,186|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,186|false|false|false|C0009214|codeine|Codeine
Event|Event|SIMPLE_SEGMENT|189,198|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|189,198|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|207,222|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|213,222|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|213,222|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|213,222|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|224,231|false|false|false|||Dyspnea
Finding|Finding|SIMPLE_SEGMENT|224,231|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|224,231|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Event|Event|SIMPLE_SEGMENT|236,242|false|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|236,242|false|false|false|C0025222|Melena|melena
Finding|Classification|SIMPLE_SEGMENT|246,251|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|252,260|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|252,260|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|264,282|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|273,282|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|273,282|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|273,282|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|273,282|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|273,282|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|291,298|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|291,298|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|291,298|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|291,298|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|291,301|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|291,317|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|291,317|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|302,309|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|302,309|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|302,317|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|310,317|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|343,350|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|343,350|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|343,350|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|343,350|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|343,353|false|false|false|C0262926|Medical History|history of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|354,359|false|false|false|C1300072|Tumor stage|stage
Event|Event|SIMPLE_SEGMENT|354,359|false|false|false|||stage
Anatomy|Cell|SIMPLE_SEGMENT|374,378|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|374,378|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|SIMPLE_SEGMENT|379,383|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|379,383|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|379,383|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|379,383|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|379,383|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|379,390|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|384,390|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|384,390|false|false|false|||cancer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|392,395|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|392,395|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|392,395|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|392,395|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|392,395|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|392,395|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|392,395|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|392,395|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|400,403|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|400,403|false|false|false|||CKD
Event|Event|SIMPLE_SEGMENT|408,416|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|422,429|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|422,429|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|422,429|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|SIMPLE_SEGMENT|432,448|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|SIMPLE_SEGMENT|443,448|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|443,448|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|443,448|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|443,448|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|453,459|false|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|453,459|false|false|false|C0025222|Melena|melena
Finding|Body Substance|SIMPLE_SEGMENT|461,468|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|461,468|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|461,468|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|461,472|false|false|false|C0332310|Has patient|Patient has
Event|Event|SIMPLE_SEGMENT|489,495|true|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|489,495|true|false|false|C0025222|Melena|melena
Anatomy|Body Location or Region|SIMPLE_SEGMENT|505,514|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|505,519|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|515,519|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|515,519|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|515,519|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|515,519|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|524,531|true|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|524,531|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|524,531|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Idea or Concept|SIMPLE_SEGMENT|537,546|true|false|false|C1546960|Patient Outcome - Worsening|worsening
Drug|Organic Chemical|SIMPLE_SEGMENT|547,552|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|547,552|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|547,552|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|547,552|true|false|false|C0010200|Coughing|cough
Finding|Idea or Concept|SIMPLE_SEGMENT|567,570|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|567,570|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|576,582|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|583,589|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|583,589|true|false|false|C0015967|Fever|fevers
Anatomy|Body Location or Region|SIMPLE_SEGMENT|593,598|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|593,598|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|593,603|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|593,603|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|599,603|true|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|599,603|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|599,603|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|599,603|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|622,629|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|630,636|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|677,680|false|false|false|||hct
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|677,680|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|677,680|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|hct
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|700,708|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|700,708|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|700,708|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|724,735|false|false|false|||transfusion
Finding|Functional Concept|SIMPLE_SEGMENT|724,735|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|724,735|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Finding|Functional Concept|SIMPLE_SEGMENT|737,746|false|false|false|C3244310|dependent|dependent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|747,753|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|747,753|false|false|false|||anemia
Event|Event|SIMPLE_SEGMENT|778,785|false|false|false|||hypoxic
Finding|Pathologic Function|SIMPLE_SEGMENT|778,785|false|false|false|C0242184|Hypoxia|hypoxic
Event|Event|SIMPLE_SEGMENT|787,790|false|false|false|||ABG
Finding|Gene or Genome|SIMPLE_SEGMENT|787,790|false|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|787,790|false|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Drug|Organic Chemical|SIMPLE_SEGMENT|814,821|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|814,821|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|814,821|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|814,821|false|false|false|C0202115|Lactic acid measurement|lactate
Finding|Body Substance|SIMPLE_SEGMENT|831,838|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|831,838|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|831,838|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|839,848|false|false|false|||responded
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|852,856|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|SIMPLE_SEGMENT|852,856|false|false|false|||nebs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|859,865|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|859,865|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|859,865|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|859,865|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|859,865|false|false|false|C0038435|Stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|871,879|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|871,879|false|false|false|C0038317|Steroids|steroids
Event|Event|SIMPLE_SEGMENT|871,879|false|false|false|||steroids
Drug|Organic Chemical|SIMPLE_SEGMENT|881,889|false|false|false|C0721336|Levaquin|levaquin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|881,889|false|false|false|C0721336|Levaquin|levaquin
Event|Event|SIMPLE_SEGMENT|881,889|false|false|false|||levaquin
Drug|Antibiotic|SIMPLE_SEGMENT|894,905|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|894,905|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|894,905|false|false|false|||ceftriaxone
Event|Event|SIMPLE_SEGMENT|911,922|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|911,922|false|false|false|C2986411|Improvement|improvement
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|931,935|false|false|false|C0312448|short-acting thyroid stimulator|sats
Drug|Hormone|SIMPLE_SEGMENT|931,935|false|false|false|C0312448|short-acting thyroid stimulator|sats
Event|Event|SIMPLE_SEGMENT|931,935|false|false|false|||sats
Event|Event|SIMPLE_SEGMENT|965,972|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|973,978|false|false|false|C3714655|On IV|on IV
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|979,982|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|979,982|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|979,982|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|992,998|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|SIMPLE_SEGMENT|992,998|false|false|false|C0018302|guaiac|guaiac
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|992,1007|false|false|false|C0744492|guaiac positive|guaiac positive
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|999,1007|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|999,1007|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|999,1007|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|999,1007|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1013,1018|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Finding|Finding|SIMPLE_SEGMENT|1013,1024|false|false|false|C5880922|Brown color of stool|brown stool
Event|Event|SIMPLE_SEGMENT|1019,1024|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|1019,1024|false|false|false|C0015733|Feces|stool
Event|Event|SIMPLE_SEGMENT|1026,1029|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1026,1029|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1030,1036|false|false|false|||showed
Finding|Gene or Genome|SIMPLE_SEGMENT|1037,1042|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Tissue|SIMPLE_SEGMENT|1045,1052|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1045,1052|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|1054,1062|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1054,1062|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1054,1062|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1054,1062|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1082,1087|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1082,1087|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1082,1092|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1088,1092|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|1088,1092|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|1093,1101|false|false|false|||collapse
Finding|Finding|SIMPLE_SEGMENT|1093,1101|false|true|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Finding|Pathologic Function|SIMPLE_SEGMENT|1093,1101|false|true|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1093,1101|false|true|false|C0332521|Collapse (morphologic abnormality)|collapse
Event|Event|SIMPLE_SEGMENT|1103,1106|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|1103,1106|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1103,1106|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|1107,1113|false|false|false|||showed
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1115,1120|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1115,1120|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|1115,1120|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1115,1120|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1115,1125|false|false|false|C0039239|Sinus Tachycardia|sinus tach
Event|Event|SIMPLE_SEGMENT|1121,1125|false|false|false|||tach
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1134,1145|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|1134,1145|false|false|false|||depressions
Event|Event|SIMPLE_SEGMENT|1155,1161|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|1165,1173|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1165,1173|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1165,1173|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1165,1173|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1182,1186|false|false|false|||MICU
Event|Event|SIMPLE_SEGMENT|1249,1256|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1257,1264|false|false|false|||feeling
Finding|Finding|SIMPLE_SEGMENT|1257,1271|false|false|false|C0424578|Psychological Well Being|feeling better
Event|Event|SIMPLE_SEGMENT|1265,1271|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|1265,1271|false|false|false|C1550462|Observation Interpretation - better|better
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1282,1291|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|1282,1291|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|1282,1291|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|1282,1291|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|1282,1291|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|1282,1291|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|1293,1303|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1293,1303|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|SIMPLE_SEGMENT|1322,1328|true|false|false|||recall
Event|Event|SIMPLE_SEGMENT|1338,1348|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|1338,1348|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|SIMPLE_SEGMENT|1350,1359|false|false|false|||breathing
Event|Event|SIMPLE_SEGMENT|1360,1367|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1376,1386|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|1376,1386|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|1376,1386|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|1380,1386|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|1380,1386|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1380,1386|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1380,1386|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1380,1386|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|1396,1406|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|1396,1406|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1396,1414|false|false|false|C1384666|hearing impairment|difficulty hearing
Finding|Finding|SIMPLE_SEGMENT|1396,1414|false|false|false|C0018772|Partial Hearing Loss|difficulty hearing
Event|Event|SIMPLE_SEGMENT|1407,1414|false|false|false|||hearing
Finding|Finding|SIMPLE_SEGMENT|1407,1414|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|1407,1414|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Finding|SIMPLE_SEGMENT|1423,1429|true|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|1423,1429|true|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|1423,1429|true|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1423,1434|true|false|false|C0002622|Amnesia|memory loss
Finding|Sign or Symptom|SIMPLE_SEGMENT|1423,1434|true|false|false|C0751295|Memory Loss|memory loss
Event|Event|SIMPLE_SEGMENT|1430,1434|true|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1430,1434|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Body Substance|SIMPLE_SEGMENT|1436,1443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1436,1443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1436,1443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1461,1468|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|1461,1468|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1461,1468|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|SIMPLE_SEGMENT|1510,1517|false|false|false|C0009214|codeine|codeine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1510,1517|false|false|false|C0009214|codeine|codeine
Drug|Clinical Drug|SIMPLE_SEGMENT|1510,1523|false|false|false|C1245651||codeine syrup
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1518,1523|false|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|syrup
Drug|Food|SIMPLE_SEGMENT|1518,1523|false|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|syrup
Event|Event|SIMPLE_SEGMENT|1518,1523|false|false|false|||syrup
Finding|Intellectual Product|SIMPLE_SEGMENT|1528,1532|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1535,1541|false|false|false|||period
Finding|Organism Function|SIMPLE_SEGMENT|1535,1541|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|SIMPLE_SEGMENT|1535,1541|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|SIMPLE_SEGMENT|1546,1557|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|1546,1557|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|1563,1572|true|false|false|||developed
Event|Event|SIMPLE_SEGMENT|1583,1590|true|false|false|||dypsnea
Drug|Organic Chemical|SIMPLE_SEGMENT|1595,1600|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1595,1600|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1595,1600|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1595,1600|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|1620,1626|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1620,1626|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1628,1634|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1628,1634|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1638,1643|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1638,1643|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1638,1648|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1638,1648|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1644,1648|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1644,1648|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1644,1648|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1644,1648|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1654,1660|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1667,1674|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1667,1674|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1667,1674|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1667,1674|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|1679,1685|true|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|1679,1685|true|false|false|C0025222|Melena|melena
Event|Event|SIMPLE_SEGMENT|1698,1704|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1698,1704|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1705,1711|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1705,1711|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1705,1711|false|false|false|C0027497|Nausea|nausea
Finding|Intellectual Product|SIMPLE_SEGMENT|1716,1720|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1716,1729|false|false|false|C5671122||poor appetite
Finding|Intellectual Product|SIMPLE_SEGMENT|1716,1729|false|false|false|C0232462;C4282406|Decrease in appetite;Poor appetite question|poor appetite
Finding|Sign or Symptom|SIMPLE_SEGMENT|1716,1729|false|false|false|C0232462;C4282406|Decrease in appetite;Poor appetite question|poor appetite
Event|Event|SIMPLE_SEGMENT|1721,1729|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|1721,1729|false|false|false|C0003618|Desire for food|appetite
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1746,1755|true|false|false|C0017168|Gastroesophageal reflux disease|heartburn
Event|Event|SIMPLE_SEGMENT|1746,1755|true|false|false|||heartburn
Finding|Sign or Symptom|SIMPLE_SEGMENT|1746,1755|true|false|false|C0018834|Heartburn|heartburn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1759,1768|true|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|SIMPLE_SEGMENT|1759,1768|true|false|false|||dysphagia
Finding|Finding|SIMPLE_SEGMENT|1775,1795|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1780,1787|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1780,1787|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1780,1787|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1780,1787|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1780,1787|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1780,1795|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1788,1795|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1788,1795|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1788,1795|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1797,1802|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|SIMPLE_SEGMENT|1797,1805|false|false|false|C0441772|Stage level 4|Stage IV
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1797,1831|false|false|false|C0278987|Metastatic non-small cell lung cancer|Stage IV nonsmall cell lung cancer
Anatomy|Cell|SIMPLE_SEGMENT|1815,1819|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|1815,1819|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1820,1824|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1820,1824|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1820,1824|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1820,1824|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1820,1831|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1820,1847|false|false|false|C0152013|Adenocarcinoma of lung (disorder)|lung cancer, adenocarcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1825,1831|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1825,1831|false|false|false|||cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1833,1847|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|SIMPLE_SEGMENT|1833,1847|false|false|false|||adenocarcinoma
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1849,1853|false|false|false|C0034802;C1368111;C1739039|EGFR protein, human;Epidermal Growth Factor Receptor;Soluble ErbB-1|EGFR
Drug|Enzyme|SIMPLE_SEGMENT|1849,1853|false|false|false|C0034802;C1368111;C1739039|EGFR protein, human;Epidermal Growth Factor Receptor;Soluble ErbB-1|EGFR
Event|Event|SIMPLE_SEGMENT|1849,1853|false|false|false|||EGFR
Finding|Gene or Genome|SIMPLE_SEGMENT|1849,1853|false|false|false|C0034802;C1150617;C1368111;C1414313;C1739039|EGFR gene;EGFR protein, human;Epidermal Growth Factor Receptor;Soluble ErbB-1;epidermal growth factor receptor activity|EGFR
Finding|Molecular Function|SIMPLE_SEGMENT|1849,1853|false|false|false|C0034802;C1150617;C1368111;C1414313;C1739039|EGFR gene;EGFR protein, human;Epidermal Growth Factor Receptor;Soluble ErbB-1;epidermal growth factor receptor activity|EGFR
Finding|Receptor|SIMPLE_SEGMENT|1849,1853|false|false|false|C0034802;C1150617;C1368111;C1414313;C1739039|EGFR gene;EGFR protein, human;Epidermal Growth Factor Receptor;Soluble ErbB-1;epidermal growth factor receptor activity|EGFR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1849,1853|false|false|false|C3811844|Estimated Glomerular Filtration Rate|EGFR
Event|Event|SIMPLE_SEGMENT|1860,1864|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|1860,1864|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|1860,1864|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1866,1870|false|false|false|C0763464|KRAS protein, human|KRAS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1866,1870|false|false|false|C0763464|KRAS protein, human|KRAS
Event|Event|SIMPLE_SEGMENT|1866,1870|false|false|false|||KRAS
Finding|Gene or Genome|SIMPLE_SEGMENT|1866,1870|false|false|false|C0022457;C1537502;C5441977|Human Oncogene K-Ras;K-ras Oncogene;KRAS gene|KRAS
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1871,1878|false|false|false|C1705285|Mutation Abnormality|mutated
Event|Event|SIMPLE_SEGMENT|1871,1878|false|false|false|||mutated
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1871,1878|false|false|false|C5444829|Gene Variant Positive|mutated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1881,1884|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1881,1884|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1881,1884|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1881,1884|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1881,1884|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1881,1884|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1881,1884|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1881,1884|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|1889,1893|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1889,1893|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1913,1916|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1913,1916|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|1913,1916|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|1913,1916|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|1913,1916|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1913,1916|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1920,1923|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1920,1923|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|1920,1923|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1920,1923|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Intellectual Product|SIMPLE_SEGMENT|1927,1934|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|1927,1934|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1927,1954|false|false|false|C0403447|Chronic Kidney Insufficiency|Chronic renal insufficiency
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1935,1940|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1935,1940|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1935,1954|false|false|false|C0035078;C1565489|Kidney Failure;Renal Insufficiency|renal insufficiency
Event|Event|SIMPLE_SEGMENT|1941,1954|false|false|false|||insufficiency
Finding|Functional Concept|SIMPLE_SEGMENT|1941,1954|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Body Substance|SIMPLE_SEGMENT|1957,1964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1957,1964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1957,1964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1970,1973|false|false|false|||GFR
Finding|Gene or Genome|SIMPLE_SEGMENT|1970,1973|false|false|false|C1424601|RAPGEF5 gene|GFR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1982,1985|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1982,1985|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|1982,1985|false|false|false|||CVA
Finding|Functional Concept|SIMPLE_SEGMENT|1994,1998|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1999,2008|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|SIMPLE_SEGMENT|2017,2024|false|false|false|||infarct
Finding|Pathologic Function|SIMPLE_SEGMENT|2017,2024|false|false|false|C0021308|Infarction|infarct
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2035,2055|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|SIMPLE_SEGMENT|2035,2055|false|false|false|||Hypercholesterolemia
Finding|Finding|SIMPLE_SEGMENT|2035,2055|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2059,2079|false|false|false|C0024437;C0242383|Age related macular degeneration;Macular degeneration|Macular Degeneration
Event|Event|SIMPLE_SEGMENT|2067,2079|false|false|false|||Degeneration
Finding|Functional Concept|SIMPLE_SEGMENT|2067,2079|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degeneration
Finding|Pathologic Function|SIMPLE_SEGMENT|2067,2079|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degeneration
Finding|Functional Concept|SIMPLE_SEGMENT|2085,2091|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2085,2099|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2092,2099|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2092,2099|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2092,2099|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2092,2099|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2105,2111|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2105,2111|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2105,2111|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2105,2111|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2105,2119|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2112,2119|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2112,2119|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2112,2119|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2112,2119|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2125,2131|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|2125,2131|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|SIMPLE_SEGMENT|2132,2136|false|false|false|||died
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2144,2147|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2144,2147|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2144,2147|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2144,2147|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2144,2147|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2144,2147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2144,2147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2144,2147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2151,2154|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2151,2154|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|2151,2154|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|SIMPLE_SEGMENT|2151,2154|false|false|false|||age
Finding|Idea or Concept|SIMPLE_SEGMENT|2164,2170|false|false|false|C1546508|Relationship - Mother|mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2175,2182|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2175,2182|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2175,2182|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|2175,2182|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|2175,2182|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2175,2182|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2185,2191|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2185,2191|false|false|false|||cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2196,2208|false|false|false|C0029463;C0585442|Osteosarcoma;Osteosarcoma of bone|osteosarcoma
Event|Event|SIMPLE_SEGMENT|2196,2208|false|false|false|||osteosarcoma
Finding|Gene or Genome|SIMPLE_SEGMENT|2196,2208|false|false|false|C0694889|RB1 gene|osteosarcoma
Event|Event|SIMPLE_SEGMENT|2215,2223|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2215,2223|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2215,2223|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2215,2223|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2215,2228|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2215,2228|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2224,2228|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2224,2228|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2224,2228|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2230,2237|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|2230,2237|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|2230,2237|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2248,2263|false|false|false|C0008715|Chronically Ill|chronically ill
Finding|Finding|SIMPLE_SEGMENT|2248,2263|false|false|false|C2051413|Patient appears chronically ill|chronically ill
Finding|Sign or Symptom|SIMPLE_SEGMENT|2260,2263|false|false|false|C0231218|Malaise|ill
Event|Event|SIMPLE_SEGMENT|2264,2273|false|false|false|||appearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2284,2287|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2284,2287|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2284,2287|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2284,2287|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2284,2287|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2284,2287|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2284,2287|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2290,2295|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2304,2308|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2310,2316|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2310,2316|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|2310,2316|false|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2310,2316|false|false|false|C2228481|examination of sclera|sclera
Event|Event|SIMPLE_SEGMENT|2317,2326|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2317,2326|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2328,2331|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2328,2331|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2334,2338|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2334,2338|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|2334,2338|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|2340,2346|true|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|2340,2346|true|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|2348,2351|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2348,2351|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|2356,2364|true|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|2384,2397|true|false|false|||submandibular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2399,2402|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2399,2402|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2399,2402|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2399,2402|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2405,2410|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|2422,2432|false|false|false|||percussion
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2422,2432|false|false|false|C0030987;C1880282|Dental Percussion;Percussion|percussion
Finding|Functional Concept|SIMPLE_SEGMENT|2444,2449|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2444,2454|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2450,2454|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2450,2454|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2450,2454|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|2450,2454|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|2450,2454|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|2460,2469|false|false|false|||decreased
Finding|Body Substance|SIMPLE_SEGMENT|2471,2477|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2471,2484|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|2478,2484|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2478,2484|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|2496,2504|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2496,2504|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2512,2517|false|false|false|C0796494|lobe|lobes
Finding|Intellectual Product|SIMPLE_SEGMENT|2528,2532|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|2534,2542|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2534,2542|false|false|false|C0043144|Wheezing|wheezing
Event|Activity|SIMPLE_SEGMENT|2557,2561|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|2557,2561|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|2557,2561|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|2566,2572|true|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2566,2572|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2566,2572|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|2593,2600|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2593,2600|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2602,2606|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2602,2606|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2617,2628|true|false|false|||appreciated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2631,2638|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2631,2638|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|2631,2638|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|2631,2638|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2640,2644|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2640,2644|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2673,2678|true|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2673,2685|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|2679,2685|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2679,2685|true|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|2686,2693|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|2686,2693|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|SIMPLE_SEGMENT|2699,2717|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|SIMPLE_SEGMENT|2707,2717|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2707,2717|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2707,2717|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2721,2729|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2721,2729|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|SIMPLE_SEGMENT|2734,2746|true|false|false|||organomegaly
Finding|Finding|SIMPLE_SEGMENT|2734,2746|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|SIMPLE_SEGMENT|2756,2761|true|false|false|||foley
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2764,2767|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|2764,2767|true|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2764,2767|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|2769,2773|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|2769,2773|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2769,2773|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|2775,2779|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2780,2788|true|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|2793,2799|true|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2793,2799|true|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2793,2799|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2793,2799|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2804,2812|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|2804,2812|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|2814,2822|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2814,2822|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2827,2832|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2827,2832|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2827,2832|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2836,2845|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|2836,2845|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2836,2845|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2836,2845|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2836,2845|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|2847,2854|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|expired
Finding|Organism Function|SIMPLE_SEGMENT|2847,2854|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|expired
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2888,2893|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2888,2893|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2888,2893|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2894,2897|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2903,2906|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2903,2906|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2903,2906|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2913,2916|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2913,2916|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2913,2916|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2913,2916|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2922,2925|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2922,2925|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2933,2936|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2933,2936|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2933,2936|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2933,2936|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2933,2936|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2940,2943|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2940,2943|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2940,2943|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2940,2943|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2940,2943|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2940,2943|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2949,2953|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2949,2953|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2969,2972|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2989,2994|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2989,2994|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2989,2994|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3007,3013|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|3019,3024|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3019,3024|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3019,3024|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3029,3032|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3029,3032|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3029,3032|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3059,3064|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3059,3064|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3059,3064|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3069,3072|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3069,3072|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3069,3072|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3094,3099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3094,3099|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3094,3099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3094,3107|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3094,3107|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3094,3107|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3100,3107|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3100,3107|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3100,3107|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3100,3107|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3100,3107|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3100,3107|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|3145,3146|false|false|false|||5
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3186,3191|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3186,3191|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3186,3191|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3192,3195|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3192,3195|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3192,3195|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3192,3195|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3192,3195|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3192,3195|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3192,3195|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3192,3195|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3199,3202|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3199,3202|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3199,3202|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3199,3202|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3199,3202|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3209,3212|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|3209,3212|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|3209,3212|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|3209,3212|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3209,3212|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3222,3225|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|3222,3225|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|3222,3225|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|3222,3225|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3222,3225|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3231,3238|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|3231,3238|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3266,3271|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3266,3271|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3266,3271|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3272,3277|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3272,3277|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3272,3277|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3272,3277|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3306,3311|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3306,3311|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3306,3311|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3312,3317|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3312,3317|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3312,3317|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3312,3317|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3361,3366|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3361,3366|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3361,3366|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3361,3374|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3367,3374|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3367,3374|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3367,3374|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3367,3374|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3367,3374|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3367,3374|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3367,3374|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3367,3374|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3408,3413|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3408,3413|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3408,3413|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3439,3444|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3439,3444|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3439,3444|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|3449,3452|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|3449,3452|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|3449,3452|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3449,3452|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3457,3461|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3457,3461|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3488,3492|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3488,3492|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3488,3492|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3488,3492|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|3488,3492|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|3488,3492|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Intellectual Product|SIMPLE_SEGMENT|3498,3505|false|false|false|C0282411;C0947611|Comment;Published Comment|Comment
Event|Event|SIMPLE_SEGMENT|3512,3515|false|false|false|||TOP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3528,3533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3528,3533|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3528,3533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3528,3538|false|false|false|C1383165|Blood Type|BLOOD Type
Finding|Classification|SIMPLE_SEGMENT|3528,3538|false|false|false|C0005810;C2911644|Blood Group Systems;Encounter due to blood type|BLOOD Type
Finding|Finding|SIMPLE_SEGMENT|3528,3538|false|false|false|C0005810;C2911644|Blood Group Systems;Encounter due to blood type|BLOOD Type
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3528,3538|false|false|false|C0005844|Blood group typing (procedure)|BLOOD Type
Finding|Gene or Genome|SIMPLE_SEGMENT|3534,3538|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|SIMPLE_SEGMENT|3534,3538|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Drug|Organic Chemical|SIMPLE_SEGMENT|3539,3542|false|false|false|C0052432|artesunate|ART
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3539,3542|false|false|false|C0052432|artesunate|ART
Event|Event|SIMPLE_SEGMENT|3539,3542|false|false|false|||ART
Finding|Gene or Genome|SIMPLE_SEGMENT|3539,3542|false|false|false|C1412286;C3890191|AGRP gene;AGRP wt Allele|ART
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3539,3542|false|false|false|C0872104;C1963724|Antiretroviral therapy;Assisted Reproductive Technologies|ART
Event|Event|SIMPLE_SEGMENT|3543,3546|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|3543,3546|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|3543,3546|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3543,3546|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3551,3555|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3551,3555|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3580,3584|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3580,3584|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3580,3584|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3580,3584|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|3580,3584|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|3580,3584|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3603,3608|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3603,3608|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3603,3608|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3603,3616|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|3609,3616|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3609,3616|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|3609,3616|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3609,3616|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3634,3639|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3634,3639|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3634,3639|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3634,3647|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|3640,3647|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3640,3647|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|3640,3647|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3640,3647|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3665,3670|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3665,3670|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3665,3670|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3665,3678|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|3671,3678|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3671,3678|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|3671,3678|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3671,3678|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3696,3701|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3696,3701|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3696,3701|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3696,3709|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|3702,3709|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3702,3709|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3702,3709|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|SIMPLE_SEGMENT|3727,3732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3727,3732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3727,3732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|3727,3738|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3733,3738|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3733,3738|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|SIMPLE_SEGMENT|3739,3744|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|SIMPLE_SEGMENT|3752,3757|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|3777,3782|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3777,3782|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3777,3782|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3777,3788|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3783,3788|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|3783,3788|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|SIMPLE_SEGMENT|3789,3792|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3789,3792|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3793,3800|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3793,3800|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3793,3800|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|SIMPLE_SEGMENT|3801,3804|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3801,3804|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3805,3812|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3805,3812|false|false|false|C0033684|Proteins|Protein
Event|Event|SIMPLE_SEGMENT|3805,3812|false|false|false|||Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|3805,3812|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3805,3812|false|false|false|C0202202|Protein measurement|Protein
Event|Event|SIMPLE_SEGMENT|3813,3815|false|false|false|||TR
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3817,3824|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3817,3824|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3817,3824|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3817,3824|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3817,3824|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3817,3824|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|3825,3828|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3825,3828|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|3829,3835|false|false|false|C0022634|Ketones|Ketone
Event|Event|SIMPLE_SEGMENT|3836,3839|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3836,3839|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|3848,3851|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|3860,3863|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3877,3880|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3877,3880|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|3893,3898|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3893,3898|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3893,3898|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3893,3902|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|SIMPLE_SEGMENT|3899,3902|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3899,3902|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3899,3902|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|3905,3908|true|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|3908,3909|true|false|false|||-
Drug|Food|SIMPLE_SEGMENT|3925,3930|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|3925,3930|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3925,3930|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3925,3930|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|SIMPLE_SEGMENT|3925,3930|true|false|false|||Yeast
Event|Event|SIMPLE_SEGMENT|3931,3935|true|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3937,3940|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3937,3940|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3937,3940|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|3937,3940|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|3937,3940|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3937,3940|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|SIMPLE_SEGMENT|3937,3940|true|false|false|||Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|3937,3940|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|3937,3940|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3937,3940|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|SIMPLE_SEGMENT|3956,3961|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3956,3961|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3956,3961|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|SIMPLE_SEGMENT|3994,3999|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|3994,3999|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|3994,3999|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|SIMPLE_SEGMENT|4051,4056|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|4051,4056|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|4051,4056|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|SIMPLE_SEGMENT|4070,4074|false|false|false|||PCXR
Finding|Intellectual Product|SIMPLE_SEGMENT|4076,4084|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4085,4096|false|false|false|C2711450|Enlargement (morphologic abnormality)|enlargement
Event|Event|SIMPLE_SEGMENT|4085,4096|false|false|false|||enlargement
Finding|Pathologic Function|SIMPLE_SEGMENT|4085,4096|false|false|false|C0020564|Hypertrophy|enlargement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4085,4096|false|false|false|C1293134|Enlargement procedure|enlargement
Finding|Functional Concept|SIMPLE_SEGMENT|4116,4121|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|SIMPLE_SEGMENT|4122,4129|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4122,4129|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|4131,4139|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|4131,4139|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|4131,4139|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|4131,4139|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4161,4174|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4161,4174|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|4182,4186|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4182,4191|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4187,4191|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4187,4191|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4187,4191|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4187,4191|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|4193,4201|false|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|4203,4212|false|false|false|||extension
Finding|Conceptual Entity|SIMPLE_SEGMENT|4203,4212|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Finding|Functional Concept|SIMPLE_SEGMENT|4203,4212|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4216,4221|false|false|false|C0027651|Neoplasms|tumor
Event|Event|SIMPLE_SEGMENT|4216,4221|false|false|false|||tumor
Finding|Finding|SIMPLE_SEGMENT|4216,4221|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|SIMPLE_SEGMENT|4216,4221|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Event|Event|SIMPLE_SEGMENT|4225,4230|false|false|false|||focal
Finding|Intellectual Product|SIMPLE_SEGMENT|4232,4237|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|4238,4248|false|false|false|||infiltrate
Finding|Functional Concept|SIMPLE_SEGMENT|4238,4248|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|SIMPLE_SEGMENT|4238,4248|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|SIMPLE_SEGMENT|4238,4248|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|SIMPLE_SEGMENT|4253,4264|false|false|false|||combination
Finding|Finding|SIMPLE_SEGMENT|4253,4264|false|false|false|C3811910|combination - answer to question|combination
Event|Event|SIMPLE_SEGMENT|4266,4273|false|false|false|||thereof
Finding|Intellectual Product|SIMPLE_SEGMENT|4279,4284|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4285,4293|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4285,4300|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4285,4300|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Body Substance|SIMPLE_SEGMENT|4306,4313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4306,4313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4306,4313|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|4318,4326|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|4334,4338|false|false|false|||MICU
Event|Event|SIMPLE_SEGMENT|4343,4349|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|4353,4358|false|false|false|||BiPAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4353,4358|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|BiPAP
Drug|Organic Chemical|SIMPLE_SEGMENT|4364,4371|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4364,4371|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|4364,4371|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|4364,4371|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|4399,4408|false|false|false|||contacted
Event|Event|SIMPLE_SEGMENT|4409,4418|false|false|false|||overnight
Event|Event|SIMPLE_SEGMENT|4435,4448|false|false|false|||thoracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4435,4448|false|false|false|C0189477|Thoracentesis|thoracentesis
Event|Event|SIMPLE_SEGMENT|4453,4463|false|false|false|||palliation
Finding|Idea or Concept|SIMPLE_SEGMENT|4469,4480|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|4481,4487|false|false|false|||volume
Finding|Intellectual Product|SIMPLE_SEGMENT|4481,4487|false|false|false|C1705102|Volume (publication)|volume
Finding|Finding|SIMPLE_SEGMENT|4500,4515|false|false|false|C0700049|Encounter due to palliative care|Palliative care
Procedure|Health Care Activity|SIMPLE_SEGMENT|4500,4515|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative care
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4500,4515|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative care
Event|Activity|SIMPLE_SEGMENT|4511,4515|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|4511,4515|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|4511,4515|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|4511,4515|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|4520,4529|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|4538,4546|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|4538,4546|false|false|false|C0679006|Decision|decision
Event|Event|SIMPLE_SEGMENT|4552,4556|false|false|false|||made
Event|Event|SIMPLE_SEGMENT|4560,4565|false|false|false|||focus
Finding|Functional Concept|SIMPLE_SEGMENT|4560,4565|false|false|false|C1285542|Has focus|focus
Drug|Organic Chemical|SIMPLE_SEGMENT|4569,4576|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4569,4576|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|4569,4576|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|4569,4576|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|4593,4600|false|false|false|||visited
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4615,4625|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|4615,4625|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|4615,4625|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|4619,4625|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|4619,4625|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|4619,4625|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|4619,4625|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|4619,4625|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|4635,4647|false|false|false|||transitioned
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4659,4662|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|4659,4662|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|4667,4674|false|false|false|||expired
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4683,4688|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4704,4715|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4704,4715|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|4704,4715|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4704,4715|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|4704,4728|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|4719,4728|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4719,4728|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|4730,4740|false|false|false|C0723110|Robitussin|Robitussin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4730,4740|false|false|false|C0723110|Robitussin|Robitussin
Event|Event|SIMPLE_SEGMENT|4730,4740|false|false|false|||Robitussin
Drug|Organic Chemical|SIMPLE_SEGMENT|4746,4753|false|false|false|C0009214|codeine|codeine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4746,4753|false|false|false|C0009214|codeine|codeine
Event|Event|SIMPLE_SEGMENT|4746,4753|false|false|false|||codeine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4758,4761|false|false|false|C0030481|Tropical Spastic Paraparesis|tsp
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4758,4761|false|false|false|C0076560;C4307536|Thrombospondins;thrombospondin-1, human|tsp
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4758,4761|false|false|false|C0076560;C4307536|Thrombospondins;thrombospondin-1, human|tsp
Event|Event|SIMPLE_SEGMENT|4758,4761|false|false|false|||tsp
Finding|Gene or Genome|SIMPLE_SEGMENT|4758,4761|false|false|false|C1336626;C1710292|THBS1 gene;THBS1 wt Allele|tsp
Drug|Organic Chemical|SIMPLE_SEGMENT|4768,4780|false|false|false|C0286651|atorvastatin|ATORVASTATIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4768,4780|false|false|false|C0286651|atorvastatin|ATORVASTATIN
Event|Event|SIMPLE_SEGMENT|4768,4780|false|false|false|||ATORVASTATIN
Drug|Organic Chemical|SIMPLE_SEGMENT|4782,4789|false|false|false|C0593906|Lipitor|LIPITOR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4782,4789|false|false|false|C0593906|Lipitor|LIPITOR
Event|Event|SIMPLE_SEGMENT|4782,4789|false|false|false|||LIPITOR
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4799,4805|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4812,4818|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|4822,4830|true|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4825,4830|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4825,4830|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|4833,4842|true|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4833,4842|true|false|false|C1170480|One Daily|one daily
Drug|Vitamin|SIMPLE_SEGMENT|4833,4842|true|false|false|C1170480|One Daily|one daily
Event|Activity|SIMPLE_SEGMENT|4848,4860|true|false|false|C1706204|Substitution - change|Substitution
Event|Event|SIMPLE_SEGMENT|4848,4860|true|false|false|||Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|4848,4860|true|false|false|C1555721|Substitution - ActClass|Substitution
Drug|Organic Chemical|SIMPLE_SEGMENT|4863,4874|true|false|false|C0053229|benzonatate|BENZONATATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4863,4874|true|false|false|C0053229|benzonatate|BENZONATATE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4884,4891|true|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|4884,4891|true|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4884,4891|true|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4896,4903|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|4896,4903|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4896,4903|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|SIMPLE_SEGMENT|4907,4915|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4910,4915|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4910,4915|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4922,4927|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|4933,4936|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|4933,4936|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|4939,4949|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|CALCITRIOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4939,4949|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|CALCITRIOL
Drug|Vitamin|SIMPLE_SEGMENT|4939,4949|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|CALCITRIOL
Event|Event|SIMPLE_SEGMENT|4939,4949|false|false|false|||CALCITRIOL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4961,4968|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|4961,4968|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4961,4968|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4973,4980|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|4973,4980|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4973,4980|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|SIMPLE_SEGMENT|4984,4992|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4987,4992|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4987,4992|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|4993,4998|false|false|false|C1720374|Every - dosing instruction fragment|every
Finding|Idea or Concept|SIMPLE_SEGMENT|5008,5011|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5008,5011|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|5014,5024|false|false|false|C0008845|citalopram|CITALOPRAM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5014,5024|false|false|false|C0008845|citalopram|CITALOPRAM
Event|Event|SIMPLE_SEGMENT|5014,5024|false|false|false|||CITALOPRAM
Event|Event|SIMPLE_SEGMENT|5028,5038|false|false|false|||Prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|5048,5056|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5048,5056|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5066,5072|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5079,5085|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5079,5085|false|false|false|||Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5089,5097|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5092,5097|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5092,5097|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|5098,5102|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5098,5108|false|false|false|C3537736|Once A Day|once a day
Event|Event|SIMPLE_SEGMENT|5105,5108|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|5105,5108|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5105,5108|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|5111,5122|false|false|false|C0070166|clopidogrel|CLOPIDOGREL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5111,5122|false|false|false|C0070166|clopidogrel|CLOPIDOGREL
Drug|Organic Chemical|SIMPLE_SEGMENT|5124,5130|false|false|false|C0633084|Plavix|PLAVIX
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5124,5130|false|false|false|C0633084|Plavix|PLAVIX
Event|Event|SIMPLE_SEGMENT|5135,5145|false|false|false|||Prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|5155,5163|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5155,5163|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5175,5181|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5175,5181|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5186,5192|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5196,5204|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5199,5204|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5199,5204|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|5205,5209|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5205,5215|false|false|false|C3537736|Once A Day|once a day
Event|Event|SIMPLE_SEGMENT|5212,5215|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|5212,5215|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5212,5215|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|5218,5228|false|false|false|C0016410|folic acid|FOLIC ACID
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5218,5228|false|false|false|C0016410|folic acid|FOLIC ACID
Drug|Vitamin|SIMPLE_SEGMENT|5218,5228|false|false|false|C0016410|folic acid|FOLIC ACID
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5218,5228|false|false|false|C0523631|Folic acid measurement|FOLIC ACID
Event|Event|SIMPLE_SEGMENT|5224,5228|false|false|false|||ACID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5236,5242|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5249,5255|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5259,5267|true|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5262,5267|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5262,5267|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|5268,5277|true|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5268,5277|true|false|false|C1170480|One Daily|one daily
Drug|Vitamin|SIMPLE_SEGMENT|5268,5277|true|false|false|C1170480|One Daily|one daily
Event|Activity|SIMPLE_SEGMENT|5286,5298|true|false|false|C1706204|Substitution - change|Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|5286,5298|true|false|false|C1555721|Substitution - ActClass|Substitution
Drug|Organic Chemical|SIMPLE_SEGMENT|5301,5310|true|false|false|C0024002|lorazepam|LORAZEPAM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5301,5310|true|false|false|C0024002|lorazepam|LORAZEPAM
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5320,5326|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5333,5339|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5343,5351|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5346,5351|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5346,5351|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|5366,5372|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5377,5383|false|false|false|C4255480||Nausea
Event|Event|SIMPLE_SEGMENT|5377,5383|false|false|false|||Nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5377,5383|false|false|false|C0027497|Nausea|Nausea
Drug|Organic Chemical|SIMPLE_SEGMENT|5386,5396|false|false|false|C0025859|metoprolol|METOPROLOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5386,5396|false|false|false|C0025859|metoprolol|METOPROLOL
Drug|Organic Chemical|SIMPLE_SEGMENT|5386,5405|false|false|false|C0700548|metoprolol tartrate|METOPROLOL TARTRATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5386,5405|false|false|false|C0700548|metoprolol tartrate|METOPROLOL TARTRATE
Drug|Organic Chemical|SIMPLE_SEGMENT|5397,5405|false|false|false|C0039328;C0144544|Tartrates;tartrate|TARTRATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5397,5405|false|false|false|C0039328;C0144544|Tartrates;tartrate|TARTRATE
Drug|Organic Chemical|SIMPLE_SEGMENT|5407,5416|false|false|false|C0700776|Lopressor|LOPRESSOR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5407,5416|false|false|false|C0700776|Lopressor|LOPRESSOR
Event|Event|SIMPLE_SEGMENT|5421,5431|false|false|false|||Prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|5441,5449|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5441,5449|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5462,5468|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5475,5481|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5485,5493|true|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5488,5493|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5488,5493|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5498,5501|true|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5498,5501|true|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5498,5501|true|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|5498,5501|true|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|5498,5501|true|false|false|C1332410|BID gene|BID
Event|Activity|SIMPLE_SEGMENT|5508,5520|true|false|false|C1706204|Substitution - change|Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|5508,5520|true|false|false|C1555721|Substitution - ActClass|Substitution
Drug|Organic Chemical|SIMPLE_SEGMENT|5523,5531|true|false|false|C0040610|tramadol|TRAMADOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5523,5531|true|false|false|C0040610|tramadol|TRAMADOL
Event|Event|SIMPLE_SEGMENT|5523,5531|true|false|false|||TRAMADOL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5523,5531|true|false|false|C1266765|Tramadol measurement (procedure)|TRAMADOL
Event|Event|SIMPLE_SEGMENT|5535,5545|true|false|false|||Prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|5555,5563|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5555,5563|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5573,5579|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5599,5605|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5599,5605|false|false|false|||Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5609,5617|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5612,5617|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5612,5617|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5624,5629|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|5632,5635|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5632,5635|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5639,5645|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5652,5656|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|5652,5656|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5652,5656|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|SIMPLE_SEGMENT|5659,5668|false|false|false|C0040805|trazodone|TRAZODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5659,5668|false|false|false|C0040805|trazodone|TRAZODONE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5677,5683|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5690,5696|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5700,5708|true|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5703,5708|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5703,5708|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|5709,5718|true|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5709,5718|true|false|false|C1170480|One Daily|one daily
Drug|Vitamin|SIMPLE_SEGMENT|5709,5718|true|false|false|C1170480|One Daily|one daily
Event|Event|SIMPLE_SEGMENT|5724,5730|true|false|false|||needed
Event|Activity|SIMPLE_SEGMENT|5736,5748|true|false|false|C1706204|Substitution - change|Substitution
Event|Event|SIMPLE_SEGMENT|5736,5748|true|false|false|||Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|5736,5748|true|false|false|C1555721|Substitution - ActClass|Substitution
Drug|Organic Chemical|SIMPLE_SEGMENT|5751,5758|true|false|false|C0004057|aspirin|ASPIRIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5751,5758|true|false|false|C0004057|aspirin|ASPIRIN
Event|Event|SIMPLE_SEGMENT|5751,5758|true|false|false|||ASPIRIN
Event|Event|SIMPLE_SEGMENT|5762,5772|true|false|false|||Prescribed
Finding|Functional Concept|SIMPLE_SEGMENT|5782,5790|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5782,5790|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5809,5815|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5809,5815|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5809,5825|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5830,5836|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5840,5848|true|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5843,5848|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5843,5848|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|5849,5858|true|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5849,5858|true|false|false|C1170480|One Daily|one daily
Drug|Vitamin|SIMPLE_SEGMENT|5849,5858|true|false|false|C1170480|One Daily|one daily
Event|Activity|SIMPLE_SEGMENT|5866,5878|true|false|false|C1706204|Substitution - change|Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|5866,5878|true|false|false|C1555721|Substitution - ActClass|Substitution
Drug|Organic Chemical|SIMPLE_SEGMENT|5881,5891|true|false|false|C0034665|ranitidine|RANITIDINE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5881,5891|true|false|false|C0034665|ranitidine|RANITIDINE
Drug|Organic Chemical|SIMPLE_SEGMENT|5881,5895|true|false|false|C0700466|ranitidine hydrochloride|RANITIDINE HCL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5881,5895|true|false|false|C0700466|ranitidine hydrochloride|RANITIDINE HCL
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5892,5895|true|false|false|C0023443|Hairy Cell Leukemia|HCL
Drug|Immunologic Factor|SIMPLE_SEGMENT|5892,5895|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5892,5895|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5892,5895|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Event|Event|SIMPLE_SEGMENT|5892,5895|true|false|false|||HCL
Drug|Organic Chemical|SIMPLE_SEGMENT|5897,5909|true|false|false|C4765118|Acid Control|ACID CONTROL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5897,5909|true|false|false|C4765118|Acid Control|ACID CONTROL
Drug|Organic Chemical|SIMPLE_SEGMENT|5902,5909|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|CONTROL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5902,5909|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|CONTROL
Drug|Substance|SIMPLE_SEGMENT|5902,5909|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|CONTROL
Event|Event|SIMPLE_SEGMENT|5902,5909|false|false|false|||CONTROL
Finding|Conceptual Entity|SIMPLE_SEGMENT|5902,5909|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|CONTROL
Finding|Functional Concept|SIMPLE_SEGMENT|5902,5909|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|CONTROL
Finding|Idea or Concept|SIMPLE_SEGMENT|5902,5909|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|CONTROL
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5920,5926|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5933,5939|false|false|false|C0039225|Tablet Dosage Form|Tablet
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5949,5954|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5949,5954|true|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|5955,5964|true|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5955,5964|true|false|false|C1170480|One Daily|one daily
Drug|Vitamin|SIMPLE_SEGMENT|5955,5964|true|false|false|C1170480|One Daily|one daily
Event|Activity|SIMPLE_SEGMENT|5970,5982|true|false|false|C1706204|Substitution - change|Substitution
Event|Event|SIMPLE_SEGMENT|5970,5982|true|false|false|||Substitution
Finding|Idea or Concept|SIMPLE_SEGMENT|5970,5982|true|false|false|C1555721|Substitution - ActClass|Substitution
Event|Event|SIMPLE_SEGMENT|5987,5996|true|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5987,5996|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5987,5996|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5987,5996|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5987,5996|true|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5987,6008|true|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5997,6008|true|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5997,6008|true|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5997,6008|true|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5997,6008|true|false|false|C4284232|Medications|Medications
Event|Event|SIMPLE_SEGMENT|6010,6011|false|false|false|||N
Event|Event|SIMPLE_SEGMENT|6016,6025|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6016,6025|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6016,6025|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6016,6025|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6016,6025|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6016,6037|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6016,6037|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6026,6037|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|6026,6037|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6026,6037|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|6039,6046|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Finding|Organism Function|SIMPLE_SEGMENT|6039,6046|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Event|Event|SIMPLE_SEGMENT|6049,6058|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6049,6058|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6049,6058|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6049,6058|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6049,6058|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6049,6068|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6059,6068|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|6059,6068|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6059,6068|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6059,6068|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6059,6068|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6077,6099|false|false|false|C0149925|Small cell carcinoma of lung|small cell lung cancer
Anatomy|Cell|SIMPLE_SEGMENT|6083,6087|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|6083,6087|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6088,6092|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6088,6092|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6088,6092|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|6088,6092|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6088,6099|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6093,6099|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|6093,6099|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|6103,6109|false|false|false|||Melena
Finding|Pathologic Function|SIMPLE_SEGMENT|6103,6109|false|false|false|C0025222|Melena|Melena
Event|Event|SIMPLE_SEGMENT|6112,6121|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6112,6121|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6112,6121|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6112,6121|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6112,6121|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6122,6131|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6122,6131|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|6122,6131|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6122,6131|false|false|false|C1705253|Logical Condition|Condition
Finding|Idea or Concept|SIMPLE_SEGMENT|6133,6140|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Finding|Organism Function|SIMPLE_SEGMENT|6133,6140|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Event|Event|SIMPLE_SEGMENT|6143,6152|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6143,6152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6143,6152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6143,6152|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6143,6152|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6143,6165|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6143,6165|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|6143,6165|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6153,6165|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6153,6165|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6153,6165|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|6167,6168|false|false|false|||N
Procedure|Health Care Activity|SIMPLE_SEGMENT|6173,6181|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6182,6194|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6182,6194|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6182,6194|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

