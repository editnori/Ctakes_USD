 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
Codeine|179,186
<EOL>|186,187
<EOL>|188,189
Attending|189,198
:|198,199
_|200,201
_|201,202
_|202,203
.|203,204
<EOL>|204,205
<EOL>|206,207
Chief|207,212
Complaint|213,222
:|222,223
<EOL>|223,224
chest|224,229
pressure|230,238
<EOL>|238,239
<EOL>|240,241
Major|241,246
Surgical|247,255
or|256,258
Invasive|259,267
Procedure|268,277
:|277,278
<EOL>|278,279
Cardiac|279,286
cathetherization|287,303
<EOL>|303,304
<EOL>|304,305
<EOL>|306,307
History|307,314
of|315,317
Present|318,325
Illness|326,333
:|333,334
<EOL>|334,335
_|335,336
_|336,337
_|337,338
is|339,341
a|342,343
_|344,345
_|345,346
_|346,347
yo|348,350
female|351,357
with|358,362
a|363,364
past|365,369
medical|370,377
history|378,385
of|386,388
<EOL>|389,390
CAD|390,393
with|394,398
a|399,400
1|401,402
vessel|403,409
CABG|410,414
(|415,416
SVG|416,419
to|420,422
LAD|423,426
)|426,427
in|428,430
_|431,432
_|432,433
_|433,434
who|435,438
presents|439,447
with|448,452
<EOL>|453,454
chest|454,459
pressure|460,468
.|468,469
She|471,474
woke|475,479
up|480,482
at|483,485
8|486,487
am|488,490
with|491,495
substernal|496,506
chest|507,512
<EOL>|513,514
pressure|514,522
.|522,523
It|525,527
was|528,531
severe|532,538
initially|539,548
.|548,549
She|551,554
took|555,559
SL|560,562
NTG|563,566
x3|567,569
with|570,574
<EOL>|575,576
relief|576,582
of|583,585
CP|586,588
for|589,592
a|593,594
short|595,600
period|601,607
of|608,610
time|611,615
.|615,616
The|618,621
CP|622,624
radiated|625,633
to|634,636
her|637,640
<EOL>|641,642
right|642,647
side|648,652
and|653,656
eventually|657,667
down|668,672
both|673,677
arms|678,682
.|682,683
She|685,688
reports|689,696
<EOL>|697,698
diaphoresis|698,709
,|709,710
but|711,714
denied|715,721
associated|722,732
nausea|733,739
,|739,740
vomiting|741,749
,|749,750
<EOL>|751,752
lightheadedness|752,767
or|768,770
dizziness|771,780
.|780,781
She|783,786
reports|787,794
that|795,799
she|800,803
has|804,807
felt|808,812
<EOL>|813,814
mildly|814,820
SOB|821,824
since|825,830
her|831,834
recent|835,841
pneumonia|842,851
(|852,853
first|853,858
diagnosed|859,868
appox|869,874
_|875,876
_|876,877
_|877,878
<EOL>|879,880
weeks|880,885
ago|886,889
)|889,890
.|890,891
She|893,896
denied|897,903
worsening|904,913
dyspnea|914,921
.|921,922
Her|924,927
cough|928,933
has|934,937
<EOL>|938,939
improved|939,947
substantially|948,961
and|962,965
is|966,968
very|969,973
minimal|974,981
at|982,984
this|985,989
time|990,994
.|994,995
She|997,1000
<EOL>|1001,1002
went|1002,1006
to|1007,1009
her|1010,1013
PCP|1014,1017
's|1017,1019
office|1020,1026
and|1027,1030
was|1031,1034
found|1035,1040
to|1041,1043
have|1044,1048
a|1049,1050
new|1051,1054
LBBB|1055,1059
and|1060,1063
<EOL>|1064,1065
anterior|1065,1073
ST|1074,1076
elevations|1077,1087
.|1087,1088
She|1090,1093
was|1094,1097
transferred|1098,1109
to|1110,1112
the|1113,1116
ED|1117,1119
.|1119,1120
She|1121,1124
<EOL>|1125,1126
received|1126,1134
Plavix|1135,1141
300mg|1142,1147
,|1147,1148
Aspirin|1149,1156
,|1156,1157
boluses|1158,1165
of|1166,1168
heparin|1169,1176
and|1177,1180
<EOL>|1181,1182
integrillin|1182,1193
.|1193,1194
Code|1195,1199
STEMI|1200,1205
was|1206,1209
called|1210,1216
and|1217,1220
went|1221,1225
to|1226,1228
the|1229,1232
cath|1233,1237
lab|1238,1241
.|1241,1242
<EOL>|1244,1245
Cath|1245,1249
showed|1250,1256
occluded|1257,1265
SVG|1266,1269
,|1269,1270
Native|1271,1277
3vd|1278,1281
,|1281,1282
occluded|1283,1291
proximal|1292,1300
LAD|1301,1304
.|1304,1305
<EOL>|1306,1307
Wiring|1307,1313
the|1314,1317
LAD|1318,1321
was|1322,1325
difficult|1326,1335
and|1336,1339
there|1340,1345
was|1346,1349
concern|1350,1357
about|1358,1363
a|1364,1365
<EOL>|1366,1367
possible|1367,1375
dissection|1376,1386
.|1386,1387
One|1388,1391
BMS|1392,1395
was|1396,1399
placed|1400,1406
in|1407,1409
the|1410,1413
proximal|1414,1422
LAD|1423,1426
.|1426,1427
<EOL>|1428,1429
Distal|1429,1435
LAD|1436,1439
is|1440,1442
diminutive|1443,1453
past|1454,1458
_|1459,1460
_|1460,1461
_|1461,1462
septal|1463,1469
and|1470,1473
diag|1474,1478
branches|1479,1487
.|1487,1488
<EOL>|1491,1492
She|1492,1495
has|1496,1499
been|1500,1504
hemodynamically|1505,1520
stable|1521,1527
with|1528,1532
HR|1533,1535
60|1536,1538
-|1538,1539
70s|1539,1542
and|1543,1546
SBP|1547,1550
<EOL>|1551,1552
120|1552,1555
-|1555,1556
130s|1556,1560
.|1560,1561
On|1563,1565
the|1566,1569
floor|1570,1575
,|1575,1576
she|1577,1580
is|1581,1583
currently|1584,1593
chest|1594,1599
pain|1600,1604
free|1605,1609
and|1610,1613
<EOL>|1614,1615
feels|1615,1620
well|1621,1625
.|1625,1626
<EOL>|1626,1627
.|1627,1628
<EOL>|1631,1632
.|1632,1633
<EOL>|1635,1636
On|1636,1638
review|1639,1645
of|1646,1648
systems|1649,1656
,|1656,1657
she|1658,1661
denies|1662,1668
any|1669,1672
prior|1673,1678
history|1679,1686
of|1687,1689
deep|1690,1694
<EOL>|1695,1696
venous|1696,1702
thrombosis|1703,1713
,|1713,1714
pulmonary|1715,1724
embolism|1725,1733
,|1733,1734
bleeding|1735,1743
at|1744,1746
the|1747,1750
time|1751,1755
of|1756,1758
<EOL>|1759,1760
surgery|1760,1767
,|1767,1768
myalgias|1769,1777
,|1777,1778
joint|1779,1784
pains|1785,1790
,|1790,1791
cough|1792,1797
,|1797,1798
hemoptysis|1799,1809
,|1809,1810
black|1811,1816
stools|1817,1823
<EOL>|1824,1825
or|1825,1827
red|1828,1831
stools|1832,1838
.|1838,1839
She|1840,1843
denies|1844,1850
recent|1851,1857
fevers|1858,1864
,|1864,1865
chills|1866,1872
or|1873,1875
rigors|1876,1882
.|1882,1883
All|1884,1887
<EOL>|1888,1889
of|1889,1891
the|1892,1895
other|1896,1901
review|1902,1908
of|1909,1911
systems|1912,1919
were|1920,1924
negative|1925,1933
.|1933,1934
<EOL>|1936,1937
.|1937,1938
<EOL>|1940,1941
Cardiac|1941,1948
review|1949,1955
of|1956,1958
systems|1959,1966
is|1967,1969
notable|1970,1977
for|1978,1981
absence|1982,1989
of|1990,1992
chest|1993,1998
pain|1999,2003
,|2003,2004
<EOL>|2005,2006
dyspnea|2006,2013
on|2014,2016
exertion|2017,2025
,|2025,2026
paroxysmal|2027,2037
nocturnal|2038,2047
dyspnea|2048,2055
,|2055,2056
orthopnea|2057,2066
,|2066,2067
<EOL>|2068,2069
ankle|2069,2074
edema|2075,2080
,|2080,2081
palpitations|2082,2094
,|2094,2095
syncope|2096,2103
or|2104,2106
presyncope|2107,2117
.|2117,2118
<EOL>|2120,2121
<EOL>|2121,2122
<EOL>|2123,2124
Past|2124,2128
Medical|2129,2136
History|2137,2144
:|2144,2145
<EOL>|2145,2146
1.|2146,2148
CARDIAC|2149,2156
RISK|2157,2161
FACTORS|2162,2169
:|2169,2170
-|2171,2172
Diabetes|2173,2181
,|2181,2182
+|2183,2184
Dyslipidemia|2185,2197
,|2197,2198
+|2199,2200
<EOL>|2201,2202
Hypertension|2202,2214
<EOL>|2216,2217
2.|2217,2219
CARDIAC|2220,2227
HISTORY|2228,2235
:|2235,2236
<EOL>|2238,2239
-|2239,2240
CABG|2240,2244
:|2244,2245
Pt|2246,2248
with|2249,2253
MI|2254,2256
in|2257,2259
_|2260,2261
_|2261,2262
_|2262,2263
and|2264,2267
subsequent|2268,2278
1|2279,2280
vessel|2281,2287
CABG|2288,2292
SVG|2293,2296
-|2297,2298
>|2298,2299
LAD|2299,2302
<EOL>|2302,2303
-|2303,2304
PERCUTANEOUS|2304,2316
CORONARY|2317,2325
INTERVENTIONS|2326,2339
:|2339,2340
none|2342,2346
<EOL>|2346,2347
-|2347,2348
PACING|2348,2354
/|2354,2355
ICD|2355,2358
:|2358,2359
none|2361,2365
<EOL>|2365,2366
3.|2366,2368
OTHER|2369,2374
PAST|2375,2379
MEDICAL|2380,2387
HISTORY|2388,2395
:|2395,2396
<EOL>|2398,2399
#|2399,2400
CVA|2401,2404
-|2405,2406
small|2407,2412
left|2413,2417
posterior|2418,2427
frontal|2428,2435
infarct|2436,2443
in|2444,2446
_|2447,2448
_|2448,2449
_|2449,2450
<EOL>|2451,2452
for|2452,2455
which|2456,2461
she|2462,2465
is|2466,2468
on|2469,2471
_|2472,2473
_|2473,2474
_|2474,2475
tab|2476,2479
of|2480,2482
plavix|2483,2489
daily|2490,2495
<EOL>|2495,2496
#|2496,2497
hypercholesterolemia|2498,2518
.|2518,2519
<EOL>|2521,2522
#|2522,2523
small|2524,2529
PFO|2530,2533
.|2533,2534
<EOL>|2534,2535
#|2535,2536
Macular|2537,2544
Degereration|2545,2557
<EOL>|2557,2558
<EOL>|2559,2560
Social|2560,2566
History|2567,2574
:|2574,2575
<EOL>|2575,2576
_|2576,2577
_|2577,2578
_|2578,2579
<EOL>|2579,2580
Family|2580,2586
History|2587,2594
:|2594,2595
<EOL>|2595,2596
Her|2596,2599
father|2600,2606
died|2607,2611
due|2612,2615
to|2616,2618
CAD|2619,2622
at|2623,2625
age|2626,2629
_|2630,2631
_|2631,2632
_|2632,2633
.|2633,2634
Her|2636,2639
mother|2640,2646
had|2647,2650
<EOL>|2650,2651
stomach|2651,2658
cancer|2659,2665
and|2666,2669
bone|2670,2674
cancer|2675,2681
.|2681,2682
<EOL>|2682,2683
<EOL>|2684,2685
Physical|2685,2693
Exam|2694,2698
:|2698,2699
<EOL>|2699,2700
GENERAL|2700,2707
:|2707,2708
WDWN|2709,2713
in|2714,2716
NAD|2717,2720
.|2720,2721
Oriented|2722,2730
x3|2731,2733
.|2733,2734
Mood|2735,2739
,|2739,2740
affect|2741,2747
appropriate|2748,2759
.|2759,2760
<EOL>|2762,2763
HEENT|2763,2768
:|2768,2769
NCAT|2770,2774
.|2774,2775
Sclera|2776,2782
anicteric|2783,2792
.|2792,2793
PERRL|2794,2799
,|2799,2800
EOMI|2801,2805
.|2805,2806
Conjunctiva|2807,2818
were|2819,2823
<EOL>|2824,2825
pink|2825,2829
,|2829,2830
no|2831,2833
pallor|2834,2840
or|2841,2843
cyanosis|2844,2852
of|2853,2855
the|2856,2859
oral|2860,2864
mucosa|2865,2871
.|2871,2872
No|2873,2875
xanthalesma|2876,2887
.|2887,2888
<EOL>|2890,2891
<EOL>|2891,2892
NECK|2892,2896
:|2896,2897
Supple|2898,2904
with|2905,2909
JVP|2910,2913
of|2914,2916
8|2917,2918
cm|2919,2921
.|2921,2922
<EOL>|2924,2925
CARDIAC|2925,2932
:|2932,2933
PMI|2934,2937
located|2938,2945
in|2946,2948
_|2949,2950
_|2950,2951
_|2951,2952
intercostal|2953,2964
space|2965,2970
,|2970,2971
midclavicular|2972,2985
<EOL>|2986,2987
line|2987,2991
.|2991,2992
RR|2993,2995
,|2995,2996
normal|2997,3003
S1|3004,3006
,|3006,3007
S2|3008,3010
.|3010,3011
No|3012,3014
m|3015,3016
/|3016,3017
r|3017,3018
/|3018,3019
g|3019,3020
.|3020,3021
No|3022,3024
thrills|3025,3032
,|3032,3033
lifts|3034,3039
.|3039,3040
No|3041,3043
S3|3044,3046
or|3047,3049
<EOL>|3050,3051
S4|3051,3053
.|3053,3054
<EOL>|3056,3057
LUNGS|3057,3062
:|3062,3063
No|3064,3066
chest|3067,3072
wall|3073,3077
deformities|3078,3089
,|3089,3090
scoliosis|3091,3100
or|3101,3103
kyphosis|3104,3112
.|3112,3113
Resp|3114,3118
<EOL>|3119,3120
were|3120,3124
unlabored|3125,3134
,|3134,3135
no|3136,3138
accessory|3139,3148
muscle|3149,3155
use|3156,3159
.|3159,3160
CTA|3161,3164
anteriorly|3165,3175
,|3175,3176
no|3177,3179
<EOL>|3180,3181
crackles|3181,3189
,|3189,3190
wheezes|3191,3198
or|3199,3201
rhonchi|3202,3209
.|3209,3210
<EOL>|3212,3213
ABDOMEN|3213,3220
:|3220,3221
Soft|3222,3226
,|3226,3227
NTND|3228,3232
.|3232,3233
No|3234,3236
HSM|3237,3240
or|3241,3243
tenderness|3244,3254
.|3254,3255
Abd|3256,3259
aorta|3260,3265
not|3266,3269
<EOL>|3270,3271
enlarged|3271,3279
by|3280,3282
palpation|3283,3292
.|3292,3293
No|3294,3296
abdominial|3297,3307
bruits|3308,3314
.|3314,3315
<EOL>|3317,3318
EXTREMITIES|3318,3329
:|3329,3330
No|3331,3333
c|3334,3335
/|3335,3336
c|3336,3337
/|3337,3338
e|3338,3339
.|3339,3340
Femoral|3341,3348
sheath|3349,3355
in|3356,3358
place|3359,3364
in|3365,3367
right|3368,3373
groin|3374,3379
.|3379,3380
<EOL>|3382,3383
SKIN|3383,3387
:|3387,3388
No|3389,3391
stasis|3392,3398
dermatitis|3399,3409
,|3409,3410
ulcers|3411,3417
,|3417,3418
scars|3419,3424
,|3424,3425
or|3426,3428
xanthomas|3429,3438
.|3438,3439
<EOL>|3441,3442
PULSES|3442,3448
:|3448,3449
<EOL>|3451,3452
Right|3452,3457
:|3457,3458
Carotid|3459,3466
2|3467,3468
+|3468,3469
DP|3470,3472
2|3473,3474
+|3474,3475
_|3476,3477
_|3477,3478
_|3478,3479
2|3480,3481
+|3481,3482
<EOL>|3484,3485
Left|3485,3489
:|3489,3490
Carotid|3491,3498
2|3499,3500
+|3500,3501
DP|3502,3504
2|3505,3506
+|3506,3507
_|3508,3509
_|3509,3510
_|3510,3511
2|3512,3513
+|3513,3514
<EOL>|3516,3517
<EOL>|3518,3519
Pertinent|3519,3528
Results|3529,3536
:|3536,3537
<EOL>|3537,3538
EKG|3538,3541
:|3541,3542
new|3544,3547
LBBB|3548,3552
with|3553,3557
STE|3558,3561
in|3562,3564
V1|3565,3567
-|3568,3569
V3|3569,3571
&|3572,3573
V5|3574,3576
that|3577,3581
in|3582,3584
some|3585,3589
leads|3590,3595
are|3596,3599
<EOL>|3600,3601
>|3601,3602
5mm|3602,3605
.|3605,3606
<EOL>|3607,3608
TELEMETRY|3608,3617
:|3617,3618
NSR|3619,3622
75|3623,3625
,|3625,3626
few|3627,3630
NSVTs|3631,3636
.|3636,3637
<EOL>|3640,3641
2D|3641,3643
-|3643,3644
ECHOCARDIOGRAM|3644,3658
:|3658,3659
pending|3661,3668
<EOL>|3668,3669
ETT|3669,3672
:|3672,3673
n|3675,3676
/|3676,3677
a|3677,3678
<EOL>|3678,3679
.|3679,3680
<EOL>|3682,3683
CARDIAC|3683,3690
CATH|3691,3695
:|3695,3696
<EOL>|3698,3699
LMCA|3699,3703
:|3703,3704
40|3705,3707
%|3707,3708
distal|3709,3715
<EOL>|3715,3716
LAD|3716,3719
:|3719,3720
Occluded|3721,3729
difficult|3730,3739
to|3740,3742
cross|3743,3748
;|3748,3749
was|3750,3753
crossed|3754,3761
and|3762,3765
stented|3766,3773
in|3774,3776
<EOL>|3777,3778
proximal|3778,3786
LAD|3787,3790
.|3790,3791
Distal|3793,3799
LAD|3800,3803
diffuse|3804,3811
diseased|3812,3820
.|3820,3821
<EOL>|3823,3824
LCX|3824,3827
:|3827,3828
occluded|3829,3837
OM2|3838,3841
,|3841,3842
50|3843,3845
%|3845,3846
LCX|3847,3850
<EOL>|3850,3851
RCA|3851,3854
:|3854,3855
Occluded|3856,3864
<EOL>|3864,3865
<EOL>|3866,3867
Brief|3867,3872
Hospital|3873,3881
Course|3882,3888
:|3888,3889
<EOL>|3889,3890
_|3890,3891
_|3891,3892
_|3892,3893
is|3894,3896
a|3897,3898
_|3899,3900
_|3900,3901
_|3901,3902
yo|3903,3905
female|3906,3912
with|3913,3917
a|3918,3919
history|3920,3927
of|3928,3930
CAD|3931,3934
who|3935,3938
<EOL>|3939,3940
presented|3940,3949
with|3950,3954
an|3955,3957
STEMI|3958,3963
s|3964,3965
/|3965,3966
p|3966,3967
catheterization|3968,3983
and|3984,3987
was|3988,3991
incidentally|3992,4004
<EOL>|4005,4006
found|4006,4011
to|4012,4014
have|4015,4019
multiple|4020,4028
pulmonary|4029,4038
nodules|4039,4046
consistent|4047,4057
with|4058,4062
<EOL>|4063,4064
adenocarcinoma|4064,4078
.|4078,4079
<EOL>|4081,4082
<EOL>|4082,4083
#|4083,4084
.|4084,4085
STEMI|4086,4091
:|4091,4092
Pt|4093,4095
presented|4096,4105
with|4106,4110
an|4111,4113
anterior|4114,4122
STEMI|4123,4128
.|4128,4129
Her|4131,4134
TIMI|4135,4139
risk|4140,4144
<EOL>|4145,4146
score|4146,4151
was|4152,4155
7|4156,4157
indicating|4158,4168
a|4169,4170
41|4171,4173
%|4173,4174
risk|4175,4179
at|4180,4182
14|4183,4185
days|4186,4190
of|4191,4193
mortality|4194,4203
,|4203,4204
new|4205,4208
<EOL>|4209,4210
or|4210,4212
recurrent|4213,4222
MI|4223,4225
,|4225,4226
or|4227,4229
severe|4230,4236
recurrent|4237,4246
ischemia|4247,4255
requiring|4256,4265
urgent|4266,4272
<EOL>|4273,4274
revascularization|4274,4291
.|4291,4292
Her|4294,4297
SVG|4298,4301
found|4302,4307
to|4308,4310
be|4311,4313
completely|4314,4324
occluded|4325,4333
and|4334,4337
<EOL>|4338,4339
a|4339,4340
BMS|4341,4344
was|4345,4348
placed|4349,4355
in|4356,4358
the|4359,4362
proximal|4363,4371
LAD|4372,4375
.|4375,4376
Due|4378,4381
to|4382,4384
the|4385,4388
timing|4389,4395
of|4396,4398
the|4399,4402
<EOL>|4403,4404
SVG|4404,4407
placement|4408,4417
over|4418,4422
_|4423,4424
_|4424,4425
_|4425,4426
years|4427,4432
ago|4433,4436
,|4436,4437
it|4438,4440
was|4441,4444
thought|4445,4452
that|4453,4457
her|4458,4461
LAD|4462,4465
had|4466,4469
<EOL>|4470,4471
managed|4471,4478
to|4479,4481
self|4482,4486
revascularize|4487,4500
and|4501,4504
was|4505,4508
partially|4509,4518
supplied|4519,4527
by|4528,4530
the|4531,4534
<EOL>|4535,4536
RCA|4536,4539
.|4539,4540
She|4542,4545
was|4546,4549
started|4550,4557
on|4558,4560
routine|4561,4568
ACS|4569,4572
medications|4573,4584
:|4584,4585
eptifibatide|4586,4598
<EOL>|4599,4600
for|4600,4603
18|4604,4606
hrs|4607,4610
,|4610,4611
plavix|4612,4618
75|4619,4621
and|4622,4625
aspirin|4626,4633
325mg|4634,4639
,|4639,4640
metoprolol|4641,4651
,|4651,4652
captopril|4653,4662
,|4662,4663
<EOL>|4664,4665
and|4665,4668
atorvastatin|4669,4681
.|4681,4682
Cardiac|4684,4691
enzymes|4692,4699
trended|4700,4707
down|4708,4712
appropriately|4713,4726
<EOL>|4727,4728
with|4728,4732
peak|4733,4737
Ck|4738,4740
and|4741,4744
CKMB|4745,4749
at|4750,4752
107|4753,4756
and|4757,4760
18.2|4761,4765
.|4765,4766
There|4768,4773
was|4774,4777
concern|4778,4785
for|4786,4789
<EOL>|4790,4791
acute|4791,4796
heart|4797,4802
failure|4803,4810
from|4811,4815
ischemic|4816,4824
insult|4825,4831
oxygen|4832,4838
requirement|4839,4850
.|4850,4851
<EOL>|4853,4854
However|4854,4861
,|4861,4862
she|4863,4866
was|4867,4870
noted|4871,4876
to|4877,4879
also|4880,4884
have|4885,4889
a|4890,4891
RLL|4892,4895
pneumonia|4896,4905
and|4906,4909
no|4910,4912
<EOL>|4913,4914
significant|4914,4925
pulmonary|4926,4935
edema|4936,4941
(|4942,4943
see|4943,4946
below|4947,4952
)|4952,4953
.|4953,4954
ECHO|4956,4960
showed|4961,4967
moderate|4968,4976
<EOL>|4977,4978
to|4978,4980
severe|4981,4987
regional|4988,4996
left|4997,5001
ventricular|5002,5013
systolic|5014,5022
dysfunction|5023,5034
with|5035,5039
<EOL>|5040,5041
anterior|5041,5049
and|5050,5053
anterospetal|5054,5066
akinesis|5067,5075
and|5076,5079
inferior|5080,5088
/|5088,5089
inferolateral|5089,5102
<EOL>|5103,5104
hypokinesis|5104,5115
.|5115,5116
Initially|5118,5127
,|5127,5128
patient|5129,5136
was|5138,5141
started|5142,5149
on|5150,5152
coumadin|5153,5161
for|5162,5165
<EOL>|5166,5167
ventricular|5167,5178
thrombus|5179,5187
prophylaxis|5188,5199
,|5199,5200
but|5201,5204
this|5205,5209
was|5210,5213
subsequantly|5214,5226
<EOL>|5227,5228
discontinued|5228,5240
as|5241,5243
risk|5244,5248
of|5249,5251
bleeding|5252,5260
outweighed|5261,5271
benefit|5272,5279
.|5279,5280
<EOL>|5281,5282
<EOL>|5282,5283
#|5283,5284
Hypoxia|5285,5292
:|5292,5293
Upon|5295,5299
hospitalization|5300,5315
,|5315,5316
patient|5317,5324
was|5325,5328
maintaing|5329,5338
<EOL>|5339,5340
saturations|5340,5351
in|5352,5354
low|5355,5358
_|5359,5360
_|5360,5361
_|5361,5362
on|5363,5365
6L|5366,5368
from|5369,5373
baseline|5374,5382
92|5383,5385
%|5385,5386
on|5387,5389
RA|5390,5392
.|5392,5393
CXR|5395,5398
<EOL>|5399,5400
showed|5400,5406
RLL|5407,5410
pneumonia|5411,5420
,|5420,5421
and|5422,5425
patient|5426,5433
was|5434,5437
subsequantly|5438,5450
started|5451,5458
on|5459,5461
<EOL>|5462,5463
ceftriaxone|5463,5474
,|5474,5475
azithromycin|5476,5488
,|5488,5489
metronidazole|5490,5503
.|5503,5504
As|5506,5508
the|5509,5512
patient|5513,5520
had|5521,5524
<EOL>|5525,5526
history|5526,5533
recurrent|5534,5543
RLL|5544,5547
pneumonia|5548,5557
,|5557,5558
a|5559,5560
CT|5561,5563
scan|5564,5568
was|5569,5572
obtained|5573,5581
which|5582,5587
<EOL>|5588,5589
showed|5589,5595
severe|5596,5602
right|5603,5608
lower|5609,5614
lobe|5615,5619
consolidation|5620,5633
and|5634,5637
extensive|5638,5647
,|5647,5648
new|5649,5652
<EOL>|5653,5654
diffuse|5654,5661
lung|5662,5666
nodules|5667,5674
with|5675,5679
sputum|5681,5687
cytology|5688,5696
positive|5697,5705
for|5706,5709
<EOL>|5710,5711
adenocarcinoma|5711,5725
.|5725,5726
Hypoxia|5728,5735
was|5736,5739
initially|5740,5749
felt|5750,5754
to|5755,5757
be|5758,5760
a|5761,5762
combination|5763,5774
<EOL>|5775,5776
of|5776,5778
postobstructive|5779,5794
pneumonia|5795,5804
and|5805,5808
tumor|5809,5814
burden|5815,5821
from|5822,5826
<EOL>|5827,5828
adenocarcinoma|5828,5842
.|5842,5843
Antibiotics|5845,5856
were|5857,5861
changed|5862,5869
to|5870,5872
vancomycin|5873,5883
,|5883,5884
<EOL>|5885,5886
levofloxacin|5886,5898
and|5899,5902
flagyl|5903,5909
of|5910,5912
which|5913,5918
she|5919,5922
completed|5923,5932
a|5933,5934
10|5935,5937
day|5938,5941
course|5942,5948
.|5948,5949
<EOL>|5951,5952
Repeat|5952,5958
CT|5959,5961
scan|5962,5966
showed|5967,5973
little|5974,5980
interval|5981,5989
improvement|5990,6001
in|6002,6004
right|6005,6010
lower|6011,6016
<EOL>|6017,6018
lobe|6018,6022
infiltrate|6023,6033
.|6033,6034
Respiratory|6036,6047
status|6048,6054
remained|6055,6063
tenuous|6064,6071
,|6071,6072
patient|6073,6080
<EOL>|6081,6082
requiring|6082,6091
high|6092,6096
flow|6097,6101
O2|6102,6104
with|6105,6109
6LNC|6110,6114
with|6115,6119
desaturations|6120,6133
to|6134,6136
high|6137,6141
_|6142,6143
_|6143,6144
_|6144,6145
<EOL>|6146,6147
with|6147,6151
activity|6152,6160
.|6160,6161
Prior|6163,6168
to|6169,6171
discharge|6172,6181
O2|6182,6184
requirement|6185,6196
was|6197,6200
5L|6201,6203
by|6204,6206
<EOL>|6207,6208
nasal|6208,6213
cannula|6214,6221
.|6221,6222
She|6224,6227
was|6228,6231
breathing|6232,6241
comfortably|6242,6253
with|6254,6258
oxygen|6259,6265
<EOL>|6266,6267
saturation|6267,6277
in|6278,6280
the|6281,6284
low|6285,6288
_|6289,6290
_|6290,6291
_|6291,6292
.|6292,6293
Likely|6295,6301
this|6302,6306
will|6307,6311
continue|6312,6320
to|6321,6323
be|6324,6326
<EOL>|6327,6328
necessary|6328,6337
for|6338,6341
some|6342,6346
time|6347,6351
.|6351,6352
A|6354,6355
shovel|6356,6362
mask|6363,6367
may|6368,6371
be|6372,6374
used|6375,6379
to|6380,6382
assist|6383,6389
<EOL>|6390,6391
with|6391,6395
oxygenation|6396,6407
as|6408,6410
needed|6411,6417
.|6417,6418
<EOL>|6423,6424
<EOL>|6424,6425
#|6425,6426
Lung|6427,6431
nodules|6432,6439
/|6439,6440
Broncheoalveolar|6441,6457
carcinoma|6458,6467
:|6467,6468
CT|6469,6471
scan|6472,6476
with|6477,6481
diffuse|6482,6489
<EOL>|6490,6491
pulmonary|6491,6500
nodules|6501,6508
and|6509,6512
sputum|6513,6519
cytology|6520,6528
positive|6529,6537
for|6538,6541
<EOL>|6542,6543
adenocarcinoma|6543,6557
.|6557,6558
Etiology|6560,6568
was|6569,6572
felt|6573,6577
to|6578,6580
be|6581,6583
primary|6584,6591
<EOL>|6592,6593
bronchioalveolar|6593,6609
vs|6610,6612
metastatic|6613,6623
thyroid|6624,6631
dx|6632,6634
(|6635,6636
prior|6636,6641
dx|6642,6644
of|6645,6647
possible|6648,6656
<EOL>|6657,6658
microfollicular|6658,6673
carcinoma|6674,6683
)|6683,6684
although|6685,6693
routine|6694,6701
cancer|6702,6708
screening|6709,6718
was|6719,6722
<EOL>|6723,6724
not|6724,6727
up|6728,6730
-|6730,6731
to|6731,6733
-|6733,6734
date|6734,6738
.|6738,6739
A|6741,6742
tissue|6743,6749
diagnosis|6750,6759
was|6760,6763
not|6764,6767
attained|6768,6776
given|6777,6782
the|6783,6786
<EOL>|6787,6788
patient|6788,6795
's|6795,6797
high|6798,6802
oxygen|6803,6809
requirement|6810,6821
and|6822,6825
anticoagulation|6826,6841
with|6842,6846
<EOL>|6847,6848
plavix|6848,6854
/|6854,6855
asa|6855,6858
in|6859,6861
the|6862,6865
setting|6866,6873
of|6874,6876
recent|6877,6883
_|6884,6885
_|6885,6886
_|6886,6887
placement|6888,6897
.|6897,6898
Although|6900,6908
<EOL>|6909,6910
patient|6910,6917
did|6918,6921
not|6922,6925
have|6926,6930
imaging|6931,6938
of|6939,6941
her|6942,6945
head|6946,6950
,|6950,6951
staging|6952,6959
based|6960,6965
on|6966,6968
CT|6969,6971
<EOL>|6972,6973
torso|6973,6978
was|6979,6982
IIIa|6983,6987
with|6988,6992
pulmonary|6993,7002
nodules|7003,7010
in|7011,7013
both|7014,7018
lung|7019,7023
fields|7024,7030
<EOL>|7031,7032
without|7032,7039
obvious|7040,7047
distal|7048,7054
LAD|7055,7058
or|7059,7061
metastasis|7062,7072
.|7072,7073
Empiric|7075,7082
therapy|7083,7090
with|7091,7095
<EOL>|7096,7097
single|7097,7103
agent|7104,7109
chemotherapy|7110,7122
was|7123,7126
initiated|7127,7136
on|7137,7139
_|7140,7141
_|7141,7142
_|7142,7143
with|7144,7148
<EOL>|7149,7150
Pemetrexed|7150,7160
.|7160,7161
She|7163,7166
tolerated|7167,7176
this|7177,7181
well|7182,7186
.|7186,7187
She|7189,7192
received|7193,7201
<EOL>|7202,7203
dexamethasone|7203,7216
on|7217,7219
_|7220,7221
_|7221,7222
_|7222,7223
to|7224,7226
prevent|7227,7234
rash|7235,7239
.|7239,7240
<EOL>|7243,7244
<EOL>|7244,7245
#|7245,7246
Chronic|7247,7254
renal|7255,7260
insufficiency|7261,7274
-|7275,7276
Patient|7277,7284
with|7285,7289
GFR|7290,7293
48|7294,7296
.|7296,7297
<EOL>|7299,7300
Medications|7300,7311
were|7312,7316
renally|7317,7324
dosed|7325,7330
and|7331,7334
renal|7335,7340
function|7341,7349
was|7350,7353
carefully|7354,7363
<EOL>|7364,7365
followed|7365,7373
.|7373,7374
She|7376,7379
was|7380,7383
treated|7384,7391
prophylactically|7392,7408
with|7409,7413
mucomyst|7414,7422
prior|7423,7428
<EOL>|7429,7430
to|7430,7432
and|7433,7436
post|7437,7441
IV|7442,7444
contrast|7445,7453
dose|7454,7458
.|7458,7459
Creatinine|7461,7471
remained|7472,7480
stable|7481,7487
at|7488,7490
<EOL>|7491,7492
_|7492,7493
_|7493,7494
_|7494,7495
.|7495,7496
<EOL>|7498,7499
<EOL>|7499,7500
#|7500,7501
Hyperkalemia|7502,7514
:|7514,7515
The|7517,7520
patient|7521,7528
was|7529,7532
mildly|7533,7539
hyperkalemic|7540,7552
the|7553,7556
day|7557,7560
<EOL>|7561,7562
prior|7562,7567
to|7568,7570
discharge|7571,7580
to|7581,7583
5.6|7584,7587
without|7588,7595
EKG|7596,7599
changes|7600,7607
.|7607,7608
This|7611,7615
responded|7616,7625
<EOL>|7626,7627
promptly|7627,7635
to|7636,7638
kayexalate|7639,7649
.|7649,7650
Electrolytes|7652,7664
should|7665,7671
be|7672,7674
checked|7675,7682
daily|7683,7688
<EOL>|7689,7690
until|7690,7695
stable|7696,7702
.|7702,7703
If|7705,7707
necessary|7708,7717
ACEI|7718,7722
could|7723,7728
be|7729,7731
stopped|7732,7739
.|7739,7740
<EOL>|7740,7741
<EOL>|7741,7742
#|7742,7743
HTN|7744,7747
:|7747,7748
She|7750,7753
was|7754,7757
normotensive|7758,7770
on|7771,7773
ACEI|7774,7778
and|7779,7782
b|7783,7784
-|7784,7785
blocker|7785,7792
.|7792,7793
<EOL>|7795,7796
<EOL>|7796,7797
<EOL>|7798,7799
Medications|7799,7810
on|7811,7813
Admission|7814,7823
:|7823,7824
<EOL>|7824,7825
#|7825,7826
Clopidogrel|7827,7838
[|7839,7840
Plavix|7840,7846
]|7846,7847
75|7848,7850
mg|7851,7853
Tablet|7854,7860
PO|7861,7863
Daily|7864,7869
<EOL>|7869,7870
#|7870,7871
Ezetimibe|7872,7881
-|7881,7882
Simvastatin|7882,7893
[|7894,7895
Vytorin|7895,7902
_|7903,7904
_|7904,7905
_|7905,7906
10|7907,7909
mg|7910,7912
-|7912,7913
20|7913,7915
mg|7916,7918
PO|7919,7921
daily|7922,7927
<EOL>|7932,7933
<EOL>|7934,7935
#|7935,7936
Nifedipine|7937,7947
30|7948,7950
mg|7951,7953
SR|7954,7956
PO|7957,7959
qday|7960,7964
<EOL>|7964,7965
#|7965,7966
Nitroglycerin|7967,7980
0.4|7981,7984
mg|7985,7987
/|7987,7988
hour|7988,7992
Patch|7993,7998
24|7999,8001
hr|8002,8004
1|8005,8006
patch|8007,8012
once|8013,8017
a|8018,8019
day|8020,8023
<EOL>|8026,8027
#|8027,8028
Nitroglycern|8029,8041
sublingual|8042,8052
tabs|8053,8057
PRN|8058,8061
-|8062,8063
has|8064,8067
not|8068,8071
used|8072,8076
recently|8077,8085
prior|8086,8091
<EOL>|8092,8093
to|8093,8095
today|8096,8101
<EOL>|8101,8102
#|8102,8103
Propranolol|8104,8115
80|8116,8118
mg|8119,8121
Tablet|8122,8128
PO|8129,8131
once|8132,8136
a|8137,8138
day|8139,8142
<EOL>|8152,8153
#|8153,8154
Multivitamin|8155,8167
<EOL>|8167,8168
<EOL>|8169,8170
Discharge|8170,8179
Disposition|8180,8191
:|8191,8192
<EOL>|8192,8193
Extended|8193,8201
Care|8202,8206
<EOL>|8206,8207
<EOL>|8208,8209
Facility|8209,8217
:|8217,8218
<EOL>|8218,8219
_|8219,8220
_|8220,8221
_|8221,8222
<EOL>|8222,8223
<EOL>|8224,8225
Discharge|8225,8234
Diagnosis|8235,8244
:|8244,8245
<EOL>|8245,8246
Primary|8246,8253
:|8253,8254
<EOL>|8254,8255
ST|8255,8257
elevation|8258,8267
myocardial|8268,8278
infarction|8279,8289
<EOL>|8289,8290
Presumed|8290,8298
broncheoalveolar|8299,8315
carcinoma|8316,8325
<EOL>|8325,8326
<EOL>|8326,8327
<EOL>|8328,8329
Discharge|8329,8338
Condition|8339,8348
:|8348,8349
<EOL>|8349,8350
stable|8350,8356
,|8356,8357
with|8358,8362
5L|8363,8365
oxygen|8366,8372
requirement|8373,8384
and|8385,8388
O2|8389,8391
Sat|8392,8395
in|8396,8398
the|8399,8402
low|8403,8406
_|8407,8408
_|8408,8409
_|8409,8410
<EOL>|8410,8411
<EOL>|8411,8412
<EOL>|8413,8414
Discharge|8414,8423
Instructions|8424,8436
:|8436,8437
<EOL>|8437,8438
You|8438,8441
were|8442,8446
admitted|8447,8455
to|8456,8458
the|8459,8462
hospital|8463,8471
for|8472,8475
chest|8476,8481
pressure|8482,8490
and|8491,8494
found|8495,8500
<EOL>|8501,8502
to|8502,8504
have|8505,8509
a|8510,8511
heart|8512,8517
attack|8518,8524
.|8524,8525
You|8527,8530
had|8531,8534
a|8535,8536
cardiac|8537,8544
catheterization|8545,8560
and|8561,8564
<EOL>|8565,8566
had|8566,8569
a|8570,8571
bare|8572,8576
metal|8577,8582
stent|8583,8588
placed|8589,8595
.|8595,8596
After|8598,8603
this|8604,8608
,|8608,8609
you|8610,8613
had|8614,8617
some|8618,8622
trouble|8623,8630
<EOL>|8631,8632
breathing|8632,8641
and|8642,8645
had|8646,8649
a|8650,8651
scan|8652,8656
that|8657,8661
showed|8662,8668
some|8669,8673
nodules|8674,8681
in|8682,8684
your|8685,8689
lungs|8690,8695
.|8695,8696
<EOL>|8697,8698
A|8699,8700
sputum|8701,8707
sample|8708,8714
was|8715,8718
sent|8719,8723
and|8724,8727
malignant|8728,8737
cells|8738,8743
were|8744,8748
seen|8749,8753
.|8753,8754
This|8755,8759
<EOL>|8760,8761
was|8761,8764
thought|8765,8772
to|8773,8775
be|8776,8778
broncheoalveolar|8779,8795
lung|8796,8800
cancer|8801,8807
,|8807,8808
and|8809,8812
you|8813,8816
were|8817,8821
<EOL>|8822,8823
treated|8823,8830
with|8831,8835
one|8836,8839
dose|8840,8844
of|8845,8847
chemotherapy|8848,8860
for|8861,8864
this|8865,8869
.|8869,8870
Please|8872,8878
<EOL>|8879,8880
follow|8880,8886
-|8886,8887
up|8887,8889
with|8890,8894
Dr.|8895,8898
_|8899,8900
_|8900,8901
_|8901,8902
to|8903,8905
determine|8906,8915
if|8916,8918
further|8919,8926
<EOL>|8927,8928
treatment|8928,8937
will|8938,8942
be|8943,8945
needed|8946,8952
.|8952,8953
<EOL>|8953,8954
<EOL>|8954,8955
Weigh|8955,8960
yourself|8961,8969
every|8970,8975
morning|8976,8983
,|8983,8984
call|8985,8989
MD|8990,8992
if|8993,8995
weight|8996,9002
goes|9003,9007
up|9008,9010
more|9011,9015
<EOL>|9016,9017
than|9017,9021
3|9022,9023
lbs|9024,9027
.|9027,9028
<EOL>|9028,9029
<EOL>|9029,9030
The|9030,9033
following|9034,9043
changes|9044,9051
were|9052,9056
made|9057,9061
to|9062,9064
your|9065,9069
medications|9070,9081
:|9081,9082
<EOL>|9082,9083
1|9083,9084
.|9084,9085
You|9086,9089
were|9090,9094
started|9095,9102
on|9103,9105
plavix|9106,9112
,|9112,9113
a|9114,9115
medication|9116,9126
to|9127,9129
thin|9130,9134
your|9135,9139
blood|9140,9145
.|9145,9146
<EOL>|9147,9148
You|9148,9151
must|9152,9156
take|9157,9161
this|9162,9166
medication|9167,9177
for|9178,9181
1|9182,9183
month|9184,9189
to|9190,9192
ensure|9193,9199
that|9200,9204
your|9205,9209
<EOL>|9210,9211
heart|9211,9216
stent|9217,9222
does|9223,9227
not|9228,9231
become|9232,9238
blocked|9239,9246
.|9246,9247
<EOL>|9247,9248
<EOL>|9248,9249
<EOL>|9250,9251
Followup|9251,9259
Instructions|9260,9272
:|9272,9273
<EOL>|9273,9274
_|9274,9275
_|9275,9276
_|9276,9277
<EOL>|9277,9278

