 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
Codeine|179,186
<EOL>|186,187
<EOL>|188,189
Attending|189,198
:|198,199
_|200,201
_|201,202
_|202,203
.|203,204
<EOL>|204,205
<EOL>|206,207
Chief|207,212
Complaint|213,222
:|222,223
<EOL>|223,224
Dyspnea|224,231
and|232,235
melena|236,242
<EOL>|243,244
<EOL>|245,246
Major|246,251
Surgical|252,260
or|261,263
Invasive|264,272
Procedure|273,282
:|282,283
<EOL>|283,284
None|284,288
<EOL>|288,289
<EOL>|290,291
History|291,298
of|299,301
Present|302,309
Illness|310,317
:|317,318
<EOL>|318,319
Ms.|319,322
_|323,324
_|324,325
_|325,326
is|327,329
a|330,331
_|332,333
_|333,334
_|334,335
F|336,337
with|338,342
history|343,350
of|351,353
stage|354,359
IV|360,362
non-small|363,372
<EOL>|373,374
cell|374,378
lung|379,383
cancer|384,390
,|390,391
CAD|392,395
and|396,399
CKD|400,403
who|404,407
presents|408,416
with|417,421
dyspnea|422,429
,|429,430
<EOL>|431,432
productive|432,442
cough|443,448
and|449,452
melena|453,459
.|459,460
Patient|461,468
has|469,472
had|473,476
_|477,478
_|478,479
_|479,480
days|481,485
of|486,488
melena|489,495
<EOL>|496,497
without|497,504
abdominal|505,514
pain|515,519
and|520,523
dyspnea|524,531
with|532,536
worsening|537,546
cough|547,552
for|553,556
the|557,560
<EOL>|561,562
past|562,566
day|567,570
.|570,571
She|572,575
denies|576,582
fevers|583,589
or|590,592
chest|593,598
pain|599,603
.|603,604
<EOL>|606,607
.|607,608
<EOL>|610,611
In|611,613
the|614,617
ER|618,620
,|620,621
initial|622,629
vitals|630,636
were|637,641
97.2|642,646
,|646,647
89|648,650
,|650,651
156|652,655
/|655,656
53|656,658
,|658,659
22|660,662
,|662,663
86|664,666
%|666,667
4L|668,670
.|670,671
Her|672,675
<EOL>|676,677
hct|677,680
was|681,684
22|685,687
from|688,692
recent|693,699
baseline|700,708
of|709,711
25|712,714
(|715,716
she|716,719
has|720,723
transfusion|724,735
<EOL>|736,737
dependent|737,746
anemia|747,753
)|753,754
,|754,755
and|756,759
she|760,763
initially|764,773
was|774,777
hypoxic|778,785
.|785,786
ABG|787,790
was|791,794
<EOL>|795,796
7.29|796,800
/|800,801
64|801,803
/|803,804
42|804,806
/|806,807
32|807,809
and|810,813
lactate|814,821
was|822,825
2.4|826,829
.|829,830
Patient|831,838
responded|839,848
to|849,851
nebs|852,856
,|856,857
<EOL>|858,859
stress|859,865
dose|866,870
steroids|871,879
,|879,880
levaquin|881,889
and|890,893
ceftriaxone|894,905
with|906,910
improvement|911,922
<EOL>|923,924
in|924,926
her|927,930
sats|931,935
to|936,938
mid|939,942
_|943,944
_|944,945
_|945,946
on|947,949
5L|950,952
NC|953,955
.|955,956
She|957,960
was|961,964
started|965,972
on|973,975
IV|976,978
PPI|979,982
for|983,986
<EOL>|987,988
her|988,991
guaiac|992,998
positive|999,1007
dark|1008,1012
brown|1013,1018
stool|1019,1024
.|1024,1025
CXR|1026,1029
showed|1030,1036
large|1037,1042
R|1043,1044
pleural|1045,1052
<EOL>|1053,1054
effusion|1054,1062
and|1063,1066
questionable|1067,1079
L|1080,1081
lower|1082,1087
lobe|1088,1092
collapse|1093,1101
.|1101,1102
EKG|1103,1106
showed|1107,1113
<EOL>|1114,1115
sinus|1115,1120
tach|1121,1125
with|1126,1130
ST|1131,1133
depressions|1134,1145
in|1146,1148
V2|1149,1151
-|1151,1152
6|1152,1153
.|1153,1154
Vitals|1155,1161
on|1162,1164
transfer|1165,1173
to|1174,1176
<EOL>|1177,1178
the|1178,1181
MICU|1182,1186
were|1187,1191
97.2|1192,1196
,|1196,1197
105|1198,1201
,|1201,1202
127|1203,1206
/|1206,1207
50|1207,1209
,|1209,1210
29|1211,1213
,|1213,1214
96|1215,1217
%|1217,1218
5L|1219,1221
NC|1222,1224
.|1224,1225
<EOL>|1227,1228
.|1228,1229
<EOL>|1231,1232
In|1232,1234
the|1235,1238
MICU|1239,1243
,|1243,1244
she|1245,1248
reports|1249,1256
feeling|1257,1264
better|1265,1271
after|1272,1277
her|1278,1281
breathing|1282,1291
<EOL>|1292,1293
treatments|1293,1303
today|1304,1309
.|1309,1310
She|1311,1314
can|1315,1318
not|1318,1321
recall|1322,1328
when|1329,1333
her|1334,1337
difficulty|1338,1348
<EOL>|1349,1350
breathing|1350,1359
started|1360,1367
and|1368,1371
per|1372,1375
her|1376,1379
family|1380,1386
,|1386,1387
she|1388,1391
has|1392,1395
difficulty|1396,1406
hearing|1407,1414
<EOL>|1415,1416
but|1416,1419
no|1420,1422
memory|1423,1429
loss|1430,1434
.|1434,1435
Patient|1436,1443
had|1444,1447
intermittent|1448,1460
dyspnea|1461,1468
for|1469,1472
weeks|1473,1478
<EOL>|1479,1480
for|1480,1483
which|1484,1489
she|1490,1493
previously|1494,1504
took|1505,1509
codeine|1510,1517
syrup|1518,1523
but|1524,1527
then|1528,1532
a|1533,1534
period|1535,1541
of|1542,1544
<EOL>|1545,1546
improvement|1546,1557
.|1557,1558
She|1559,1562
developed|1563,1572
worsening|1573,1582
dypsnea|1583,1590
and|1591,1594
cough|1595,1600
yesterday|1601,1610
<EOL>|1611,1612
without|1612,1619
fevers|1620,1626
,|1626,1627
chills|1628,1634
or|1635,1637
chest|1638,1643
pain|1644,1648
.|1648,1649
She|1650,1653
denies|1654,1660
prior|1661,1666
history|1667,1674
<EOL>|1675,1676
of|1676,1678
melena|1679,1685
but|1686,1689
has|1690,1693
had|1694,1697
stable|1698,1704
nausea|1705,1711
and|1712,1715
poor|1716,1720
appetite|1721,1729
for|1730,1733
<EOL>|1734,1735
months|1735,1741
.|1741,1742
No|1743,1745
heartburn|1746,1755
or|1756,1758
dysphagia|1759,1768
.|1768,1769
<EOL>|1771,1772
<EOL>|1772,1773
<EOL>|1774,1775
Past|1775,1779
Medical|1780,1787
History|1788,1795
:|1795,1796
<EOL>|1796,1797
Stage|1797,1802
IV|1803,1805
nonsmall|1806,1814
cell|1815,1819
lung|1820,1824
cancer|1825,1831
,|1831,1832
adenocarcinoma|1833,1847
,|1847,1848
EGFR|1849,1853
<EOL>|1854,1855
wild|1855,1859
-|1859,1860
type|1860,1864
,|1864,1865
KRAS|1866,1870
mutated|1871,1878
<EOL>|1880,1881
CAD|1881,1884
s|1885,1886
/|1886,1887
p|1887,1888
CABG|1889,1893
in|1894,1896
_|1897,1898
_|1898,1899
_|1899,1900
,|1900,1901
MI|1902,1904
_|1905,1906
_|1906,1907
_|1907,1908
s|1909,1910
/|1910,1911
p|1911,1912
PCI|1913,1916
to|1917,1919
LAD|1920,1923
.|1923,1924
<EOL>|1926,1927
Chronic|1927,1934
renal|1935,1940
insufficiency|1941,1954
-|1955,1956
Patient|1957,1964
with|1965,1969
GFR|1970,1973
<|1974,1975
50|1976,1978
.|1978,1979
<EOL>|1981,1982
CVA|1982,1985
-|1986,1987
small|1988,1993
left|1994,1998
posterior|1999,2008
frontal|2009,2016
infarct|2017,2024
in|2025,2027
_|2028,2029
_|2029,2030
_|2030,2031
.|2031,2032
<EOL>|2034,2035
Hypercholesterolemia|2035,2055
.|2055,2056
<EOL>|2058,2059
Macular|2059,2066
Degeneration|2067,2079
<EOL>|2081,2082
<EOL>|2082,2083
<EOL>|2084,2085
Social|2085,2091
History|2092,2099
:|2099,2100
<EOL>|2100,2101
_|2101,2102
_|2102,2103
_|2103,2104
<EOL>|2104,2105
Family|2105,2111
History|2112,2119
:|2119,2120
<EOL>|2120,2121
Her|2121,2124
father|2125,2131
died|2132,2136
due|2137,2140
to|2141,2143
CAD|2144,2147
at|2148,2150
age|2151,2154
_|2155,2156
_|2156,2157
_|2157,2158
.|2158,2159
Her|2160,2163
mother|2164,2170
had|2171,2174
stomach|2175,2182
<EOL>|2184,2185
cancer|2185,2191
and|2192,2195
osteosarcoma|2196,2208
.|2208,2209
<EOL>|2211,2212
<EOL>|2212,2213
<EOL>|2214,2215
Physical|2215,2223
Exam|2224,2228
:|2228,2229
<EOL>|2229,2230
General|2230,2237
:|2237,2238
Elderly|2239,2246
,|2246,2247
chronically|2248,2259
ill|2260,2263
appearing|2264,2273
female|2274,2280
in|2281,2283
NAD|2284,2287
<EOL>|2289,2290
HEENT|2290,2295
:|2295,2296
NC|2297,2299
/|2299,2300
AT|2300,2302
,|2302,2303
EOMI|2304,2308
,|2308,2309
sclera|2310,2316
anicteric|2317,2326
,|2326,2327
MMM|2328,2331
<EOL>|2333,2334
Neck|2334,2338
:|2338,2339
supple|2340,2346
,|2346,2347
JVP|2348,2351
not|2352,2355
elevated|2356,2364
,|2364,2365
1|2366,2367
+|2367,2368
firm|2369,2373
bilateral|2374,2383
submandibular|2384,2397
<EOL>|2398,2399
LAD|2399,2402
<EOL>|2404,2405
Lungs|2405,2410
:|2410,2411
Decreased|2412,2421
percussion|2422,2432
_|2433,2434
_|2434,2435
_|2435,2436
way|2437,2440
up|2441,2443
right|2444,2449
lung|2450,2454
with|2455,2459
decreased|2460,2469
<EOL>|2470,2471
breath|2471,2477
sounds|2478,2484
,|2484,2485
L|2486,2487
basalar|2488,2495
crackles|2496,2504
,|2504,2505
upper|2506,2511
lobes|2512,2517
with|2518,2522
some|2523,2527
mild|2528,2532
<EOL>|2533,2534
wheezing|2534,2542
<EOL>|2544,2545
CV|2545,2547
:|2547,2548
Regular|2549,2556
rate|2557,2561
and|2562,2565
rhythm|2566,2572
,|2572,2573
normal|2574,2580
S1|2581,2583
+|2584,2585
S2|2586,2588
,|2588,2589
no|2590,2592
murmurs|2593,2600
,|2600,2601
rubs|2602,2606
,|2606,2607
<EOL>|2608,2609
gallops|2609,2616
appreciated|2617,2628
<EOL>|2630,2631
Abdomen|2631,2638
:|2638,2639
soft|2640,2644
,|2644,2645
non-tender|2646,2656
,|2656,2657
non-distended|2658,2671
,|2671,2672
bowel|2673,2678
sounds|2679,2685
present|2686,2693
,|2693,2694
<EOL>|2695,2696
no|2696,2698
rebound|2699,2706
tenderness|2707,2717
or|2718,2720
guarding|2721,2729
,|2729,2730
no|2731,2733
organomegaly|2734,2746
<EOL>|2748,2749
GU|2749,2751
:|2751,2752
no|2753,2755
foley|2756,2761
<EOL>|2763,2764
Ext|2764,2767
:|2767,2768
warm|2769,2773
,|2773,2774
well|2775,2779
perfused|2780,2788
,|2788,2789
2|2790,2791
+|2791,2792
pulses|2793,2799
,|2799,2800
no|2801,2803
clubbing|2804,2812
,|2812,2813
cyanosis|2814,2822
or|2823,2825
<EOL>|2826,2827
edema|2827,2832
<EOL>|2834,2835
<EOL>|2835,2836
Discharge|2836,2845
:|2845,2846
<EOL>|2846,2847
expired|2847,2854
<EOL>|2854,2855
<EOL>|2856,2857
Pertinent|2857,2866
Results|2867,2874
:|2874,2875
<EOL>|2875,2876
_|2876,2877
_|2877,2878
_|2878,2879
07|2880,2882
:|2882,2883
42PM|2883,2887
BLOOD|2888,2893
WBC|2894,2897
-|2897,2898
9|2898,2899
.|2899,2900
8|2900,2901
#|2901,2902
RBC|2903,2906
-|2906,2907
2|2907,2908
.|2908,2909
60|2909,2911
*|2911,2912
Hgb|2913,2916
-|2916,2917
7|2917,2918
.|2918,2919
5|2919,2920
*|2920,2921
Hct|2922,2925
-|2925,2926
22|2926,2928
.|2928,2929
4|2929,2930
*|2930,2931
<EOL>|2932,2933
MCV|2933,2936
-|2936,2937
86|2937,2939
MCH|2940,2943
-|2943,2944
28.7|2944,2948
MCHC|2949,2953
-|2953,2954
33.3|2954,2958
RDW|2959,2962
-|2962,2963
18|2963,2965
.|2965,2966
8|2966,2967
*|2967,2968
Plt|2969,2972
_|2973,2974
_|2974,2975
_|2975,2976
<EOL>|2976,2977
_|2977,2978
_|2978,2979
_|2979,2980
07|2981,2983
:|2983,2984
42PM|2984,2988
BLOOD|2989,2994
Neuts|2995,3000
-|3000,3001
83|3001,3003
.|3003,3004
0|3004,3005
*|3005,3006
Lymphs|3007,3013
-|3013,3014
8|3014,3015
.|3015,3016
5|3016,3017
*|3017,3018
Monos|3019,3024
-|3024,3025
5.7|3025,3028
Eos|3029,3032
-|3032,3033
2.4|3033,3036
<EOL>|3037,3038
Baso|3038,3042
-|3042,3043
0.4|3043,3046
<EOL>|3046,3047
_|3047,3048
_|3048,3049
_|3049,3050
07|3051,3053
:|3053,3054
42PM|3054,3058
BLOOD|3059,3064
_|3065,3066
_|3066,3067
_|3067,3068
PTT|3069,3072
-|3072,3073
24.5|3073,3077
_|3078,3079
_|3079,3080
_|3080,3081
<EOL>|3081,3082
_|3082,3083
_|3083,3084
_|3084,3085
07|3086,3088
:|3088,3089
42PM|3089,3093
BLOOD|3094,3099
Glucose|3100,3107
-|3107,3108
133|3108,3111
*|3111,3112
UreaN|3113,3118
-|3118,3119
45|3119,3121
*|3121,3122
Creat|3123,3128
-|3128,3129
1|3129,3130
.|3130,3131
4|3131,3132
*|3132,3133
Na|3134,3136
-|3136,3137
120|3137,3140
*|3140,3141
<EOL>|3142,3143
K|3143,3144
-|3144,3145
5|3145,3146
.|3146,3147
7|3147,3148
*|3148,3149
Cl|3150,3152
-|3152,3153
85|3153,3155
*|3155,3156
HCO3|3157,3161
-|3161,3162
26|3162,3164
AnGap|3165,3170
-|3170,3171
15|3171,3173
<EOL>|3173,3174
_|3174,3175
_|3175,3176
_|3176,3177
07|3178,3180
:|3180,3181
42PM|3181,3185
BLOOD|3186,3191
ALT|3192,3195
-|3195,3196
20|3196,3198
AST|3199,3202
-|3202,3203
24|3203,3205
LD|3206,3208
(|3208,3209
LDH|3209,3212
)|3212,3213
-|3213,3214
297|3214,3217
*|3217,3218
CK|3219,3221
(|3221,3222
CPK|3222,3225
)|3225,3226
-|3226,3227
73|3227,3229
<EOL>|3230,3231
AlkPhos|3231,3238
-|3238,3239
81|3239,3241
TotBili|3242,3249
-|3249,3250
0.3|3250,3253
<EOL>|3253,3254
_|3254,3255
_|3255,3256
_|3256,3257
07|3258,3260
:|3260,3261
42PM|3261,3265
BLOOD|3266,3271
CK|3272,3274
-|3274,3275
MB|3275,3277
-|3277,3278
4|3278,3279
cTropnT|3280,3287
-|3287,3288
<|3288,3289
0|3289,3290
.|3290,3291
01|3291,3293
<EOL>|3293,3294
_|3294,3295
_|3295,3296
_|3296,3297
02|3298,3300
:|3300,3301
04AM|3301,3305
BLOOD|3306,3311
CK|3312,3314
-|3314,3315
MB|3315,3317
-|3317,3318
10|3318,3320
MB|3321,3323
Indx|3324,3328
-|3328,3329
10|3329,3331
.|3331,3332
1|3332,3333
*|3333,3334
cTropnT|3335,3342
-|3342,3343
0|3343,3344
.|3344,3345
05|3345,3347
*|3347,3348
<EOL>|3348,3349
_|3349,3350
_|3350,3351
_|3351,3352
11|3353,3355
:|3355,3356
02PM|3356,3360
BLOOD|3361,3366
Calcium|3367,3374
-|3374,3375
8.4|3375,3378
Phos|3379,3383
-|3383,3384
2|3384,3385
.|3385,3386
6|3386,3387
*|3387,3388
Mg|3389,3391
-|3391,3392
1.8|3392,3395
<EOL>|3395,3396
_|3396,3397
_|3397,3398
_|3398,3399
07|3400,3402
:|3402,3403
42PM|3403,3407
BLOOD|3408,3413
Osmolal|3414,3421
-|3421,3422
268|3422,3425
*|3425,3426
<EOL>|3426,3427
_|3427,3428
_|3428,3429
_|3429,3430
07|3431,3433
:|3433,3434
42PM|3434,3438
BLOOD|3439,3444
_|3445,3446
_|3446,3447
_|3447,3448
pO2|3449,3452
-|3452,3453
42|3453,3455
*|3455,3456
pCO2|3457,3461
-|3461,3462
64|3462,3464
*|3464,3465
pH|3466,3468
-|3468,3469
7|3469,3470
.|3470,3471
29|3471,3473
*|3473,3474
<EOL>|3475,3476
calTCO2|3476,3483
-|3483,3484
32|3484,3486
*|3486,3487
Base|3488,3492
XS|3493,3495
-|3495,3496
1|3496,3497
Comment|3498,3505
-|3505,3506
GREEN|3506,3511
TOP|3512,3515
<EOL>|3515,3516
_|3516,3517
_|3517,3518
_|3518,3519
12|3520,3522
:|3522,3523
15AM|3523,3527
BLOOD|3528,3533
Type|3534,3538
-|3538,3539
ART|3539,3542
pO2|3543,3546
-|3546,3547
55|3547,3549
*|3549,3550
pCO2|3551,3555
-|3555,3556
43|3556,3558
pH|3559,3561
-|3561,3562
7|3562,3563
.|3563,3564
32|3564,3566
*|3566,3567
<EOL>|3568,3569
calTCO2|3569,3576
-|3576,3577
23|3577,3579
Base|3580,3584
XS|3585,3587
-|3587,3588
-|3588,3589
3|3589,3590
<EOL>|3590,3591
_|3591,3592
_|3592,3593
_|3593,3594
04|3595,3597
:|3597,3598
39AM|3598,3602
BLOOD|3603,3608
Lactate|3609,3616
-|3616,3617
4|3617,3618
.|3618,3619
2|3619,3620
*|3620,3621
<EOL>|3621,3622
_|3622,3623
_|3623,3624
_|3624,3625
01|3626,3628
:|3628,3629
46AM|3629,3633
BLOOD|3634,3639
Lactate|3640,3647
-|3647,3648
5|3648,3649
.|3649,3650
9|3650,3651
*|3651,3652
<EOL>|3652,3653
_|3653,3654
_|3654,3655
_|3655,3656
12|3657,3659
:|3659,3660
15AM|3660,3664
BLOOD|3665,3670
Lactate|3671,3678
-|3678,3679
7|3679,3680
.|3680,3681
7|3681,3682
*|3682,3683
<EOL>|3683,3684
_|3684,3685
_|3685,3686
_|3686,3687
07|3688,3690
:|3690,3691
42PM|3691,3695
BLOOD|3696,3701
Lactate|3702,3709
-|3709,3710
2|3710,3711
.|3711,3712
4|3712,3713
*|3713,3714
<EOL>|3714,3715
_|3715,3716
_|3716,3717
_|3717,3718
12|3719,3721
:|3721,3722
58AM|3722,3726
URINE|3727,3732
Color|3733,3738
-|3738,3739
Straw|3739,3744
Appear|3745,3751
-|3751,3752
Clear|3752,3757
Sp|3758,3760
_|3761,3762
_|3762,3763
_|3763,3764
<EOL>|3764,3765
_|3765,3766
_|3766,3767
_|3767,3768
12|3769,3771
:|3771,3772
58AM|3772,3776
URINE|3777,3782
Blood|3783,3788
-|3788,3789
NEG|3789,3792
Nitrite|3793,3800
-|3800,3801
NEG|3801,3804
Protein|3805,3812
-|3812,3813
TR|3813,3815
<EOL>|3816,3817
Glucose|3817,3824
-|3824,3825
NEG|3825,3828
Ketone|3829,3835
-|3835,3836
NEG|3836,3839
Bilirub|3840,3847
-|3847,3848
NEG|3848,3851
Urobiln|3852,3859
-|3859,3860
NEG|3860,3863
pH|3864,3866
-|3866,3867
5.0|3867,3870
Leuks|3871,3876
-|3876,3877
NEG|3877,3880
<EOL>|3880,3881
_|3881,3882
_|3882,3883
_|3883,3884
12|3885,3887
:|3887,3888
58AM|3888,3892
URINE|3893,3898
RBC|3899,3902
-|3902,3903
1|3903,3904
WBC|3905,3908
-|3908,3909
<|3909,3910
1|3910,3911
Bacteri|3912,3919
-|3919,3920
NONE|3920,3924
Yeast|3925,3930
-|3930,3931
NONE|3931,3935
<EOL>|3936,3937
Epi|3937,3940
-|3940,3941
<|3941,3942
1|3942,3943
<EOL>|3943,3944
_|3944,3945
_|3945,3946
_|3946,3947
12|3948,3950
:|3950,3951
58AM|3951,3955
URINE|3956,3961
CastGr|3962,3968
-|3968,3969
1|3969,3970
*|3970,3971
CastHy|3972,3978
-|3978,3979
1|3979,3980
*|3980,3981
<EOL>|3981,3982
_|3982,3983
_|3983,3984
_|3984,3985
12|3986,3988
:|3988,3989
58AM|3989,3993
URINE|3994,3999
Hours|4000,4005
-|4005,4006
RANDOM|4006,4012
Creat|4013,4018
-|4018,4019
65|4019,4021
Na|4022,4024
-|4024,4025
21|4025,4027
K|4028,4029
-|4029,4030
37|4030,4032
Cl|4033,4035
-|4035,4036
19|4036,4038
<EOL>|4038,4039
_|4039,4040
_|4040,4041
_|4041,4042
12|4043,4045
:|4045,4046
58AM|4046,4050
URINE|4051,4056
Osmolal|4057,4064
-|4064,4065
469|4065,4068
<EOL>|4068,4069
<EOL>|4069,4070
PCXR|4070,4074
:|4074,4075
Interval|4076,4084
enlargement|4085,4096
of|4097,4099
the|4100,4103
now|4104,4107
massive|4108,4115
right|4116,4121
pleural|4122,4129
<EOL>|4130,4131
effusion|4131,4139
.|4139,4140
<EOL>|4142,4143
Denser|4143,4149
and|4150,4153
larger|4154,4160
consolidation|4161,4174
of|4175,4177
the|4178,4181
left|4182,4186
lung|4187,4191
,|4191,4192
possibly|4193,4201
<EOL>|4202,4203
extension|4203,4212
of|4213,4215
tumor|4216,4221
or|4222,4224
focal|4225,4230
,|4230,4231
acute|4232,4237
infiltrate|4238,4248
,|4248,4249
or|4250,4252
combination|4253,4264
<EOL>|4265,4266
thereof|4266,4273
.|4273,4274
<EOL>|4275,4276
<EOL>|4276,4277
<EOL>|4278,4279
Brief|4279,4284
Hospital|4285,4293
Course|4294,4300
:|4300,4301
<EOL>|4301,4302
The|4302,4305
patient|4306,4313
was|4314,4317
admitted|4318,4326
to|4327,4329
the|4330,4333
MICU|4334,4338
and|4339,4342
placed|4343,4349
on|4350,4352
BiPAP|4353,4358
for|4359,4362
<EOL>|4363,4364
comfort|4364,4371
.|4371,4372
Her|4373,4376
outpt|4377,4382
.|4382,4383
oncologist|4384,4394
was|4395,4398
contacted|4399,4408
overnight|4409,4418
.|4418,4419
She|4420,4423
<EOL>|4424,4425
underwent|4425,4434
thoracentesis|4435,4448
for|4449,4452
palliation|4453,4463
with|4464,4468
significant|4469,4480
volume|4481,4487
<EOL>|4488,4489
taken|4489,4494
off|4495,4498
.|4498,4499
Palliative|4500,4510
care|4511,4515
was|4516,4519
consulted|4520,4529
and|4530,4533
the|4534,4537
decision|4538,4546
was|4547,4550
<EOL>|4551,4552
made|4552,4556
to|4557,4559
focus|4560,4565
on|4566,4568
comfort|4569,4576
.|4576,4577
Her|4578,4581
oncologist|4582,4592
visited|4593,4600
with|4601,4605
her|4606,4609
and|4610,4613
<EOL>|4614,4615
her|4615,4618
family|4619,4625
.|4625,4626
SHe|4627,4630
was|4631,4634
transitioned|4635,4647
out|4648,4651
of|4652,4654
the|4655,4658
ICU|4659,4662
and|4663,4666
expired|4667,4674
on|4675,4677
<EOL>|4678,4679
the|4679,4682
floor|4683,4688
soon|4689,4693
after|4694,4699
.|4699,4700
<EOL>|4701,4702
<EOL>|4703,4704
Medications|4704,4715
on|4716,4718
Admission|4719,4728
:|4728,4729
<EOL>|4729,4730
Robitussin|4730,4740
with|4741,4745
codeine|4746,4753
_|4754,4755
_|4755,4756
_|4756,4757
tsp|4758,4761
QHS|4762,4765
<EOL>|4767,4768
ATORVASTATIN|4768,4780
[|4781,4782
LIPITOR|4782,4789
]|4789,4790
-|4791,4792
80|4793,4795
mg|4796,4798
Tablet|4799,4805
-|4806,4807
one|4808,4811
Tablet|4812,4818
(|4818,4819
s|4819,4820
)|4820,4821
by|4822,4824
mouth|4825,4830
<EOL>|4832,4833
one|4833,4836
daily|4837,4842
-|4843,4844
No|4845,4847
Substitution|4848,4860
<EOL>|4862,4863
BENZONATATE|4863,4874
-|4875,4876
100|4877,4880
mg|4881,4883
Capsule|4884,4891
-|4892,4893
1|4894,4895
Capsule|4896,4903
(|4903,4904
s|4904,4905
)|4905,4906
by|4907,4909
mouth|4910,4915
three|4916,4921
times|4922,4927
<EOL>|4928,4929
<EOL>|4930,4931
a|4931,4932
day|4933,4936
<EOL>|4938,4939
CALCITRIOL|4939,4949
-|4950,4951
0.25|4952,4956
mcg|4957,4960
Capsule|4961,4968
-|4969,4970
1|4971,4972
Capsule|4973,4980
(|4980,4981
s|4981,4982
)|4982,4983
by|4984,4986
mouth|4987,4992
every|4993,4998
<EOL>|4999,5000
other|5000,5005
<EOL>|5007,5008
day|5008,5011
<EOL>|5013,5014
CITALOPRAM|5014,5024
-|5025,5026
(|5027,5028
Prescribed|5028,5038
by|5039,5041
Other|5042,5047
Provider|5048,5056
)|5056,5057
-|5058,5059
10|5060,5062
mg|5063,5065
Tablet|5066,5072
-|5073,5074
1|5075,5076
<EOL>|5078,5079
Tablet|5079,5085
(|5085,5086
s|5086,5087
)|5087,5088
by|5089,5091
mouth|5092,5097
once|5098,5102
a|5103,5104
day|5105,5108
<EOL>|5110,5111
CLOPIDOGREL|5111,5122
[|5123,5124
PLAVIX|5124,5130
]|5130,5131
-|5132,5133
(|5134,5135
Prescribed|5135,5145
by|5146,5148
Other|5149,5154
Provider|5155,5163
)|5163,5164
-|5165,5166
75|5167,5169
mg|5170,5172
<EOL>|5174,5175
Tablet|5175,5181
-|5182,5183
1|5184,5185
Tablet|5186,5192
(|5192,5193
s|5193,5194
)|5194,5195
by|5196,5198
mouth|5199,5204
once|5205,5209
a|5210,5211
day|5212,5215
<EOL>|5217,5218
FOLIC|5218,5223
ACID|5224,5228
-|5229,5230
1|5231,5232
mg|5233,5235
Tablet|5236,5242
-|5243,5244
one|5245,5248
Tablet|5249,5255
(|5255,5256
s|5256,5257
)|5257,5258
by|5259,5261
mouth|5262,5267
one|5268,5271
daily|5272,5277
-|5278,5279
No|5280,5282
<EOL>|5283,5284
<EOL>|5285,5286
Substitution|5286,5298
<EOL>|5300,5301
LORAZEPAM|5301,5310
-|5311,5312
0.5|5313,5316
mg|5317,5319
Tablet|5320,5326
-|5327,5328
_|5329,5330
_|5330,5331
_|5331,5332
Tablet|5333,5339
(|5339,5340
s|5340,5341
)|5341,5342
by|5343,5345
mouth|5346,5351
q6|5352,5354
hours|5355,5360
as|5361,5363
<EOL>|5365,5366
needed|5366,5372
for|5373,5376
Nausea|5377,5383
<EOL>|5385,5386
METOPROLOL|5386,5396
TARTRATE|5397,5405
[|5406,5407
LOPRESSOR|5407,5416
]|5416,5417
-|5418,5419
(|5420,5421
Prescribed|5421,5431
by|5432,5434
Other|5435,5440
Provider|5441,5449
)|5449,5450
<EOL>|5451,5452
<EOL>|5453,5454
-|5454,5455
50|5456,5458
mg|5459,5461
Tablet|5462,5468
-|5469,5470
one|5471,5474
Tablet|5475,5481
(|5481,5482
s|5482,5483
)|5483,5484
by|5485,5487
mouth|5488,5493
_|5494,5495
_|5495,5496
_|5496,5497
BID|5498,5501
-|5502,5503
No|5504,5506
<EOL>|5507,5508
Substitution|5508,5520
<EOL>|5522,5523
TRAMADOL|5523,5531
-|5532,5533
(|5534,5535
Prescribed|5535,5545
by|5546,5548
Other|5549,5554
Provider|5555,5563
)|5563,5564
-|5565,5566
50|5567,5569
mg|5570,5572
Tablet|5573,5579
-|5580,5581
0.5|5582,5585
<EOL>|5587,5588
(|5588,5589
One|5589,5592
half|5593,5597
)|5597,5598
Tablet|5599,5605
(|5605,5606
s|5606,5607
)|5607,5608
by|5609,5611
mouth|5612,5617
three|5618,5623
times|5624,5629
a|5630,5631
day|5632,5635
as|5636,5638
needed|5639,5645
for|5646,5649
<EOL>|5651,5652
Pain|5652,5656
<EOL>|5658,5659
TRAZODONE|5659,5668
-|5669,5670
50|5671,5673
mg|5674,5676
Tablet|5677,5683
-|5684,5685
one|5686,5689
Tablet|5690,5696
(|5696,5697
s|5697,5698
)|5698,5699
by|5700,5702
mouth|5703,5708
one|5709,5712
daily|5713,5718
as|5719,5721
<EOL>|5723,5724
needed|5724,5730
-|5731,5732
No|5733,5735
Substitution|5736,5748
<EOL>|5750,5751
ASPIRIN|5751,5758
-|5759,5760
(|5761,5762
Prescribed|5762,5772
by|5773,5775
Other|5776,5781
Provider|5782,5790
:|5790,5791
_|5792,5793
_|5793,5794
_|5794,5795
.|5795,5796
)|5796,5797
-|5798,5799
81|5800,5802
<EOL>|5803,5804
<EOL>|5805,5806
mg|5806,5808
Tablet|5809,5815
,|5815,5816
Chewable|5817,5825
-|5826,5827
1|5828,5829
Tablet|5830,5836
(|5836,5837
s|5837,5838
)|5838,5839
by|5840,5842
mouth|5843,5848
one|5849,5852
daily|5853,5858
-|5859,5860
No|5861,5863
<EOL>|5865,5866
Substitution|5866,5878
<EOL>|5880,5881
RANITIDINE|5881,5891
HCL|5892,5895
[|5896,5897
ACID|5897,5901
CONTROL|5902,5909
]|5909,5910
-|5911,5912
150|5913,5916
mg|5917,5919
Tablet|5920,5926
-|5927,5928
one|5929,5932
Tablet|5933,5939
(|5939,5940
s|5940,5941
)|5941,5942
by|5943,5945
<EOL>|5946,5947
<EOL>|5948,5949
mouth|5949,5954
one|5955,5958
daily|5959,5964
-|5965,5966
No|5967,5969
Substitution|5970,5982
<EOL>|5984,5985
<EOL>|5986,5987
Discharge|5987,5996
Medications|5997,6008
:|6008,6009
<EOL>|6009,6010
N|6010,6011
/|6011,6012
A|6012,6013
<EOL>|6013,6014
<EOL>|6015,6016
Discharge|6016,6025
Disposition|6026,6037
:|6037,6038
<EOL>|6038,6039
Expired|6039,6046
<EOL>|6046,6047
<EOL>|6048,6049
Discharge|6049,6058
Diagnosis|6059,6068
:|6068,6069
<EOL>|6069,6070
1.|6070,6072
Non|6073,6076
small|6077,6082
cell|6083,6087
lung|6088,6092
cancer|6093,6099
<EOL>|6099,6100
2.|6100,6102
Melena|6103,6109
<EOL>|6109,6110
<EOL>|6111,6112
Discharge|6112,6121
Condition|6122,6131
:|6131,6132
<EOL>|6132,6133
Expired|6133,6140
<EOL>|6140,6141
<EOL>|6142,6143
Discharge|6143,6152
Instructions|6153,6165
:|6165,6166
<EOL>|6166,6167
N|6167,6168
/|6168,6169
A|6169,6170
<EOL>|6170,6171
<EOL>|6172,6173
Followup|6173,6181
Instructions|6182,6194
:|6194,6195
<EOL>|6195,6196
_|6196,6197
_|6197,6198
_|6198,6199
<EOL>|6199,6200

