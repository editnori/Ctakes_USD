CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Role Class - access|Finding|false|false||accessnull|Access|Modifier|false|false||accessnull|Intra-Aortic Balloon Pumping|Procedure|false|false||IABPnull|null|Device|false|false||IABPnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Hypertensive disease|Disorder|false|false||HTNnull|null|Time|false|false||priornull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Catheterization|Procedure|false|false||cathnull|Catheterization|Procedure|false|false||catheterizationnull|Concern|Finding|false|false||concernnull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Angina Pectoris|Finding|false|false||angina painnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Exertion|Finding|false|false||exertionnull|Night time|Time|false|false||nightnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||acute onsetnull|Sudden onset (attribute)|Time|false|false||acute onset
null|acute|Time|false|false||acute onsetnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Morning|Time|false|false||morningnull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Episode of|Time|false|false||episodesnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Malaise|Finding|false|false||malaisenull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Palpitations|Finding|false|false||palpitationsnull|Dyspnea|Finding|false|false||SOBnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Chest Pain|Finding|false|false||Chest painnull|null|Attribute|false|false||Chest painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Laboratory test finding|Lab|false|false||Labsnull|Leukocytes|Anatomy|false|false||WBCnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|CR1 protein, human|Drug|false|false||Cr1
null|Complement 3b Receptor|Drug|false|false||Cr1
null|Complement 3b Receptor|Drug|false|false||Cr1
null|CR1 protein, human|Drug|false|false||Cr1null|CR1 protein, human|Finding|false|false||Cr1
null|Complement 3b Receptor|Finding|false|false||Cr1
null|CR1 gene|Finding|false|false||Cr1null|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Elevation|Modifier|false|false||elevationsnull|aVR|Modifier|false|false||AVRnull|Borderline|Modifier|false|false||borderlinenull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Diffuse|Modifier|false|false||diffusenull|Mental Depression|Disorder|false|false||depressionsnull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Septal|Modifier|false|false||septalnull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|ticagrelor|Drug|false|false||Ticagrelor
null|ticagrelor|Drug|false|false||Ticagrelornull|vancomycin|Drug|false|false||Vanco
null|vancomycin|Drug|false|false||Vanconull|Cardiac Catheterization Procedures|Procedure|false|false||cardiac cathnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||cathnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Apyrexial|Finding|false|false||afebrilenull|Catheterization|Procedure|false|false||Cathnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Still|Disorder|false|false||stillnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Catheterization|Procedure|false|false||Catheterizationnull|Septal|Modifier|false|false||septalnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Diffuse|Modifier|false|false||diffusenull|Disease|Disorder|false|false||diseasenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Circumflex|Modifier|false|false||circumflexnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Main|Modifier|false|false||main
null|Primary|Modifier|false|false||mainnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Role Class - access|Finding|false|false||accessnull|Access|Modifier|false|false||accessnull|Hypotensive|Finding|false|false||Hypotensivenull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false||IVFnull|SCN5A wt Allele|Finding|false|false||IVF
null|SCN5A gene|Finding|false|false||IVFnull|Assisted Reproductive Technologies|Procedure|false|false||IVF
null|Fertilization in Vitro|Procedure|false|false||IVFnull|Structure of interventricular foramen|Anatomy|false|false||IVFnull|Coughing|Finding|false|false||Coughingnull|Post-Procedure|Time|false|false||post-procedurenull|Left ventricular end-diastolic pressure|Finding|false|false||LVEDPnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Hypertensive (finding)|Finding|false|false||hypertensivenull|Further|Modifier|false|false||furthernull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Coronary Care Units|Device|false|false||CCUnull|Coronary Care Units|Entity|false|false||CCUnull|Hypotension|Finding|false|false||hypotensionnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Leukocytes|Anatomy|false|false||WBCnull|Lacking|Modifier|false|false||lacknull|Beds|Device|false|false||bedsnull|Coronary Care Units|Device|false|false||CCUnull|Coronary Care Units|Entity|false|false||CCUnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Productive Cough|Finding|false|false||productive coughnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Two weeks|Time|false|false||two weeksnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|Current (present time)|Time|false|false||Currentlynull|clarithromycin|Drug|false|false||clarithromycin
null|clarithromycin|Drug|false|false||clarithromycinnull|amoxicillin|Drug|false|false||amoxicillin
null|amoxicillin|Drug|false|false||amoxicillinnull|Night time|Time|false|false||nightnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Weight Loss|Finding|false|false||weight loss
null|Losing Weight (question)|Finding|false|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|false|false||weight lossnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|month|Time|false|false||monthsnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||HTNnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Management procedure|Event|false|false||managednull|Spinal canal stenosis|Disorder|false|false||Spinal stenosis
null|Spinal Stenosis|Disorder|false|false||Spinal stenosisnull|Spinal|Modifier|false|false||Spinalnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Cardiomyopathies|Disorder|false|false||cardiomyopathynull|Family Medical History|Finding|true|false||family history ofnull|Family Medical History|Finding|true|false||family historynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|true|true||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Early|Time|false|false||earlynull|Cardiac Arrhythmia|Disorder|true|false||arrhythmianull|Sudden (qualifier value)|Modifier|false|false||suddennull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Event Consequence - Death|Finding|false|false||death
null|Death (finding)|Finding|false|false||death
null|Cessation of life|Finding|false|false||deathnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Apyrexial|Finding|false|false||afebrilenull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|Telephone Number|Finding|false|false||Tele
null|TCAP gene|Finding|false|false||Telenull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Slightly (qualifier value)|Modifier|false|false||Slightly
null|Slight (qualifier value)|Modifier|false|false||Slightlynull|Tachypnea|Finding|false|false||tachypneicnull|Male population group|Subject|false|false||man
null|Homo sapiens|Subject|false|false||man
null|Males|Subject|false|false||mannull|Mandinka Language|Entity|false|false||mannull|Wheezing|Finding|false|false||wheezingnull|Sentence|Finding|false|false||sentencesnull|HEENT|Anatomy|false|false||HEENTnull|PERRLA|Finding|false|false||PERRLAnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Jugular venous engorgement|Finding|true|false||JVDnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Heart Sounds|Finding|false|false||heart soundsnull|auscultation of heart sounds|Procedure|false|false||heart soundsnull|null|Attribute|false|false||heart soundsnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Rhonchi|Finding|false|false||rhonchinull|Lung|Anatomy|false|false||LUNGSnull|Rhonchi|Finding|false|false||rhonchinull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Expiratory wheezing|Finding|false|false||expiratory wheezingnull|Expiration, Respiratory|Finding|false|false||expiratorynull|Wheezing|Finding|false|false||wheezingnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Right arm|Anatomy|false|false||R armnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Bands|Device|false|false||bandnull|Band form|Modifier|false|false||bandnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Sensory perception|Finding|false|false||sensory functionnull|Sensory (qualifier value)|Modifier|false|false||sensorynull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Full|Modifier|false|false||fullnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Rupture of Membranes|Finding|false|false||ROM
null|ROM1 gene|Finding|false|false||ROMnull|Range of motion technique (procedure)|Procedure|false|false||ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Chronic - Admission Level of Care Code|Finding|true|false||chronicnull|Provision of recurring care for chronic illness|Procedure|true|false||chronicnull|chronic|Time|false|false||chronicnull|Edema|Finding|false|false||edematousnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|At discharge|Time|false|false||At dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|HEENT|Anatomy|false|false||HEENTnull|PERRLA|Finding|false|false||PERRLAnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Jugular venous engorgement|Finding|true|false||JVDnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Heart Sounds|Finding|false|false||heart soundsnull|auscultation of heart sounds|Procedure|false|false||heart soundsnull|null|Attribute|false|false||heart soundsnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Lung|Anatomy|false|false||LUNGSnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Right arm|Anatomy|false|false||R armnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Sensory perception|Finding|false|false||sensory functionnull|Sensory (qualifier value)|Modifier|false|false||sensorynull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Full|Modifier|false|false||fullnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Rupture of Membranes|Finding|false|false||ROM
null|ROM1 gene|Finding|false|false||ROMnull|Range of motion technique (procedure)|Procedure|false|false||ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Chronic - Admission Level of Care Code|Finding|true|false||chronicnull|Provision of recurring care for chronic illness|Procedure|true|false||chronicnull|chronic|Time|false|false||chronicnull|Edema|Finding|false|false||edematousnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Laboratory test finding|Lab|false|false||Labsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Mandibular left lateral incisor mesial prosthesis|Device|false|false||23PMnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Megakaryocyte-Potentiating Factor, human|Drug|false|false||SMR
null|Megakaryocyte-Potentiating Factor, human|Drug|false|false||SMRnull|MSLN wt Allele|Finding|false|false||SMR
null|MSLN gene|Finding|false|false||SMRnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Bands|Device|false|false||BANDSnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Mandibular left lateral incisor mesial prosthesis|Device|false|false||23PMnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular left lateral incisor mesial prosthesis|Device|false|false||23PMnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|calcium|Drug|false|false||CALCIUM
null|CALCIUM SUPPLEMENTS|Drug|false|false||CALCIUM
null|Calcium, Dietary|Drug|false|false||CALCIUM
null|Calcium [EPC]|Drug|false|false||CALCIUM
null|Calcium Drug Class|Drug|false|false||CALCIUMnull|Calcium metabolic function|Finding|false|false||CALCIUMnull|Calcium measurement|Procedure|false|false||CALCIUMnull|phosphate ion|Drug|false|false||PHOSPHATE
null|Phosphates|Drug|false|false||PHOSPHATE
null|phosphate ion|Drug|false|false||PHOSPHATEnull|Phosphate measurement|Procedure|false|false||PHOSPHATEnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|magnesium|Drug|false|false||MAGNESIUM
null|Magnesium Drug Class|Drug|false|false||MAGNESIUM
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||MAGNESIUMnull|Magnesium measurement|Procedure|false|false||MAGNESIUMnull|Glycosylated hemoglobin A|Drug|false|false||HbA1c
null|Glycosylated hemoglobin A|Drug|false|false||HbA1cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1cnull|KCNH1 gene|Finding|false|false||eAGnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Mandibular left lateral incisor mesial prosthesis|Device|false|false||23PMnull|High Density Lipoproteins|Drug|false|false||HDL
null|High Density Lipoproteins|Drug|false|false||HDLnull|HSD11B1 wt Allele|Finding|false|false||HDLnull|High density lipoprotein measurement|Procedure|false|false||HDLnull|High Density Lipoproteins|Drug|false|false||HDL
null|High Density Lipoproteins|Drug|false|false||HDLnull|HSD11B1 wt Allele|Finding|false|false||HDLnull|High density lipoprotein measurement|Procedure|false|false||HDLnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|MICU1 gene|Finding|false|false||CALCnull|Intracalcarine cortex|Anatomy|false|false||CALCnull|Mandibular left lateral incisor mesial prosthesis|Device|false|false||23PMnull|Bur - medical device|Device|false|false||BURRnull|Burr - plant|Entity|false|false||BURRnull|Laboratory test finding|Lab|false|false||Labsnull|At discharge|Time|false|false||at Dischargenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bands|Device|false|false||Bandsnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Relevance|Modifier|false|false||Relevantnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Left atrial structure|Anatomy|false|false||left atriumnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false||atriumnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Heart Atrium|Anatomy|false|false||atrialnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mmHgnull|Wall of left ventricle|Anatomy|false|false||Left ventricular wallnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Wall of ventricle|Anatomy|false|false||ventricular wallnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Overall Publication Type|Finding|false|false||Overallnull|Overall|Modifier|false|false||Overallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Moderate Response|Finding|false|false||moderately
null|Moderate|Finding|false|false||moderately
null|Moderate Effect|Finding|false|false||moderatelynull|Moderate (severity modifier)|Modifier|false|false||moderately
null|Moderation|Modifier|false|false||moderatelynull|Depressed mood|Disorder|false|false||depressednull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Knowledge acquisition using a method of assessment|Finding|false|false||assessmentnull|assessment of cognitive functions|Procedure|false|false||assessment
null|Physical Examination|Procedure|false|false||assessment
null|Nutrition Assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Personal care assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Evaluation procedure|Procedure|false|false||assessment
null|Evaluation|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessmentnull|Assessed|Event|false|false||assessmentnull|Suboptimal Image Reason|Finding|false|false||suboptimal imagenull|Suboptimal|Modifier|false|false||suboptimalnull|Image Quality|Modifier|false|false||image qualitynull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false||imagenull|Image (foundation metadata concept)|Finding|false|false||image
null|Image|Finding|false|false||image
null|Medical Image|Finding|false|false||image
null|image - dosage form|Finding|false|false||imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Quality|Modifier|false|false||qualitynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Variability|Finding|false|false||variabilitynull|Hypokinesia|Finding|false|false||hypokinesisnull|APEX1 protein, human|Drug|false|false||apex
null|APEX1 protein, human|Drug|false|false||apexnull|APEX1 gene|Finding|false|false||apexnull|dinoflagellate apex|Anatomy|false|false||apexnull|Highest|Modifier|false|false||apexnull|Ventricular Septal Defects|Disorder|true|false||ventricular septal defectnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Congenital septal defect of heart|Disorder|true|false||septal defect
null|Heart Septal Defects|Disorder|true|false||septal defectnull|Septal|Modifier|false|false||septalnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|true|false||defectnull|Defect|Finding|true|false||defectnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Ascending aorta structure|Anatomy|false|false||ascending aortanull|Sequencing - Ascending|Finding|false|false||ascending
null|Ascend (action)|Finding|false|false||ascendingnull|Ascending|Modifier|false|false||ascendingnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Valve Area|Finding|false|false||valve areanull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Chiari malformation type II|Disorder|false|false||cm2null|sq. cm|LabModifier|false|false||cm2null|Aortic Valve Insufficiency|Disorder|true|false||aortic regurgitationnull|Aorta|Anatomy|false|false||aorticnull|Regurgitation|Finding|true|false||regurgitation
null|Regurgitates after swallowing|Finding|true|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|true|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Pulmonary artery systolic pressure|Finding|false|false||pulmonary artery systolic pressurenull|Pulmonary artery structure|Anatomy|false|false||pulmonary arterynull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Systolic Pressure|Attribute|false|false||systolic pressurenull|Systole|Finding|false|false||systolicnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Physiological|Finding|false|false||physiologicnull|Pericardial effusion|Disorder|false|false||pericardial effusionnull|Pericardial effusion body substance|Finding|false|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|null|Time|false|false||priornull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Probably|Finding|false|false||probably
null|Probable diagnosis|Finding|false|false||probablynull|Similarity|Modifier|false|false||similarnull|Suboptimal Image Reason|Finding|false|false||suboptimal imagenull|Suboptimal|Modifier|false|false||suboptimalnull|Image Quality|Modifier|false|false||image qualitynull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false||imagenull|Image (foundation metadata concept)|Finding|false|false||image
null|Image|Finding|false|false||image
null|Medical Image|Finding|false|false||image
null|image - dosage form|Finding|false|false||imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Quality|Modifier|false|false||qualitynull|Scientific Study|Procedure|false|false||studiesnull|Definite|Modifier|false|false||definite
null|Definitely Related to Intervention|Modifier|false|false||definitenull|Comparison|Event|false|false||comparisonnull|Plain chest X-ray|Procedure|false|false||CXRnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Generalized|Modifier|false|false||Generalizednull|Improvement|Finding|false|false||improvementnull|Bilateral lungs|Anatomy|false|false||both lungsnull|Lung|Anatomy|false|false||lungsnull|Probably|Finding|false|false||probably
null|Probable diagnosis|Finding|false|false||probablynull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Still|Disorder|false|false||stillnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Structure of right upper lobe of lung|Anatomy|false|false||right upper lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of upper lobe of lung|Anatomy|false|false||upper lobenull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Probably|Finding|false|false||probably
null|Probable diagnosis|Finding|false|false||probablynull|Pneumonia|Disorder|false|false||pneumonianull|Bilateral|Modifier|false|false||bilateralnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Component object|Device|false|false||componentsnull|heart size|Finding|false|false||Heart sizenull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Micro (prefix)|Finding|false|false||MICRO
null|Microbiology - Laboratory Class|Finding|false|false||MICROnull|Microbiology procedure|Procedure|false|false||MICROnull|Unit Of Measure Prefix - micro|LabModifier|false|false||MICROnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|dna amplification|Finding|false|false||DNA amplificationnull|DNA|Drug|false|false||DNA
null|DNA|Drug|false|false||DNAnull|Gene Amplification Abnormality|Disorder|false|false||amplificationnull|Gene Amplification Technique|Procedure|false|false||amplificationnull|Amplification|Phenomenon|false|false||amplificationnull|Biological Assay|Procedure|false|false||assay
null|Assay|Procedure|false|false||assaynull|assay qualifier|Modifier|false|false||assaynull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Clostridioides difficile|Entity|false|false||CLOSTRIDIUM DIFFICILEnull|Genus Clostridium (organism)|Entity|false|false||CLOSTRIDIUMnull|Positive|Finding|false|false||Positive fornull|BRAF Gene Rearrangement|Disorder|false|false||Positivenull|Rh Positive Blood Group|Finding|false|false||Positive
null|Positive Finding|Finding|false|false||Positive
null|Positive|Finding|false|false||Positivenull|Positive Charge|Modifier|false|false||Positivenull|Positive Number|LabModifier|false|false||Positivenull|Toxigenic|Finding|false|false||toxigenicnull|DNA|Drug|false|false||DNA
null|DNA|Drug|false|false||DNAnull|Gene Amplification Abnormality|Disorder|false|false||amplificationnull|Gene Amplification Technique|Procedure|false|false||amplificationnull|Amplification|Phenomenon|false|false||amplificationnull|Reference range (qualifier value)|Modifier|false|false||Reference Rangenull|null|LabModifier|false|false||Reference Rangenull|Reference - MdfHmdMetSourceType|Finding|false|false||Reference
null|Reference Object|Finding|false|false||Reference
null|Reference source|Finding|false|false||Reference
null|Bibliographic Reference|Finding|false|false||Reference
null|Reference - HL7UpdateMode|Finding|false|false||Referencenull|Concept model range (foundation metadata concept)|Finding|false|false||Rangenull|Sample Range|LabModifier|false|false||Range
null|Range|LabModifier|false|false||Rangenull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Specimen Type - Sputum|Finding|false|false||SPUTUM
null|null|Finding|false|false||SPUTUM
null|Sputum|Finding|false|false||SPUTUMnull|Source (property) (qualifier value)|Finding|false|false||Source
null|Term Source|Finding|false|false||Source
null|Source|Finding|false|false||Sourcenull|Does expectorate|Finding|false|false||Expectoratednull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Epithelial Cells|Anatomy|false|false||epithelial cellsnull|Epithelial|Modifier|false|false||epithelialnull|Cells|Anatomy|false|false||cellsnull|Per 100x Field|LabModifier|false|false||/100X fieldnull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|Knowledge Field|Finding|true|false||FIELD
null|Force Field|Finding|true|false||FIELD
null|Field|Finding|true|false||FIELDnull|field - patient encounter|Procedure|true|false||FIELDnull|Gram-negative bacillus|Entity|false|false||GRAM NEGATIVE RODnull|gram|LabModifier|false|false||GRAMnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Renal Osteodystrophy|Disorder|true|false||RODnull|KNTC1 gene|Finding|true|false||RODnull|Rod Photoreceptors|Anatomy|false|false||RODnull|Rod Device|Device|true|false||RODnull|Form-bacillus|Entity|true|false||RODnull|Rod Shape|Modifier|false|false||RODnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Saccharomycetales|Entity|false|false||BUDDING YEASTnull|Cell budding|Finding|false|false||BUDDINGnull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|Quality|Modifier|false|false||QUALITYnull|Specimen|Drug|false|false||SPECIMENnull|Role Class - specimen|Finding|false|false||SPECIMEN
null|Biospecimen|Finding|false|false||SPECIMENnull|Respiratory culture|Procedure|false|false||RESPIRATORY CULTUREnull|Respiratory attachment|Finding|false|false||RESPIRATORY
null|respiratory|Finding|false|false||RESPIRATORY
null|null|Finding|false|false||RESPIRATORY
null|Respiratory specimen|Finding|false|false||RESPIRATORYnull|Respiratory rate|Attribute|false|false||RESPIRATORYnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Further|Modifier|false|false||Furthernull|Incubation|Procedure|false|false||incubationnull|Providing presence (regime/therapy)|Procedure|false|false||presencenull|Presence (property)|Modifier|false|false||presencenull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Symbiotic|Finding|false|false||commensalnull|Commensal parasite|Entity|false|false||commensalnull|Pharyngeal/Respiratory Flora|Entity|false|false||respiratory floranull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|Disorder|false|false||KLEBSIELLA PNEUMONIAEnull|Klebsiella pneumoniae|Entity|false|false||KLEBSIELLA PNEUMONIAEnull|Pneumonia due to Klebsiella pneumoniae|Disorder|false|false||KLEBSIELLAnull|Klebsiella|Entity|false|false||KLEBSIELLAnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|cefazolin|Drug|false|false||Cefazolin
null|cefazolin|Drug|false|false||Cefazolinnull|criteria|Finding|false|false||criterianull|Dosage|LabModifier|false|false||dosagenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Gram-negative bacillus|Entity|false|false||GRAM NEGATIVE RODnull|gram|LabModifier|false|false||GRAMnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Renal Osteodystrophy|Disorder|false|false||RODnull|KNTC1 gene|Finding|false|false||RODnull|Rod Photoreceptors|Anatomy|false|false||RODnull|Rod Device|Device|false|false||RODnull|Form-bacillus|Entity|false|false||RODnull|Rod Shape|Modifier|false|false||RODnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|Disorder|false|false||KLEBSIELLA PNEUMONIAEnull|Klebsiella pneumoniae|Entity|false|false||KLEBSIELLA PNEUMONIAEnull|Pneumonia due to Klebsiella pneumoniae|Disorder|false|false||KLEBSIELLAnull|Klebsiella|Entity|false|false||KLEBSIELLAnull|Ampicillin / Sulbactam|Drug|false|false||AMPICILLIN/SULBACTAMnull|ampicillin|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillin|Drug|false|false||AMPICILLINnull|sulbactam|Drug|false|false||SULBACTAM
null|sulbactam|Drug|false|false||SULBACTAMnull|cefazolin|Drug|false|false||CEFAZOLIN
null|cefazolin|Drug|false|false||CEFAZOLINnull|cefepime|Drug|false|false||CEFEPIME
null|cefepime|Drug|false|false||CEFEPIMEnull|ceftazidime|Drug|false|false||CEFTAZIDIME
null|ceftazidime|Drug|false|false||CEFTAZIDIMEnull|ceftriaxone|Drug|false|false||CEFTRIAXONE
null|ceftriaxone|Drug|false|false||CEFTRIAXONEnull|ciprofloxacin|Drug|false|false||CIPROFLOXACIN
null|ciprofloxacin|Drug|false|false||CIPROFLOXACINnull|gentamicin|Drug|false|false||GENTAMICIN
null|gentamicin|Drug|false|false||GENTAMICINnull|Gentamicin measurement|Procedure|false|false||GENTAMICINnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEMnull|piperacillin|Drug|false|false||PIPERACILLIN
null|piperacillin|Drug|false|false||PIPERACILLINnull|tazobactam|Drug|false|false||TAZO
null|tazobactam|Drug|false|false||TAZOnull|tobramycin|Drug|false|false||TOBRAMYCIN
null|tobramycin|Drug|false|false||TOBRAMYCINnull|Tobramycin measurement|Procedure|false|false||TOBRAMYCINnull|trimethoprim|Drug|false|false||TRIMETHOPRIM
null|trimethoprim|Drug|false|false||TRIMETHOPRIMnull|sulfa|Drug|false|false||SULFAnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Hypertensive disease|Disorder|false|false||HTNnull|Old|Time|false|false||oldnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Diffuse|Modifier|false|false||diffusenull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|SULT1E1 wt Allele|Finding|false|false||STE
null|SULT1E1 gene|Finding|false|false||STEnull|aVR|Modifier|false|false||aVRnull|Mental Depression|Disorder|false|false||depressionsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Numerous|LabModifier|false|false||multinull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Catheterization|Procedure|false|false||cathnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|ACE protein, human|Drug|false|false||ACE
null|ACE protein, human|Drug|false|false||ACEnull|ACE gene|Finding|false|false||ACE
null|Adverse Childhood Experience questionnaire|Finding|false|false||ACEnull|cisplatin, cytarabine, and etoposide chemotherapy protocol|Procedure|false|false||ACE
null|cyclophosphamide/doxorubicin protocol|Procedure|false|false||ACE
null|CDE protocol|Procedure|false|false||ACE
null|CDE Regimen|Procedure|false|false||ACEnull|Achinese language|Entity|false|false||ACEnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|ECHO protocol|Procedure|false|false||Echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||Echonull|Echo <Calopterygidae>|Entity|false|false||Echonull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Hypokinesia|Finding|false|false||hypokinesisnull|APEX1 protein, human|Drug|false|false||apex
null|APEX1 protein, human|Drug|false|false||apexnull|APEX1 gene|Finding|false|false||apexnull|dinoflagellate apex|Anatomy|false|false||apexnull|Highest|Modifier|false|false||apexnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Hypokinesia|Finding|false|false||hypokineticnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Atrial Fibrillation|Disorder|false|false||atrial fibrillationnull|null|Attribute|false|false||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Possible|Finding|false|false||Possiblynull|Possible diagnosis|Modifier|false|false||Possiblynull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Pulmonary Wedge Pressure|Attribute|false|false||PCWPnull|Initially|Time|false|false||initiallynull|Pressors|Drug|false|false||pressorsnull|Balloon Dilatation|Procedure|false|false||balloonnull|Medical Balloon Device|Device|false|false||balloon
null|Balloon Device|Device|false|false||balloon
null|Balloon Aircraft|Device|false|false||balloonnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Atrial Fibrillation|Disorder|false|false||Atrial Fibrillationnull|null|Attribute|false|false||Atrial Fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Atrial Fibrillationnull|Heart Atrium|Anatomy|false|false||Atrialnull|Fibrillation|Disorder|false|false||Fibrillationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Paroxysmal|Time|false|false||paroxysmalnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|digoxin|Drug|false|false||digoxin
null|digoxin|Drug|false|false||digoxinnull|Digoxin measurement|Procedure|false|false||digoxinnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Daily|Time|false|false||dailynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|During admission|Time|false|false||during admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Decision|Finding|false|false||decisionnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|digoxin|Drug|false|false||digoxin
null|digoxin|Drug|false|false||digoxinnull|Digoxin measurement|Procedure|false|false||digoxinnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Hematuria|Disorder|false|false||Hematurianull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Traumatic|Finding|false|false||traumaticnull|Systemic Route of Administration|Finding|false|false||systemic
null|Systemic|Finding|false|false||systemicnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cytology--Technique|Procedure|false|false||Cytology
null|Cytological Techniques|Procedure|false|false||Cytologynull|Cytology|Title|false|false||Cytologynull|cellular aspects|Modifier|false|false||Cytologynull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Urology|Title|false|false||urologynull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Episode of|Time|false|false||episodesnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Improved - answer to question|Finding|false|false||improved
null|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Plain chest X-ray|Procedure|false|false||CXRnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Structure of right upper lobe of lung|Anatomy|false|false||RULnull|Aspiration Pneumonia|Disorder|false|false||aspiration pneumonia
null|Aspiration pneumonitis|Disorder|false|false||aspiration pneumonianull|Respiratory Aspiration|Disorder|false|false||aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Pneumonia|Disorder|false|false||pneumonianull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Focal|Modifier|false|false||focalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Peptide Nucleic Acids|Drug|false|false||pnanull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Culture (Anthropological)|Finding|false|false||culturesnull|Pneumonia due to Klebsiella pneumoniae|Disorder|false|false||Klebsiella pneumonianull|Pneumonia due to Klebsiella pneumoniae|Disorder|false|false||Klebsiellanull|Klebsiella|Entity|false|false||Klebsiellanull|Pneumonia|Disorder|false|false||pneumonianull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Biomaterial Treatment|Finding|true|false||treatment
null|Treating|Finding|true|false||treatment
null|therapeutic aspects|Finding|true|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|true|false||treatment
null|Administration (procedure)|Procedure|true|false||treatment
null|Therapeutic procedure|Procedure|true|false||treatmentnull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Daily|Time|false|false||dailynull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Electrolytes|Drug|false|false||electrolytes
null|Electrolytes|Drug|false|false||electrolytes
null|Electrolyte [EPC]|Drug|false|false||electrolytesnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Loose stool|Finding|false|false||loose stoolnull|Loose|Modifier|false|false||loosenull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Antibiotics|Drug|false|false||antibioticnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Leukocytes|Anatomy|false|false||WBCnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Four times daily|Time|false|false||qidnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Gastroesophageal reflux disease|Disorder|false|false||GASTROESOPHAGEAL REFLUX DISEASE (GERD)null|Gastroesophageal reflux disease|Disorder|false|false||GASTROESOPHAGEAL REFLUX DISEASEnull|Gastroesophageal reflux disease|Disorder|false|false||GASTROESOPHAGEAL REFLUXnull|Infantile Gastroesophageal Reflux|Finding|false|false||GASTROESOPHAGEAL REFLUX
null|Acid reflux|Finding|false|false||GASTROESOPHAGEAL REFLUXnull|gastroesophageal|Anatomy|false|false||GASTROESOPHAGEALnull|Reflux|Finding|false|false||REFLUXnull|Disease|Disorder|false|false||DISEASEnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Endoscopy, Gastrointestinal|Procedure|false|false||Endoscopy
null|Endoscopy (procedure)|Procedure|false|false||Endoscopynull|Helicobacter pylori|Entity|false|false||H Pylorinull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|clarithromycin|Drug|false|false||clarithromycin
null|clarithromycin|Drug|false|false||clarithromycinnull|amoxicillin|Drug|false|false||amoxicillin
null|amoxicillin|Drug|false|false||amoxicillinnull|14 days|Time|false|false||14 daysnull|day|Time|false|false||daysnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Clostridium difficile infection|Disorder|false|false||c.diff infectionnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Delirium|Disorder|false|false||Deliriumnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Frequently|Time|false|false||frequentnull|Sundowning|Disorder|false|false||sundowningnull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|Seroquel|Drug|false|false||Seroquel
null|Seroquel|Drug|false|false||Seroquelnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Spinal canal stenosis|Disorder|false|false||Spinal Stenosis
null|Spinal Stenosis|Disorder|false|false||Spinal Stenosisnull|Spinal|Modifier|false|false||Spinalnull|Stenosis|Finding|false|false||Stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||Stenosisnull|Stenosis Morphology|Modifier|false|false||Stenosisnull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|cephradine|Drug|false|false||ced
null|cephradine|Drug|false|false||cednull|Camurati-Engelmann Syndrome|Disorder|false|false||ced
null|Cranioectodermal dysplasia|Disorder|false|false||cednull|Convection-Enhanced Delivery|Finding|false|false||ced
null|TGFB1 wt Allele|Finding|false|false||ced
null|TGFB1 gene|Finding|false|false||cednull|cisplatin/dexamethasone/etoposide protocol|Procedure|false|false||ced
null|CDE protocol|Procedure|false|false||cednull|naproxen|Drug|false|false||naproxen
null|naproxen|Drug|false|false||naproxennull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hospital course|Finding|true|false||hospital coursenull|null|Attribute|true|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|More|LabModifier|false|false||morenull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|false|false||NSAIDS
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDSnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Recent|Time|false|false||recentnull|ACSS2 protein, human|Drug|false|false||ACS
null|ACSS2 protein, human|Drug|false|false||ACSnull|Acrocallosal Syndrome|Disorder|false|false||ACS
null|Acute Chest Syndrome|Disorder|false|false||ACSnull|ACS - Activity Card Sort|Finding|false|false||ACS
null|American Community Survey|Finding|false|false||ACS
null|ACCS gene|Finding|false|false||ACS
null|CO-methylating acetyl-CoA synthase activity|Finding|false|false||ACS
null|PLA2G15 gene|Finding|false|false||ACS
null|ACSS2 wt Allele|Finding|false|false||ACS
null|ACSS2 gene|Finding|false|false||ACS
null|acetate-CoA ligase activity|Finding|false|false||ACSnull|anterior calcarine sulcus (human only)|Anatomy|false|false||ACSnull|Alternate Care Site|Device|false|false||ACSnull|American College of Surgeons|Entity|false|false||ACS
null|American Cancer Society|Entity|false|false||ACS
null|Alternate Care Site|Entity|false|false||ACSnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Arylsulfatase A, human|Drug|false|false||asa
null|Arylsulfatase A, human|Drug|false|false||asa
null|aspirin|Drug|false|false||asa
null|aspirin|Drug|false|false||asanull|ARSA gene|Finding|false|false||asanull|SHORT STATURE, IDIOPATHIC, X-LINKED|Disorder|false|false||ISSnull|During admission|Time|false|false||during admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|glipizide|Drug|false|false||glipizide
null|glipizide|Drug|false|false||glipizidenull|metformin|Drug|false|false||metformin
null|metformin|Drug|false|false||metforminnull|Hypertensive disease|Disorder|false|false||HTNnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|metoprolol dose|LabModifier|false|false||dose metoprololnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Urology|Title|false|false||urologynull|follow-up|Procedure|false|false||followupnull|Hematuria|Disorder|false|false||hematurianull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Urine cytology (finding)|Finding|false|false||Urine cytologynull|Urine cytology|Procedure|false|false||Urine cytologynull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Cytology--Technique|Procedure|false|false||cytology
null|Cytological Techniques|Procedure|false|false||cytologynull|Cytology|Title|false|false||cytologynull|cellular aspects|Modifier|false|false||cytologynull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Course|Time|false|false||coursenull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Electrolytes|Drug|false|false||electrolytes
null|Electrolytes|Drug|false|false||electrolytes
null|Electrolyte [EPC]|Drug|false|false||electrolytesnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Atrial Fibrillation|Disorder|false|false||atrial fibrillationnull|null|Attribute|false|false||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Daily|Time|false|false||dailynull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Recent|Time|false|false||recentnull|Stenting|Procedure|false|false||stent placementnull|null|Device|false|false||stentnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Daily|Time|false|false||dailynull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Daily|Time|false|false||dailynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|true|false||NSAIDS
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|true|false||NSAIDSnull|C4A wt Allele|Finding|false|false||SLP
null|C4A gene|Finding|false|false||SLPnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Pharyngeal structure|Anatomy|false|false||pharyngealnull|Muscular strength development exercise|Procedure|false|false||strengthening exercisesnull|Exercise|Finding|false|false||exercisesnull|Physical therapy exercises|Procedure|false|false||exercisesnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|naproxen|Drug|false|false||Naproxen
null|naproxen|Drug|false|false||Naproxennull|Daily|Time|false|false||DAILYnull|metformin|Drug|false|false||MetFORMIN
null|metformin|Drug|false|false||MetFORMINnull|Glucophage|Drug|false|false||Glucophage
null|Glucophage|Drug|false|false||Glucophagenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|glipizide|Drug|false|false||GlipiZIDE
null|glipizide|Drug|false|false||GlipiZIDEnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|digoxin|Drug|false|false||Digoxin
null|digoxin|Drug|false|false||Digoxinnull|Digoxin measurement|Procedure|false|false||Digoxinnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Aspirin EC|Drug|false|false||Aspirin EC
null|Aspirin EC|Drug|false|false||Aspirin ECnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|digoxin|Drug|false|false||Digoxin
null|digoxin|Drug|false|false||Digoxinnull|Digoxin measurement|Procedure|false|false||Digoxinnull|Daily|Time|false|false||DAILYnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|glipizide|Drug|false|false||GlipiZIDE
null|glipizide|Drug|false|false||GlipiZIDEnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|null|Drug|false|false||Vancomycin Oralnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Oral Liquid Product|Drug|false|false||Oral Liquidnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|Every six hours|Time|false|false||Q6Hnull|metformin|Drug|false|false||MetFORMIN
null|metformin|Drug|false|false||MetFORMINnull|Glucophage|Drug|false|false||Glucophage
null|Glucophage|Drug|false|false||Glucophagenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Mixed (Normal and Tumor)|Finding|false|false||mixed
null|Mixed (qualifier value)|Finding|false|false||mixednull|Hematuria|Disorder|false|false||Hematurianull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|TNF wt Allele|Finding|false|false||dif
null|TNF gene|Finding|false|false||difnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Delirium|Disorder|false|false||Deliriumnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Myocardial Infarction|Disorder|false|false||heart attacknull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Catheterization|Procedure|false|false||cathnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Partial Blockage within Medical Device|Finding|false|false||blockage
null|Blockage (obstruction - finding)|Finding|false|false||blockage
null|null|Finding|false|false||blockagenull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|null|Device|false|false||stentnull|Hypotension|Finding|false|false||low blood pressurenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Dysentery|Disorder|false|false||infectious diarrheanull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Physical trauma|Disorder|false|false||trauma
null|Traumatic injury|Disorder|false|false||trauma
null|Trauma|Disorder|false|false||traumanull|Trauma assessment and care|Procedure|false|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Anti-Inflammatory Agents|Drug|false|false||antiinflammatorynull|Pharmaceutical Preparations|Drug|false|false||drugsnull|Drugs - dental services|Procedure|false|false||drugsnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|false|false||NSAIDS
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDSnull|ibuprofen|Drug|false|false||ibuprofen
null|ibuprofen|Drug|false|false||ibuprofennull|Advil|Drug|false|false||advil
null|Advil|Drug|false|false||advilnull|AVIL gene|Finding|false|false||advilnull|Motrin|Drug|false|false||motrin
null|Motrin|Drug|false|false||motrinnull|Aleve|Drug|false|false||aleve
null|Aleve|Drug|false|false||alevenull|naproxen|Drug|false|false||naproxen
null|naproxen|Drug|false|false||naproxennull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Appointments|Event|false|false||appointmentsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions