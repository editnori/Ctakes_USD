 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|51,60|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|51,60|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|51,65|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|85,94|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|85,94|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|85,94|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|85,94|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|85,94|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|85,99|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|117,122|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|117,122|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|117,122|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|141,144|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|141,144|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|141,144|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|141,144|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|141,144|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|152,159|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|152,159|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|161,169|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|193,202|false|false|false|C1717415||Allergies
Event|Event|Allergies|193,202|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|193,202|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|205,227|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|213,217|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|213,217|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|213,227|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|218,227|false|false|false|||Reactions
Event|Event|Allergies|230,239|false|false|false|||Attending
Finding|Functional Concept|Allergies|230,239|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|265,270|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|Chief Complaint|265,276|false|false|false|C0733995|Structure of right flank|Right flank
Anatomy|Body Location or Region|Chief Complaint|271,276|false|false|false|C0230171|Flank (surface region)|flank
Disorder|Injury or Poisoning|Chief Complaint|277,285|false|false|false|C0009938|Contusions|bruising
Event|Event|Chief Complaint|277,285|false|false|false|||bruising
Finding|Finding|Chief Complaint|277,285|false|false|false|C2136686|reported bruising (history)|bruising
Attribute|Clinical Attribute|Chief Complaint|290,294|false|false|false|C2598155||pain
Event|Event|Chief Complaint|290,294|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|290,294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|290,294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Chief Complaint|299,303|false|false|false|C0085639|Falls|fall
Finding|Classification|Chief Complaint|306,311|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|312,320|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|312,320|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|324,342|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|333,342|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|333,342|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|333,342|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|333,342|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|333,342|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|History of Present Illness|402,409|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|402,409|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|402,412|false|false|false|C0262926|Medical History|history of
Finding|Conceptual Entity|History of Present Illness|413,419|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|History of Present Illness|413,419|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Intellectual Product|History of Present Illness|413,419|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Disorder|Disease or Syndrome|History of Present Illness|425,435|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|History of Present Illness|425,435|false|false|false|||deficiency
Finding|Functional Concept|History of Present Illness|425,435|false|false|false|C0011155|Deficiency|deficiency
Event|Event|History of Present Illness|441,449|false|false|false|||presents
Finding|Functional Concept|History of Present Illness|455,460|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|461,465|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|461,465|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|461,465|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|History of Present Illness|461,474|false|false|false|C0578454|Neck swelling|neck swelling
Event|Event|History of Present Illness|466,474|false|false|false|||swelling
Finding|Finding|History of Present Illness|466,474|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|466,474|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Daily or Recreational Activity|History of Present Illness|481,493|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Finding|Finding|History of Present Illness|481,493|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Event|Event|History of Present Illness|494,502|false|false|false|||accident
Event|Event|History of Present Illness|494,502|false|false|false|C1690974|Accidental event (event)|accident
Finding|Finding|History of Present Illness|494,502|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Finding|Idea or Concept|History of Present Illness|494,502|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Phenomenon|Phenomenon or Process|History of Present Illness|494,502|false|false|false|C0000924|Accidents|accident
Finding|Body Substance|History of Present Illness|509,516|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|509,516|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|509,516|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|517,524|false|false|false|||reports
Event|Event|History of Present Illness|533,537|false|false|false|||fell
Event|Event|History of Present Illness|544,556|false|false|false|||snowboarding
Event|Event|History of Present Illness|562,566|false|false|false|||loss
Finding|Finding|History of Present Illness|562,566|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|History of Present Illness|571,584|false|false|false|||consciousness
Finding|Finding|History of Present Illness|571,584|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|History of Present Illness|571,584|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Event|Event|History of Present Illness|610,614|false|false|false|||seen
Event|Event|History of Present Illness|632,639|false|false|false|||imaging
Finding|Finding|History of Present Illness|632,639|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|History of Present Illness|632,639|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Procedure|Diagnostic Procedure|History of Present Illness|632,647|false|false|false|C2711858|Imaging of head|imaging of head
Anatomy|Body Location or Region|History of Present Illness|643,647|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|643,647|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|643,647|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|643,647|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|History of Present Illness|648,652|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|648,652|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|648,652|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|History of Present Illness|653,659|false|false|false|||showed
Anatomy|Body Location or Region|History of Present Illness|664,676|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|History of Present Illness|664,676|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|History of Present Illness|664,687|false|false|false|C0151699|Intracranial Hemorrhage|intracranial hemorrhage
Event|Event|History of Present Illness|677,687|false|false|false|||hemorrhage
Finding|Pathologic Function|History of Present Illness|677,687|false|false|false|C0019080|Hemorrhage|hemorrhage
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|691,694|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|History of Present Illness|691,694|false|false|false|||CTA
Finding|Gene or Genome|History of Present Illness|691,694|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|691,694|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|History of Present Illness|695,699|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|695,699|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|695,699|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|History of Present Illness|700,706|false|false|false|||showed
Event|Event|History of Present Illness|709,718|false|false|false|||thickened
Finding|Functional Concept|History of Present Illness|719,724|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|726,734|false|false|false|C0224176|Structure of platysma muscle|platysma
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|726,741|false|false|false|C0224176|Structure of platysma muscle|platysma muscle
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|735,741|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|History of Present Illness|735,741|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|History of Present Illness|759,767|false|false|false|||hematoma
Finding|Pathologic Function|History of Present Illness|759,767|false|false|false|C0018944|Hematoma|hematoma
Event|Event|History of Present Illness|774,779|false|false|false|||focus
Finding|Functional Concept|History of Present Illness|774,779|false|false|false|C1285542|Has focus|focus
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|791,799|false|false|false|C0009924|Contrast Media|contrast
Disorder|Injury or Poisoning|History of Present Illness|800,813|false|false|false|C0015379|Extravasation of Diagnostic and Therapeutic Materials|extravasation
Event|Event|History of Present Illness|800,813|false|false|false|||extravasation
Finding|Pathologic Function|History of Present Illness|800,813|false|false|false|C0015376|Extravasation|extravasation
Finding|Functional Concept|History of Present Illness|825,830|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|825,839|false|false|false|C0921006|Right platysma|right platysma
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|825,846|false|false|false|C0921006|Right platysma|right platysma muscle
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|831,839|false|false|false|C0224176|Structure of platysma muscle|platysma
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|831,846|false|false|false|C0224176|Structure of platysma muscle|platysma muscle
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|840,846|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|History of Present Illness|840,846|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|History of Present Illness|857,866|false|false|false|||developed
Finding|Functional Concept|History of Present Illness|869,874|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|869,883|false|false|false|C0524468|Structure of right shoulder region|right shoulder
Anatomy|Body Location or Region|History of Present Illness|875,883|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|875,883|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|875,883|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|History of Present Illness|884,892|false|false|false|||hematoma
Finding|Pathologic Function|History of Present Illness|884,892|false|false|false|C0018944|Hematoma|hematoma
Anatomy|Body Location or Region|History of Present Illness|902,910|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|902,910|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|902,910|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|History of Present Illness|911,916|false|false|false|||plain
Event|Event|History of Present Illness|918,923|false|false|false|||films
Finding|Intellectual Product|History of Present Illness|918,923|false|false|false|C4019020||films
Event|Event|History of Present Illness|931,935|false|false|false|||show
Finding|Intellectual Product|History of Present Illness|936,941|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Congenital Abnormality|History of Present Illness|942,953|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|History of Present Illness|942,953|false|false|false|||abnormality
Finding|Finding|History of Present Illness|942,953|false|false|false|C1704258|Abnormality|abnormality
Event|Event|History of Present Illness|962,966|false|false|false|||seen
Event|Event|History of Present Illness|975,985|false|false|false|||Hematology
Finding|Intellectual Product|History of Present Illness|975,985|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|Hematology
Procedure|Laboratory Procedure|History of Present Illness|975,985|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|Hematology
Event|Event|History of Present Illness|990,994|false|false|false|||gave
Event|Event|History of Present Illness|1003,1007|false|false|false|||dose
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1011,1016|false|false|false|C0701195|DDAVP|DDAVP
Drug|Hormone|History of Present Illness|1011,1016|false|false|false|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|History of Present Illness|1011,1016|false|false|false|C0701195|DDAVP|DDAVP
Finding|Conceptual Entity|History of Present Illness|1023,1029|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|History of Present Illness|1023,1029|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Intellectual Product|History of Present Illness|1023,1029|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Event|Event|History of Present Illness|1036,1041|false|false|false|||assay
Procedure|Laboratory Procedure|History of Present Illness|1036,1041|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Attribute|Clinical Attribute|History of Present Illness|1076,1082|false|false|false|C4255046||report
Event|Event|History of Present Illness|1076,1082|false|false|false|||report
Finding|Intellectual Product|History of Present Illness|1076,1082|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|1076,1082|false|false|false|C0700287|Reporting|report
Attribute|Clinical Attribute|History of Present Illness|1088,1094|false|false|false|C4255046||report
Event|Event|History of Present Illness|1088,1094|false|false|false|||report
Finding|Intellectual Product|History of Present Illness|1088,1094|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|1088,1094|false|false|false|C0700287|Reporting|report
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1101,1111|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|History of Present Illness|1101,1111|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|History of Present Illness|1101,1111|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|History of Present Illness|1101,1111|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|History of Present Illness|1101,1111|false|false|false|||hemoglobin
Finding|Finding|History of Present Illness|1101,1111|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|History of Present Illness|1101,1111|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Finding|Finding|History of Present Illness|1101,1121|false|false|false|C0162119|Hemoglobin below reference range|hemoglobin decreased
Event|Event|History of Present Illness|1112,1121|false|false|false|||decreased
Finding|Functional Concept|History of Present Illness|1156,1162|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|History of Present Illness|1163,1170|false|false|false|||imaging
Finding|Finding|History of Present Illness|1163,1170|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|History of Present Illness|1163,1170|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|History of Present Illness|1186,1192|false|false|false|||showed
Finding|Intellectual Product|History of Present Illness|1193,1199|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Injury or Poisoning|History of Present Illness|1200,1208|false|false|false|C0497561;C0497571;C0497582;C3263723|Female genital injuries;Male Genital Injuries;Traumatic injury;urologic injuries|injuries
Event|Event|History of Present Illness|1200,1208|false|false|false|||injuries
Finding|Body Substance|History of Present Illness|1215,1222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1215,1222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1215,1222|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1223,1226|false|false|false|||saw
Event|Event|History of Present Illness|1259,1264|false|false|false|||found
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1276,1286|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|History of Present Illness|1276,1286|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|History of Present Illness|1276,1286|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|History of Present Illness|1276,1286|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|History of Present Illness|1276,1286|false|false|false|||hemoglobin
Finding|Finding|History of Present Illness|1276,1286|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|History of Present Illness|1276,1286|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Finding|Intellectual Product|History of Present Illness|1321,1325|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|History of Present Illness|1326,1334|false|false|false|||decrease
Finding|Finding|History of Present Illness|1326,1334|false|false|false|C0392756|Reduced|decrease
Finding|Body Substance|History of Present Illness|1341,1348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1341,1348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1341,1348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|History of Present Illness|1370,1373|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1370,1373|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1370,1373|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1370,1373|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1370,1373|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1370,1373|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1370,1373|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1370,1373|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1370,1373|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1370,1373|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1370,1373|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Finding|History of Present Illness|1391,1395|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1391,1395|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1391,1395|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1401,1411|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|History of Present Illness|1401,1411|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|History of Present Illness|1401,1411|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|History of Present Illness|1401,1411|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|History of Present Illness|1401,1411|false|false|false|||hemoglobin
Finding|Finding|History of Present Illness|1401,1411|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|History of Present Illness|1401,1411|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|History of Present Illness|1428,1433|false|false|false|||found
Anatomy|Body Location or Region|History of Present Illness|1455,1460|false|false|false|C0230171|Flank (surface region)|flank
Event|Event|History of Present Illness|1462,1470|false|false|false|||hematoma
Finding|Pathologic Function|History of Present Illness|1462,1470|false|false|false|C0018944|Hematoma|hematoma
Event|Event|History of Present Illness|1481,1489|false|false|false|||referred
Event|Event|History of Present Illness|1496,1503|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1496,1503|false|false|false|C2699424|Concern|concern
Anatomy|Body Space or Junction|History of Present Illness|1508,1523|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Event|Event|History of Present Illness|1525,1530|false|false|false|||bleed
Finding|Pathologic Function|History of Present Illness|1525,1530|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|History of Present Illness|1536,1543|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1536,1543|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1536,1543|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|1536,1547|false|false|false|C0332310|Has patient|patient has
Event|Event|History of Present Illness|1553,1558|false|false|false|||using
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1559,1564|false|false|false|C0701195|DDAVP|DDAVP
Drug|Hormone|History of Present Illness|1559,1564|false|false|false|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|History of Present Illness|1559,1564|false|false|false|C0701195|DDAVP|DDAVP
Event|Event|History of Present Illness|1559,1564|false|false|false|||DDAVP
Event|Event|History of Present Illness|1604,1612|false|false|false|||accident
Event|Event|History of Present Illness|1604,1612|false|false|false|C1690974|Accidental event (event)|accident
Finding|Finding|History of Present Illness|1604,1612|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Finding|Idea or Concept|History of Present Illness|1604,1612|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Phenomenon|Phenomenon or Process|History of Present Illness|1604,1612|false|false|false|C0000924|Accidents|accident
Event|Event|History of Present Illness|1617,1623|false|false|false|||denies
Event|Event|History of Present Illness|1624,1639|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1624,1639|true|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|1644,1656|false|false|false|||palpitations
Finding|Finding|History of Present Illness|1644,1656|false|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|1662,1670|false|false|false|||increase
Finding|Functional Concept|History of Present Illness|1662,1670|true|false|false|C0442805|Increase|increase
Anatomy|Body Location or Region|History of Present Illness|1674,1678|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|1674,1678|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|1674,1678|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|History of Present Illness|1674,1687|false|false|false|C0578454|Neck swelling|neck swelling
Event|Event|History of Present Illness|1679,1687|false|false|false|||swelling
Finding|Finding|History of Present Illness|1679,1687|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|1679,1687|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Intellectual Product|History of Present Illness|1712,1716|false|false|false|C1561540|Transaction counts and value totals - week|week
Attribute|Clinical Attribute|History of Present Illness|1734,1738|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1734,1738|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1734,1738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1734,1738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|History of Present Illness|1746,1751|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|1746,1760|false|false|false|C0524468|Structure of right shoulder region|right shoulder
Anatomy|Body Location or Region|History of Present Illness|1752,1760|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|1752,1760|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1752,1760|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|History of Present Illness|1766,1773|false|false|false|||resting
Event|Event|History of Present Illness|1779,1785|false|false|false|||moving
Event|Event|History of Present Illness|1804,1812|false|false|false|||improved
Finding|Intellectual Product|History of Present Illness|1837,1841|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|History of Present Illness|1856,1863|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1864,1869|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1864,1875|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1864,1875|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|1870,1875|false|false|false|||signs
Finding|Finding|History of Present Illness|1870,1875|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1870,1875|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Idea or Concept|History of Present Illness|1909,1916|false|false|false|C1555582|Initial (abbreviation)|Initial
Event|Event|History of Present Illness|1917,1921|false|false|false|||labs
Lab|Laboratory or Test Result|History of Present Illness|1917,1921|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|History of Present Illness|1922,1934|false|false|false|||demonstrated
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1935,1945|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|History of Present Illness|1935,1945|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|History of Present Illness|1935,1945|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|History of Present Illness|1935,1945|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|History of Present Illness|1935,1945|false|false|false|||hemoglobin
Finding|Finding|History of Present Illness|1935,1945|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|History of Present Illness|1935,1945|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|History of Present Illness|1959,1965|false|false|false|||repeat
Finding|Functional Concept|History of Present Illness|1959,1965|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|History of Present Illness|1976,1987|false|false|false|||Chemistries
Event|Event|History of Present Illness|1992,1997|false|false|false|||coags
Event|Event|History of Present Illness|2003,2015|false|false|false|||unremarkable
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2017,2022|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Drug|Pharmacologic Substance|History of Present Illness|2017,2022|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Finding|Gene or Genome|History of Present Illness|2017,2022|false|false|false|C1366370;C1704822|F8 gene;F8 wt Allele|FVIII
Event|Activity|History of Present Illness|2023,2031|false|false|false|C0441655|Activities|activity
Event|Event|History of Present Illness|2023,2031|false|false|false|||activity
Finding|Daily or Recreational Activity|History of Present Illness|2023,2031|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|History of Present Illness|2023,2031|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|History of Present Illness|2044,2048|false|false|false|||CTAP
Event|Event|History of Present Illness|2069,2081|false|false|false|||demonstrated
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2082,2090|false|false|false|C4083049|Muscle (organ)|muscular
Event|Event|History of Present Illness|2091,2101|false|false|false|||hemorrhage
Finding|Pathologic Function|History of Present Illness|2091,2101|false|false|false|C0019080|Hemorrhage|hemorrhage
Anatomy|Body Location or Region|History of Present Illness|2113,2118|false|false|false|C0230171|Flank (surface region)|flank
Anatomy|Body Space or Junction|History of Present Illness|2127,2142|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Finding|Pathologic Function|History of Present Illness|2127,2148|true|false|false|C0151705|Retroperitoneal Hemorrhage|retroperitoneal bleed
Event|Event|History of Present Illness|2143,2148|false|false|false|||bleed
Finding|Pathologic Function|History of Present Illness|2143,2148|true|false|false|C0019080|Hemorrhage|bleed
Event|Event|History of Present Illness|2152,2163|false|false|false|||preliminary
Event|Event|History of Present Illness|2165,2169|false|false|false|||read
Finding|Body Substance|History of Present Illness|2175,2182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2175,2182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2175,2182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Classification|History of Present Illness|2185,2195|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|History of Present Illness|2185,2195|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|History of Present Illness|2196,2208|false|false|false|||hematologist
Event|Event|History of Present Illness|2224,2233|false|false|false|||contacted
Event|Event|History of Present Illness|2245,2252|false|false|false|||decided
Finding|Body Substance|History of Present Illness|2265,2272|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2265,2272|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2265,2272|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2273,2285|false|false|false|C0011701|desmopressin|desmopressin
Drug|Hormone|History of Present Illness|2273,2285|false|false|false|C0011701|desmopressin|desmopressin
Drug|Pharmacologic Substance|History of Present Illness|2273,2285|false|false|false|C0011701|desmopressin|desmopressin
Event|Event|History of Present Illness|2273,2285|false|false|false|||desmopressin
Finding|Body Substance|History of Present Illness|2304,2311|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2304,2311|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2304,2311|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2316,2320|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|2321,2329|false|false|false|||admitted
Event|Event|History of Present Illness|2342,2352|false|false|false|||management
Event|Occupational Activity|History of Present Illness|2342,2352|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|2342,2352|false|false|false|C0376636|Disease Management|management
Event|Event|History of Present Illness|2360,2366|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|2360,2366|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|2360,2366|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|2360,2369|false|false|false|C0699752|Review of|review of
Event|Event|History of Present Illness|2370,2377|false|false|false|||records
Finding|Idea or Concept|History of Present Illness|2370,2377|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|History of Present Illness|2370,2377|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Body Substance|History of Present Illness|2383,2390|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2383,2390|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2383,2390|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|2383,2394|false|false|false|C0332310|Has patient|patient has
Event|Event|History of Present Illness|2397,2404|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|2397,2407|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|2408,2419|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|2408,2419|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|2421,2429|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|2421,2429|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|History of Present Illness|2440,2452|false|false|false|||circumcision
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2440,2452|false|false|false|C0008819|Male Circumcision|circumcision
Disorder|Disease or Syndrome|History of Present Illness|2464,2469|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|2464,2469|false|false|false|||blood
Finding|Body Substance|History of Present Illness|2464,2469|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2464,2481|false|false|false|C0005841|Blood Transfusion|blood transfusion
Event|Event|History of Present Illness|2470,2481|false|false|false|||transfusion
Finding|Functional Concept|History of Present Illness|2470,2481|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2470,2481|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Event|History of Present Illness|2520,2528|false|false|false|||tendency
Finding|Finding|History of Present Illness|2520,2545|false|false|false|C3889026|Tendency to bruise easily|tendency to bruise easily
Event|Event|History of Present Illness|2532,2538|false|false|false|||bruise
Finding|Finding|History of Present Illness|2539,2545|false|false|false|C0332219|Easy|easily
Event|Event|History of Present Illness|2555,2561|false|false|false|||tested
Event|Event|History of Present Illness|2566,2571|false|false|false|||found
Disorder|Disease or Syndrome|History of Present Illness|2584,2591|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|2584,2591|false|false|false|||disease
Finding|Idea or Concept|History of Present Illness|2607,2613|false|false|false|C0871611|wisdom|wisdom
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2607,2619|false|false|false|C0026369;C1305762|Structure of wisdom tooth|wisdom tooth
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2607,2630|false|false|false|C0204147|Extraction of wisdom tooth|wisdom tooth extraction
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2614,2619|false|false|false|C0040426|Tooth structure|tooth
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2614,2630|false|false|false|C0040440;C1879715|Apical Endodontic Surgery;Tooth Extraction|tooth extraction
Event|Event|History of Present Illness|2620,2630|false|false|false|||extraction
Procedure|Laboratory Procedure|History of Present Illness|2620,2630|false|false|false|C0185115;C0684295|Chemical extraction;Extraction|extraction
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2620,2630|false|false|false|C0185115;C0684295|Chemical extraction;Extraction|extraction
Finding|Body Substance|History of Present Illness|2636,2643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2636,2643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2636,2643|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2656,2660|false|false|false|||late
Event|Event|History of Present Illness|2663,2664|false|false|false|||e
Event|Event|History of Present Illness|2684,2692|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|2684,2692|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|History of Present Illness|2701,2710|false|false|false|||treatment
Finding|Conceptual Entity|History of Present Illness|2701,2710|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|History of Present Illness|2701,2710|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|History of Present Illness|2701,2710|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2701,2710|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2716,2721|false|false|false|C0701195|DDAVP|DDAVP
Drug|Hormone|History of Present Illness|2716,2721|false|false|false|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|History of Present Illness|2716,2721|false|false|false|C0701195|DDAVP|DDAVP
Event|Event|History of Present Illness|2716,2721|false|false|false|||DDAVP
Finding|Body Substance|History of Present Illness|2728,2735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2728,2735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2728,2735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2740,2748|false|false|false|||retested
Event|Event|History of Present Illness|2767,2777|false|false|false|||associated
Event|Event|History of Present Illness|2800,2809|false|false|false|||diagnosed
Disorder|Disease or Syndrome|History of Present Illness|2816,2826|false|false|false|C0019069;C0684275|Hemophilia A|hemophilia
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2834,2839|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Drug|Pharmacologic Substance|History of Present Illness|2834,2839|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Finding|Gene or Genome|History of Present Illness|2834,2839|false|false|false|C1366370;C1704822|F8 gene;F8 wt Allele|FVIII
Event|Activity|History of Present Illness|2840,2848|false|false|false|C0441655|Activities|activity
Event|Event|History of Present Illness|2840,2848|false|false|false|||activity
Finding|Daily or Recreational Activity|History of Present Illness|2840,2848|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|History of Present Illness|2840,2848|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|History of Present Illness|2858,2865|false|false|false|||checked
Event|Event|History of Present Illness|2879,2888|false|false|false|||occasions
Event|Event|History of Present Illness|2900,2907|false|false|false|||testing
Event|Event|History of Present Illness|2908,2914|false|false|false|||normal
Event|Event|History of Present Illness|2916,2922|false|false|false|||though
Finding|Finding|History of Present Illness|2936,2939|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|2936,2939|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Activity|History of Present Illness|2955,2962|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|2955,2962|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|2955,2962|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2970,2975|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|2981,2988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2981,2988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2981,2988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2992,3003|false|false|false|||comfortable
Finding|Finding|History of Present Illness|2992,3003|false|false|false|C5546696|Feeling comfortable|comfortable
Attribute|Clinical Attribute|History of Present Illness|3013,3022|false|false|false|C3864418||complaint
Event|Event|History of Present Illness|3013,3022|false|false|false|||complaint
Finding|Finding|History of Present Illness|3013,3022|false|false|false|C5441521|Complaint (finding)|complaint
Event|Event|History of Present Illness|3026,3032|false|false|false|||Review
Finding|Idea or Concept|History of Present Illness|3026,3032|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|History of Present Illness|3026,3032|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|History of Present Illness|3026,3035|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|History of Present Illness|3026,3043|false|false|false|C0488564;C0488565||Review of Systems
Procedure|Health Care Activity|History of Present Illness|3026,3043|false|false|false|C0489633|Review of systems (procedure)|Review of Systems
Event|Event|History of Present Illness|3036,3043|false|false|false|||Systems
Finding|Functional Concept|History of Present Illness|3036,3043|false|false|false|C0449913|System|Systems
Disorder|Disease or Syndrome|History of Present Illness|3055,3058|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|3055,3058|false|false|false|||HPI
Finding|Finding|History of Present Illness|3055,3058|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|3055,3058|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|3065,3070|false|false|false|||fever
Finding|Finding|History of Present Illness|3065,3070|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|3065,3070|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|3072,3078|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|3072,3078|false|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|3080,3092|false|false|false|C0028081|Night sweats|night sweats
Event|Event|History of Present Illness|3086,3092|false|false|false|||sweats
Finding|Body Substance|History of Present Illness|3086,3092|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|3086,3092|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|History of Present Illness|3094,3102|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|3094,3102|false|false|false|C0018681|Headache|headache
Attribute|Clinical Attribute|History of Present Illness|3104,3110|false|false|false|C2707266||vision
Finding|Organism Function|History of Present Illness|3104,3110|false|false|false|C0042789|Vision|vision
Event|Event|History of Present Illness|3111,3118|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|3111,3118|false|false|false|C0392747|Changing|changes
Event|Event|History of Present Illness|3121,3131|false|false|false|||rhinorrhea
Finding|Sign or Symptom|History of Present Illness|3121,3131|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|History of Present Illness|3133,3143|false|false|false|||congestion
Finding|Pathologic Function|History of Present Illness|3133,3143|false|false|false|C0700148|Congestion|congestion
Finding|Sign or Symptom|History of Present Illness|3145,3149|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|History of Present Illness|3145,3156|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|History of Present Illness|3145,3156|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|History of Present Illness|3145,3156|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|History of Present Illness|3145,3156|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|History of Present Illness|3150,3156|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3150,3156|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|History of Present Illness|3150,3156|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|History of Present Illness|3150,3156|false|false|false|||throat
Finding|Body Substance|History of Present Illness|3150,3156|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|History of Present Illness|3150,3156|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Drug|Organic Chemical|History of Present Illness|3158,3163|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|3158,3163|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|3158,3163|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|3158,3163|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|3165,3174|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|3165,3184|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|3165,3184|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|3178,3184|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|History of Present Illness|3187,3192|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|3187,3192|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|3187,3197|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|3187,3197|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|3193,3197|false|false|false|C2598155||pain
Event|Event|History of Present Illness|3193,3197|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|3193,3197|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3193,3197|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3193,3208|false|false|false|C0000737|Abdominal Pain|pain, abdominal
Anatomy|Body Location or Region|History of Present Illness|3199,3208|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|3199,3213|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|3209,3213|false|false|false|C2598155||pain
Event|Event|History of Present Illness|3209,3213|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|3209,3213|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3209,3213|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|3215,3221|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|3215,3221|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|3215,3221|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|3223,3231|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|3223,3231|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|3233,3241|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|3233,3241|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|3233,3241|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|3244,3256|false|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|3244,3256|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|History of Present Illness|3258,3263|false|false|false|C0018932|Hematochezia|BRBPR
Event|Event|History of Present Illness|3258,3263|false|false|false|||BRBPR
Event|Event|History of Present Illness|3265,3271|false|false|false|||melena
Finding|Pathologic Function|History of Present Illness|3265,3271|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|History of Present Illness|3273,3285|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|History of Present Illness|3273,3285|false|false|false|||hematochezia
Finding|Sign or Symptom|History of Present Illness|3273,3285|false|false|false|C1321898|Blood in stool|hematochezia
Event|Event|History of Present Illness|3287,3294|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|3287,3294|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|History of Present Illness|3296,3305|false|false|false|C0018965|Hematuria|hematuria
Event|Event|History of Present Illness|3296,3305|false|false|false|||hematuria
Finding|Conceptual Entity|Past Medical History|3332,3338|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|Factor
Finding|Functional Concept|Past Medical History|3332,3338|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|Factor
Finding|Intellectual Product|Past Medical History|3332,3338|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|Factor
Drug|Amino Acid, Peptide, or Protein|Past Medical History|3332,3343|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|Factor VIII
Drug|Biologically Active Substance|Past Medical History|3332,3343|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|Factor VIII
Drug|Clinical Drug|Past Medical History|3332,3343|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|Factor VIII
Drug|Pharmacologic Substance|Past Medical History|3332,3343|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|Factor VIII
Finding|Gene or Genome|Past Medical History|3332,3343|false|false|false|C1366370|F8 gene|Factor VIII
Disorder|Disease or Syndrome|Past Medical History|3332,3354|false|false|false|C0019069;C3494187|Factor VIII Deficiency;Hemophilia A|Factor VIII deficiency
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3339,3343|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|Past Medical History|3339,3343|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|Past Medical History|3339,3343|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Disorder|Disease or Syndrome|Past Medical History|3344,3354|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Past Medical History|3344,3354|false|false|false|||deficiency
Finding|Functional Concept|Past Medical History|3344,3354|false|false|false|C0011155|Deficiency|deficiency
Finding|Intellectual Product|Past Medical History|3356,3360|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Body Substance|Family Medical History|3407,3414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|3407,3414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|3407,3414|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|3417,3423|false|false|false|C1546508|Relationship - Mother|mother
Event|Event|Family Medical History|3428,3436|false|false|false|||tendency
Finding|Pathologic Function|Family Medical History|3428,3445|false|false|false|C1458140|Bleeding tendency|tendency to bleed
Event|Event|Family Medical History|3440,3445|false|false|false|||bleed
Procedure|Health Care Activity|General Exam|3470,3479|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3507,3514|false|false|false|||GENERAL
Finding|Classification|General Exam|3507,3514|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3507,3514|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|3516,3521|false|false|false|||lying
Disorder|Disease or Syndrome|General Exam|3530,3533|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|3530,3533|false|false|false|C2346952|Bachelor of Education|bed
Finding|Intellectual Product|General Exam|3538,3543|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3544,3552|false|false|false|||distress
Finding|Finding|General Exam|3544,3552|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3544,3552|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3555,3560|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3562,3566|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3568,3571|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3568,3571|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3568,3571|false|false|false|||MMM
Event|Event|General Exam|3576,3581|false|false|false|||clear
Finding|Idea or Concept|General Exam|3576,3581|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3584,3588|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3584,3588|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3584,3588|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|3590,3596|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3599,3606|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3599,3606|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3608,3611|false|false|false|||RRR
Event|Event|General Exam|3623,3630|false|false|false|||murmurs
Finding|Finding|General Exam|3623,3630|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3632,3639|false|false|false|||gallops
Event|Event|General Exam|3644,3648|false|false|false|||rubs
Finding|Finding|General Exam|3644,3648|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|General Exam|3651,3655|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|General Exam|3651,3655|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|General Exam|3651,3655|false|false|false|C0024115|Lung diseases|LUNG
Event|Event|General Exam|3651,3655|false|false|false|||LUNG
Finding|Finding|General Exam|3651,3655|false|false|false|C0740941|Lung Problem|LUNG
Drug|Amino Acid, Peptide, or Protein|General Exam|3667,3670|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|3667,3670|false|false|false|||CTA
Finding|Gene or Genome|General Exam|3667,3670|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|3667,3670|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|3677,3684|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3677,3684|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3677,3684|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3677,3684|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3686,3690|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|3686,3690|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|3720,3731|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|3733,3737|false|false|false|||Warm
Finding|Finding|General Exam|3733,3737|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3733,3737|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3739,3743|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3744,3752|false|false|false|||perfused
Drug|Food|General Exam|3755,3761|false|false|false|C5890763||PULSES
Event|Event|General Exam|3755,3761|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|3755,3761|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3755,3761|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|General Exam|3769,3775|false|false|false|C5890763||pulses
Event|Event|General Exam|3769,3775|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3769,3775|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3769,3775|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|3807,3813|false|false|false|||intact
Finding|Finding|General Exam|3807,3813|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body System|General Exam|3816,3820|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3816,3820|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3816,3820|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|3816,3820|false|false|false|||SKIN
Finding|Body Substance|General Exam|3816,3820|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3816,3820|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|3822,3831|false|false|false|||Hematomas
Finding|Pathologic Function|General Exam|3822,3831|false|false|false|C0018944|Hematoma|Hematomas
Finding|Functional Concept|General Exam|3835,3840|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|3851,3855|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|3851,3855|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|3851,3855|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|General Exam|3860,3865|false|false|false|C0230171|Flank (surface region)|flank
Finding|Body Substance|General Exam|3871,3880|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3871,3880|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3871,3880|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3871,3880|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3929,3936|false|false|false|||GENERAL
Finding|Classification|General Exam|3929,3936|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3929,3936|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|3938,3943|false|false|false|||lying
Disorder|Disease or Syndrome|General Exam|3952,3955|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|3952,3955|false|false|false|C2346952|Bachelor of Education|bed
Finding|Intellectual Product|General Exam|3960,3965|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3966,3974|false|false|false|||distress
Finding|Finding|General Exam|3966,3974|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3966,3974|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3977,3982|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3984,3988|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3990,3993|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3990,3993|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3990,3993|false|false|false|||MMM
Event|Event|General Exam|3998,4003|false|false|false|||clear
Finding|Idea or Concept|General Exam|3998,4003|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|4006,4010|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|4006,4010|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|4006,4010|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|4012,4018|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|4021,4028|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4021,4028|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|4030,4033|false|false|false|||RRR
Event|Event|General Exam|4045,4052|false|false|false|||murmurs
Finding|Finding|General Exam|4045,4052|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|4054,4061|false|false|false|||gallops
Event|Event|General Exam|4066,4070|false|false|false|||rubs
Finding|Finding|General Exam|4066,4070|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|General Exam|4073,4077|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|General Exam|4073,4077|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|General Exam|4073,4077|false|false|false|C0024115|Lung diseases|LUNG
Event|Event|General Exam|4073,4077|false|false|false|||LUNG
Finding|Finding|General Exam|4073,4077|false|false|false|C0740941|Lung Problem|LUNG
Drug|Amino Acid, Peptide, or Protein|General Exam|4089,4092|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|4089,4092|false|false|false|||CTA
Finding|Gene or Genome|General Exam|4089,4092|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|4089,4092|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|4099,4106|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4099,4106|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4099,4106|false|false|false|||ABDOMEN
Finding|Finding|General Exam|4099,4106|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4108,4112|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|4108,4112|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|4142,4153|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|4155,4159|false|false|false|||Warm
Finding|Finding|General Exam|4155,4159|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4155,4159|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4161,4165|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4166,4174|false|false|false|||perfused
Drug|Food|General Exam|4177,4183|false|false|false|C5890763||PULSES
Event|Event|General Exam|4177,4183|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|4177,4183|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|4177,4183|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|General Exam|4191,4197|false|false|false|C5890763||pulses
Event|Event|General Exam|4191,4197|false|false|false|||pulses
Finding|Physiologic Function|General Exam|4191,4197|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4191,4197|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|4229,4235|false|false|false|||intact
Finding|Finding|General Exam|4229,4235|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body System|General Exam|4238,4242|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4238,4242|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4238,4242|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4238,4242|false|false|false|||SKIN
Finding|Body Substance|General Exam|4238,4242|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4238,4242|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|4244,4253|false|false|false|||Hematomas
Finding|Pathologic Function|General Exam|4244,4253|false|false|false|C0018944|Hematoma|Hematomas
Finding|Functional Concept|General Exam|4257,4262|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|4273,4277|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|4273,4277|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|4273,4277|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|General Exam|4282,4287|false|false|false|C0230171|Flank (surface region)|flank
Procedure|Health Care Activity|General Exam|4310,4319|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Body Substance|General Exam|4321,4330|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4321,4330|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4321,4330|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4321,4330|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4342,4346|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4342,4346|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4361,4366|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4361,4366|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4361,4366|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4367,4370|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4375,4378|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4375,4378|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4375,4378|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4385,4388|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4385,4388|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4385,4388|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4385,4388|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4396,4399|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4396,4399|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4408,4411|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4408,4411|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4408,4411|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4408,4411|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4408,4411|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4415,4418|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4415,4418|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4415,4418|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4415,4418|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4415,4418|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4415,4418|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4424,4428|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4424,4428|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4444,4447|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4464,4469|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4464,4469|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4464,4469|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|4485,4490|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4485,4490|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4485,4490|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4495,4498|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|4495,4498|false|false|false|||Eos
Finding|Gene or Genome|General Exam|4495,4498|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4525,4530|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4525,4530|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4525,4530|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4535,4538|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4535,4538|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4535,4538|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4560,4565|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4560,4565|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4566,4569|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4586,4591|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4586,4591|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4586,4591|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4616,4621|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4616,4621|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4616,4621|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4616,4629|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4616,4629|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4616,4629|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4622,4629|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4622,4629|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4622,4629|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4622,4629|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4622,4629|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4622,4629|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4673,4677|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4673,4677|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4673,4677|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4702,4707|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4702,4707|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4702,4707|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4708,4711|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4716,4719|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4716,4719|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4716,4719|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4726,4729|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4726,4729|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4726,4729|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4726,4729|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4735,4738|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4735,4738|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4746,4749|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4746,4749|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4746,4749|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4746,4749|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4746,4749|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4753,4756|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4753,4756|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4753,4756|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4753,4756|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4753,4756|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4753,4756|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4762,4766|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4762,4766|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4782,4785|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4802,4807|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4802,4807|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4802,4807|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4808,4811|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4816,4819|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4816,4819|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4816,4819|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4826,4829|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4826,4829|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4826,4829|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4826,4829|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4835,4838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4835,4838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4846,4849|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4846,4849|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4846,4849|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4846,4849|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4846,4849|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4853,4856|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4853,4856|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4853,4856|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4853,4856|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4853,4856|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4853,4856|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4862,4866|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4862,4866|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4882,4885|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4902,4907|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4902,4907|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4902,4907|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4908,4911|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4916,4919|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4916,4919|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4916,4919|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4926,4929|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4926,4929|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4926,4929|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4926,4929|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4935,4938|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4935,4938|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4946,4949|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4946,4949|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4946,4949|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4946,4949|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4946,4949|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4953,4956|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4953,4956|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4953,4956|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4953,4956|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4953,4956|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4953,4956|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4962,4966|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4962,4966|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4982,4985|false|false|false|C0201617|Primed lymphocyte test|Plt
Finding|Body Substance|General Exam|5002,5007|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5002,5007|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5002,5007|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|5002,5013|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|5008,5013|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5008,5013|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Finding|Idea or Concept|General Exam|5028,5033|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|5053,5058|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5053,5058|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5053,5058|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|5053,5064|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|5059,5064|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|5059,5064|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|5065,5068|false|false|false|||NEG
Finding|Finding|General Exam|5065,5068|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|5069,5076|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|5069,5076|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|5069,5076|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|General Exam|5077,5080|false|false|false|||NEG
Finding|Finding|General Exam|5077,5080|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|5081,5088|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|5081,5088|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|5081,5088|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|5081,5088|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|5081,5088|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|General Exam|5093,5100|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5093,5100|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5093,5100|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5093,5100|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5093,5100|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5093,5100|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|5101,5104|false|false|false|||NEG
Finding|Finding|General Exam|5101,5104|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|5105,5111|false|false|false|C0022634|Ketones|Ketone
Event|Event|General Exam|5112,5115|false|false|false|||NEG
Finding|Finding|General Exam|5112,5115|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|5124,5127|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|5136,5139|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5153,5156|false|false|false|||NEG
Finding|Finding|General Exam|5153,5156|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|5169,5174|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5169,5174|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5169,5174|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|5169,5178|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|General Exam|5175,5178|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5175,5178|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5175,5178|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|5182,5185|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|General Exam|5200,5205|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|General Exam|5200,5205|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5200,5205|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|General Exam|5200,5205|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Disorder|Disease or Syndrome|General Exam|5211,5214|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|General Exam|5211,5214|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|General Exam|5211,5214|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|General Exam|5211,5214|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|General Exam|5211,5214|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|General Exam|5211,5214|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|General Exam|5211,5214|false|false|false|||Epi
Finding|Gene or Genome|General Exam|5211,5214|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|General Exam|5211,5214|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|General Exam|5211,5214|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|General Exam|5229,5234|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5229,5234|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5229,5234|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|5229,5241|false|false|false|C0455910|Mucus in urine (finding)|URINE Mucous
Finding|Body Substance|General Exam|5235,5241|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|Mucous
Event|Event|General Exam|5242,5246|false|false|false|||RARE
Finding|Gene or Genome|General Exam|5242,5246|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Event|Event|General Exam|5248,5255|false|false|false|||IMAGING
Finding|Finding|General Exam|5248,5255|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|5248,5255|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|5256,5263|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|5256,5263|false|false|false|C0947630|Scientific Study|STUDIES
Drug|Amino Acid, Peptide, or Protein|General Exam|5271,5275|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Drug|Enzyme|General Exam|5271,5275|false|false|false|C3538970|Choline-Phosphate Cytidylyltransferase A|CT A
Finding|Intellectual Product|General Exam|5278,5283|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Pathologic Function|General Exam|5278,5294|false|false|false|C0333276|Acute hemorrhage|Acute hemorrhage
Event|Event|General Exam|5284,5294|false|false|false|||hemorrhage
Finding|Pathologic Function|General Exam|5284,5294|false|false|false|C0019080|Hemorrhage|hemorrhage
Finding|Functional Concept|General Exam|5301,5306|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|General Exam|5307,5316|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Location or Region|General Exam|5307,5322|false|false|false|C0446499|Posterior abdominal surface region|posterior flank
Anatomy|Body Location or Region|General Exam|5317,5322|false|false|false|C0230171|Flank (surface region)|flank
Anatomy|Body Part, Organ, or Organ Component|General Exam|5323,5334|false|false|false|C1995013|Set of muscles|musculature
Finding|Finding|General Exam|5340,5348|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|General Exam|5340,5348|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Anatomy|Body Part, Organ, or Organ Component|General Exam|5349,5357|false|false|false|C0934502|anatomical layer|layering
Anatomy|Body Part, Organ, or Organ Component|General Exam|5411,5422|false|false|false|C1995013|Set of muscles|musculature
Event|Event|General Exam|5428,5438|false|false|false|||hemorrhage
Finding|Pathologic Function|General Exam|5428,5438|false|false|false|C0019080|Hemorrhage|hemorrhage
Disorder|Injury or Poisoning|General Exam|5450,5463|true|false|false|C0015379|Extravasation of Diagnostic and Therapeutic Materials|extravasation
Event|Event|General Exam|5450,5463|false|false|false|||extravasation
Finding|Pathologic Function|General Exam|5450,5463|true|false|false|C0015376|Extravasation|extravasation
Event|Event|General Exam|5465,5469|false|false|false|||seen
Finding|Finding|General Exam|5471,5479|false|false|false|C0332148|Probable diagnosis|Probable
Event|Event|General Exam|5484,5492|false|false|false|||hematoma
Finding|Pathologic Function|General Exam|5484,5492|false|true|false|C0018944|Hematoma|hematoma
Disorder|Disease or Syndrome|General Exam|5499,5508|false|true|false|C0751438|Posterior pituitary disease|posterior
Finding|Functional Concept|General Exam|5509,5513|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|5509,5519|false|false|false|C0733996|Structure of left flank|left flank
Anatomy|Body Location or Region|General Exam|5514,5519|false|false|false|C0230171|Flank (surface region)|flank
Event|Event|Hospital Course|5570,5577|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5570,5577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5570,5577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5570,5577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5570,5580|false|false|false|C0262926|Medical History|history of
Finding|Intellectual Product|Hospital Course|5581,5585|false|false|false|C1547225|Mild Severity of Illness Code|mild
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5586,5591|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Drug|Pharmacologic Substance|Hospital Course|5586,5591|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Event|Event|Hospital Course|5586,5591|false|false|false|||FVIII
Finding|Gene or Genome|Hospital Course|5586,5591|false|false|false|C1366370;C1704822|F8 gene;F8 wt Allele|FVIII
Disorder|Disease or Syndrome|Hospital Course|5592,5602|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Hospital Course|5592,5602|false|false|false|||deficiency
Finding|Functional Concept|Hospital Course|5592,5602|false|false|false|C0011155|Deficiency|deficiency
Event|Event|Hospital Course|5608,5616|false|false|false|||presents
Finding|Daily or Recreational Activity|Hospital Course|5623,5635|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Finding|Finding|Hospital Course|5623,5635|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Event|Event|Hospital Course|5636,5644|false|false|false|||accident
Event|Event|Hospital Course|5636,5644|false|false|false|C1690974|Accidental event (event)|accident
Finding|Finding|Hospital Course|5636,5644|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Finding|Idea or Concept|Hospital Course|5636,5644|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Phenomenon|Phenomenon or Process|Hospital Course|5636,5644|false|false|false|C0000924|Accidents|accident
Event|Event|Hospital Course|5659,5668|false|false|false|||hematomas
Finding|Pathologic Function|Hospital Course|5659,5668|false|false|false|C0018944|Hematoma|hematomas
Event|Event|Hospital Course|5674,5681|false|false|false|||falling
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5682,5692|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|5682,5692|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|5682,5692|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|5682,5692|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Hospital Course|5682,5692|false|false|false|||hemoglobin
Finding|Finding|Hospital Course|5682,5692|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|5682,5692|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|Hospital Course|5693,5703|false|false|false|||concerning
Finding|Idea or Concept|Hospital Course|5708,5715|false|false|false|C0549178|Continuous|ongoing
Event|Event|Hospital Course|5716,5724|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|5716,5724|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Conceptual Entity|Hospital Course|5729,5735|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|FACTOR
Finding|Functional Concept|Hospital Course|5729,5735|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|FACTOR
Finding|Intellectual Product|Hospital Course|5729,5735|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|FACTOR
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5729,5740|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|FACTOR VIII
Drug|Biologically Active Substance|Hospital Course|5729,5740|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|FACTOR VIII
Drug|Clinical Drug|Hospital Course|5729,5740|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|FACTOR VIII
Drug|Pharmacologic Substance|Hospital Course|5729,5740|false|false|false|C0015506;C1307126;C2732002;C2732016;C4520835|Factor viii (antihemophilic factor, human) per i.u.;Human Coagulation Factor VIII/Von Willebrand Factor Complex;antihemophilic factor, human recombinant;factor VIII;factor VIII, human|FACTOR VIII
Finding|Gene or Genome|Hospital Course|5729,5740|false|false|false|C1366370|F8 gene|FACTOR VIII
Disorder|Disease or Syndrome|Hospital Course|5729,5751|false|false|false|C0019069;C3494187|Factor VIII Deficiency;Hemophilia A|FACTOR VIII DEFICIENCY
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5736,5740|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|Hospital Course|5736,5740|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|Hospital Course|5736,5740|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Disorder|Disease or Syndrome|Hospital Course|5741,5751|false|false|false|C0162429|Malnutrition|DEFICIENCY
Event|Event|Hospital Course|5741,5751|false|false|false|||DEFICIENCY
Finding|Functional Concept|Hospital Course|5741,5751|false|false|false|C0011155|Deficiency|DEFICIENCY
Finding|Pathologic Function|Hospital Course|5762,5771|false|false|false|C0018944|Hematoma|HEMATOMAS
Finding|Body Substance|Hospital Course|5773,5780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|5773,5780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|5773,5780|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|5781,5790|false|false|false|||presented
Finding|Idea or Concept|Hospital Course|5781,5790|false|false|false|C0449450|Presentation|presented
Event|Event|Hospital Course|5805,5817|false|false|false|||snowboarding
Finding|Daily or Recreational Activity|Hospital Course|5805,5817|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Finding|Finding|Hospital Course|5805,5817|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Event|Event|Hospital Course|5818,5826|false|false|false|||accident
Event|Event|Hospital Course|5818,5826|false|false|false|C1690974|Accidental event (event)|accident
Finding|Finding|Hospital Course|5818,5826|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Finding|Idea or Concept|Hospital Course|5818,5826|false|false|false|C1546397;C2046386|Admission Type - Accident;history of accident|accident
Phenomenon|Phenomenon or Process|Hospital Course|5818,5826|false|false|false|C0000924|Accidents|accident
Event|Event|Hospital Course|5841,5848|false|false|false|||imaging
Finding|Finding|Hospital Course|5841,5848|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|5841,5848|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Hospital Course|5853,5860|false|false|false|||notable
Anatomy|Body Location or Region|Hospital Course|5865,5869|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|5865,5869|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|5865,5869|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|Hospital Course|5874,5882|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|Hospital Course|5874,5882|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5874,5882|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Event|Event|Hospital Course|5883,5892|false|false|false|||hematomas
Finding|Pathologic Function|Hospital Course|5883,5892|false|false|false|C0018944|Hematoma|hematomas
Event|Event|Hospital Course|5900,5912|false|false|false|||reevaluation
Disorder|Disease or Syndrome|Hospital Course|5920,5923|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5920,5923|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|5920,5923|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5920,5923|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|5920,5923|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|5920,5923|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|5920,5923|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|5920,5923|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|5920,5923|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|5920,5923|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|5920,5923|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|Hospital Course|5929,5936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5929,5936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5929,5936|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5941,5946|false|false|false|||found
Anatomy|Body Location or Region|Hospital Course|5958,5963|false|false|false|C0230171|Flank (surface region)|flank
Event|Event|Hospital Course|5964,5972|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|5964,5972|false|false|false|C0018944|Hematoma|hematoma
Disorder|Injury or Poisoning|Hospital Course|5980,5987|false|false|false|C0000921|Accidental Falls|falling
Event|Event|Hospital Course|5980,5987|false|false|false|||falling
Finding|Finding|Hospital Course|5980,5987|false|false|false|C0085639|Falls|falling
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5988,5998|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|5988,5998|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|5988,5998|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|5988,5998|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Hospital Course|5988,5998|false|false|false|||hemoglobin
Finding|Finding|Hospital Course|5988,5998|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|5988,5998|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|Hospital Course|6010,6017|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|6010,6017|false|false|false|C2699424|Concern|concern
Anatomy|Body Space or Junction|Hospital Course|6023,6038|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Finding|Pathologic Function|Hospital Course|6023,6044|false|false|false|C0151705|Retroperitoneal Hemorrhage|retroperitoneal bleed
Event|Event|Hospital Course|6039,6044|false|false|false|||bleed
Finding|Pathologic Function|Hospital Course|6039,6044|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|Hospital Course|6046,6050|false|false|false|||CTAP
Event|Event|Hospital Course|6061,6073|false|false|false|||demonstrated
Finding|Pathologic Function|Hospital Course|6074,6082|false|false|false|C0018944|Hematoma|hematoma
Anatomy|Body Location or Region|Hospital Course|6093,6098|false|false|false|C0230171|Flank (surface region)|flank
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6099,6110|false|false|false|C1995013|Set of muscles|musculature
Disorder|Injury or Poisoning|Hospital Course|6126,6139|true|false|false|C0015379|Extravasation of Diagnostic and Therapeutic Materials|extravasation
Event|Event|Hospital Course|6126,6139|false|false|false|||extravasation
Finding|Pathologic Function|Hospital Course|6126,6139|true|false|false|C0015376|Extravasation|extravasation
Event|Event|Hospital Course|6148,6153|false|false|false|||given
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6158,6163|false|false|false|C0701195|DDAVP|DDAVP
Drug|Hormone|Hospital Course|6158,6163|false|false|false|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|Hospital Course|6158,6163|false|false|false|C0701195|DDAVP|DDAVP
Event|Event|Hospital Course|6158,6163|false|false|false|||DDAVP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6169,6174|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Drug|Pharmacologic Substance|Hospital Course|6169,6174|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Finding|Gene or Genome|Hospital Course|6169,6174|false|false|false|C1366370;C1704822|F8 gene;F8 wt Allele|FVIII
Event|Activity|Hospital Course|6175,6183|false|false|false|C0441655|Activities|activity
Event|Event|Hospital Course|6175,6183|false|false|false|||activity
Finding|Daily or Recreational Activity|Hospital Course|6175,6183|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Hospital Course|6175,6183|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Anatomy|Cell Component|Hospital Course|6199,6202|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|6199,6202|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|Hospital Course|6212,6218|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|6212,6218|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Body Substance|Hospital Course|6224,6231|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6224,6231|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6224,6231|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6232,6240|false|false|false|||declined
Event|Event|Hospital Course|6249,6258|false|false|false|||inpatient
Finding|Idea or Concept|Hospital Course|6249,6258|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|6249,6258|false|false|false|C1555324|inpatient encounter|inpatient
Event|Activity|Hospital Course|6259,6269|false|false|false|C1283169||monitoring
Event|Event|Hospital Course|6259,6269|false|false|false|||monitoring
Procedure|Health Care Activity|Hospital Course|6259,6269|false|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|Hospital Course|6279,6289|false|false|false|||hematology
Finding|Intellectual Product|Hospital Course|6279,6289|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|Hospital Course|6279,6289|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Event|Event|Hospital Course|6290,6301|false|false|false|||recommended
Event|Event|Hospital Course|6302,6311|false|false|false|||continued
Finding|Classification|Hospital Course|6312,6322|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|6312,6322|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6323,6333|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|6323,6333|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|6323,6333|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|6323,6333|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Hospital Course|6323,6333|false|false|false|||hemoglobin
Finding|Finding|Hospital Course|6323,6333|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|6323,6333|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Activity|Hospital Course|6335,6345|false|false|false|C1283169||monitoring
Event|Event|Hospital Course|6335,6345|false|false|false|||monitoring
Procedure|Health Care Activity|Hospital Course|6335,6345|false|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|Hospital Course|6359,6364|false|false|false|||think
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6373,6378|true|false|true|C0701195|DDAVP|DDAVP
Drug|Hormone|Hospital Course|6373,6378|true|false|true|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|Hospital Course|6373,6378|true|false|true|C0701195|DDAVP|DDAVP
Event|Event|Hospital Course|6373,6378|false|false|false|||DDAVP
Event|Event|Hospital Course|6383,6392|false|false|false|||indicated
Event|Event|Hospital Course|6400,6406|false|false|false|||normal
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6407,6412|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Drug|Pharmacologic Substance|Hospital Course|6407,6412|false|false|false|C2732002|antihemophilic factor, human recombinant|FVIII
Finding|Gene or Genome|Hospital Course|6407,6412|false|false|false|C1366370;C1704822|F8 gene;F8 wt Allele|FVIII
Event|Event|Hospital Course|6413,6418|false|false|false|||level
Event|Event|Hospital Course|6440,6446|false|false|false|||ISSUES
Disorder|Disease or Syndrome|Hospital Course|6450,6453|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6450,6453|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|6450,6453|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6450,6453|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|6450,6453|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|6450,6453|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|6450,6453|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|6450,6453|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|6450,6453|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|6450,6453|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|6450,6453|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Anatomy|Cell Component|Hospital Course|6464,6467|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|6464,6467|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|Hospital Course|6498,6503|false|false|false|||avoid
Event|Activity|Hospital Course|6514,6522|false|false|false|C0441655|Activities|activity
Event|Event|Hospital Course|6514,6522|false|false|false|||activity
Finding|Daily or Recreational Activity|Hospital Course|6514,6522|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Hospital Course|6514,6522|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Hospital Course|6525,6529|false|false|false|||Code
Event|Occupational Activity|Hospital Course|6525,6529|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|6525,6529|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|Hospital Course|6549,6558|false|false|false|||Emergency
Finding|Finding|Hospital Course|6549,6558|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Hospital Course|6549,6558|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Hospital Course|6549,6558|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Hospital Course|6549,6558|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Hospital Course|6549,6558|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Hospital Course|6549,6558|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|Hospital Course|6549,6566|false|false|false|C1552023|emergency contact|Emergency Contact
Event|Activity|Hospital Course|6559,6566|false|false|false|C3812666|Personal Contact|Contact
Finding|Functional Concept|Hospital Course|6559,6566|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|Hospital Course|6559,6566|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|Hospital Course|6559,6566|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|Hospital Course|6559,6566|false|false|false|C0392367|Physical contact|Contact
Attribute|Clinical Attribute|Hospital Course|6587,6598|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6587,6598|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6587,6598|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6587,6598|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|6587,6611|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|6602,6611|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|6602,6611|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|6630,6640|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|6630,6640|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|6630,6645|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|6641,6645|false|false|false|||list
Finding|Intellectual Product|Hospital Course|6641,6645|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|6649,6657|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|6662,6670|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|6662,6670|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|6662,6670|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|6662,6670|false|false|false|||complete
Finding|Functional Concept|Hospital Course|6662,6670|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6662,6670|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6675,6687|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Hormone|Hospital Course|6675,6687|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Pharmacologic Substance|Hospital Course|6675,6687|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Clinical Drug|Hospital Course|6675,6693|false|false|false|C3212180||Desmopressin Nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6688,6693|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|6688,6693|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|6688,6693|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|6688,6693|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|6688,6693|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|6688,6693|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Disorder|Disease or Syndrome|Hospital Course|6702,6705|false|false|false|C0027609|Neonatal Abstinence Syndrome|NAS
Drug|Organic Chemical|Hospital Course|6702,6705|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Drug|Substance|Hospital Course|6702,6705|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Event|Event|Hospital Course|6702,6705|false|false|false|||NAS
Finding|Finding|Hospital Course|6702,6705|false|false|false|C5552704||NAS
Finding|Gene or Genome|Hospital Course|6706,6709|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|6710,6718|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|6710,6718|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|6723,6732|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6723,6732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6723,6732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6723,6732|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6723,6732|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6723,6744|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6733,6744|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6733,6744|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6733,6744|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6733,6744|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6749,6762|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6749,6762|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|6749,6762|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6749,6762|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Attribute|Clinical Attribute|Hospital Course|6778,6782|false|false|false|C2598155||pain
Event|Event|Hospital Course|6778,6782|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6778,6782|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6778,6782|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6787,6799|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Hormone|Hospital Course|6787,6799|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Pharmacologic Substance|Hospital Course|6787,6799|false|false|false|C0011701|desmopressin|Desmopressin
Drug|Clinical Drug|Hospital Course|6787,6805|false|false|false|C3212180||Desmopressin Nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6800,6805|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|6800,6805|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|6800,6805|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|6800,6805|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|6800,6805|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|6800,6805|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Disorder|Disease or Syndrome|Hospital Course|6814,6817|false|false|false|C0027609|Neonatal Abstinence Syndrome|NAS
Drug|Organic Chemical|Hospital Course|6814,6817|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Drug|Substance|Hospital Course|6814,6817|false|false|false|C0067783;C0068453|N-acetylserotonin;Tobacco containing mixture|NAS
Event|Event|Hospital Course|6814,6817|false|false|false|||NAS
Finding|Finding|Hospital Course|6814,6817|false|false|false|C5552704||NAS
Finding|Gene or Genome|Hospital Course|6818,6821|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|6822,6830|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|6822,6830|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Classification|Hospital Course|6835,6845|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|6835,6845|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|Hospital Course|6846,6849|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|Hospital Course|6846,6849|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|Hospital Course|6850,6854|false|false|false|||Work
Event|Occupational Activity|Hospital Course|6850,6854|false|false|false|C0043227|Work|Work
Anatomy|Cell Component|Hospital Course|6855,6858|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|Hospital Course|6855,6858|false|false|false|||CBC
Procedure|Laboratory Procedure|Hospital Course|6855,6858|false|false|false|C0009555|Complete Blood Count|CBC
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6879,6889|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|6879,6889|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|6879,6889|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|6879,6889|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Hospital Course|6879,6889|false|false|false|||hemoglobin
Finding|Finding|Hospital Course|6879,6889|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|6879,6889|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|Hospital Course|6906,6915|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6906,6915|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6906,6915|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6906,6915|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6906,6915|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6906,6927|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6906,6927|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6916,6927|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6916,6927|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6916,6927|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6929,6933|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6929,6933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6929,6933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6929,6933|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|6936,6945|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6936,6945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6936,6945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6936,6945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6936,6945|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6936,6955|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6946,6955|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6946,6955|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6946,6955|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6946,6955|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6946,6955|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Hospital Course|6968,6973|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6974,6982|false|false|false|C4083049|Muscle (organ)|muscular
Event|Event|Hospital Course|6983,6991|false|false|false|||hematoma
Finding|Pathologic Function|Hospital Course|6983,6991|false|false|false|C0018944|Hematoma|hematoma
Finding|Functional Concept|Hospital Course|6993,6998|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|6993,7004|false|false|false|C0733995|Structure of right flank|right flank
Anatomy|Body Location or Region|Hospital Course|6999,7004|false|false|false|C0230171|Flank (surface region)|flank
Disorder|Disease or Syndrome|Hospital Course|7007,7017|false|false|false|C0019069;C0684275|Hemophilia A|Hemophilia
Event|Event|Hospital Course|7007,7017|false|false|false|||Hemophilia
Event|Event|Hospital Course|7019,7025|false|false|false|||factor
Finding|Conceptual Entity|Hospital Course|7019,7025|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Functional Concept|Hospital Course|7019,7025|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Finding|Intellectual Product|Hospital Course|7019,7025|false|false|false|C1521761;C2827422;C5400797|Factor;Feelings about Genomic Testing Results;Mathematical Factor|factor
Disorder|Disease or Syndrome|Hospital Course|7031,7041|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Hospital Course|7031,7041|false|false|false|||deficiency
Finding|Functional Concept|Hospital Course|7031,7041|false|false|false|C0011155|Deficiency|deficiency
Finding|Mental Process|Discharge Condition|7066,7072|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|7066,7079|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|7066,7079|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|7073,7079|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|7073,7079|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7081,7086|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|7081,7086|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|7091,7099|false|false|false|||coherent
Finding|Finding|Discharge Condition|7091,7099|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|7101,7106|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|7101,7123|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|7101,7123|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|7110,7123|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|7110,7123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|7110,7123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|7125,7130|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|7125,7130|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|7125,7130|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|7125,7130|false|false|false|||Alert
Finding|Finding|Discharge Condition|7125,7130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|7125,7130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|7125,7130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|7135,7146|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|7135,7146|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|7148,7156|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|7148,7156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|7148,7156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|7157,7163|false|false|false|C5889824||Status
Event|Event|Discharge Condition|7157,7163|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|7157,7163|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7165,7175|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|7165,7175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|7165,7175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|7165,7175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|7165,7175|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|7178,7189|false|false|false|||Independent
Finding|Finding|Discharge Condition|7178,7189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|7178,7189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|7239,7247|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|7239,7247|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|7239,7247|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|Discharge Instructions|7285,7293|false|false|false|||admitted
Disorder|Injury or Poisoning|Discharge Instructions|7299,7307|false|false|false|C0009938|Contusions|bruising
Event|Event|Discharge Instructions|7299,7307|false|false|false|||bruising
Finding|Finding|Discharge Instructions|7299,7307|false|false|false|C2136686|reported bruising (history)|bruising
Event|Event|Discharge Instructions|7316,7321|false|false|false|||right
Finding|Functional Concept|Discharge Instructions|7316,7321|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|Discharge Instructions|7332,7335|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|7332,7335|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Disorder|Disease or Syndrome|Discharge Instructions|7336,7341|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7336,7341|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7336,7341|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7342,7348|false|false|false|||counts
Event|Event|Discharge Instructions|7357,7369|false|false|false|||snowboarding
Finding|Daily or Recreational Activity|Discharge Instructions|7357,7369|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Finding|Finding|Discharge Instructions|7357,7369|false|false|false|C1138838;C2350009|Snowboarding (activity);snowboarding (history)|snowboarding
Event|Event|Discharge Instructions|7370,7374|false|false|false|||fall
Finding|Finding|Discharge Instructions|7370,7374|false|false|false|C0085639|Falls|fall
Event|Event|Discharge Instructions|7387,7394|false|false|false|||history
Finding|Conceptual Entity|Discharge Instructions|7387,7394|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Discharge Instructions|7387,7394|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Discharge Instructions|7387,7394|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Discharge Instructions|7387,7397|false|false|false|C0262926|Medical History|history of
Attribute|Clinical Attribute|Discharge Instructions|7387,7408|false|false|false|C3176015||history of hemophilia
Disorder|Disease or Syndrome|Discharge Instructions|7398,7408|false|false|false|C0019069;C0684275|Hemophilia A|hemophilia
Event|Event|Discharge Instructions|7398,7408|false|false|false|||hemophilia
Event|Event|Discharge Instructions|7417,7426|false|false|false|||important
Event|Event|Discharge Instructions|7430,7438|false|false|false|||evaluate
Event|Event|Discharge Instructions|7449,7457|false|false|false|||bleeding
Finding|Pathologic Function|Discharge Instructions|7449,7457|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Discharge Instructions|7468,7472|false|false|false|||show
Finding|Functional Concept|Discharge Instructions|7475,7480|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7481,7489|false|false|false|C4083049|Muscle (organ)|muscular
Anatomy|Body Location or Region|Discharge Instructions|7490,7495|false|false|false|C0230171|Flank (surface region)|flank
Disorder|Disease or Syndrome|Discharge Instructions|7496,7501|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7496,7501|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7496,7501|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7502,7512|false|false|false|||collection
Finding|Conceptual Entity|Discharge Instructions|7502,7512|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Discharge Instructions|7502,7512|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Discharge Instructions|7502,7512|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Discharge Instructions|7502,7512|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7527,7531|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|Discharge Instructions|7527,7531|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|Discharge Instructions|7527,7531|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|Discharge Instructions|7532,7537|false|false|false|||level
Event|Event|Discharge Instructions|7554,7562|false|false|false|||received
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|7566,7571|false|false|false|C0701195|DDAVP|DDAVP
Drug|Hormone|Discharge Instructions|7566,7571|false|false|false|C0701195|DDAVP|DDAVP
Drug|Pharmacologic Substance|Discharge Instructions|7566,7571|false|false|false|C0701195|DDAVP|DDAVP
Event|Event|Discharge Instructions|7572,7577|false|false|false|||under
Event|Activity|Discharge Instructions|7583,7587|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|7583,7587|false|false|false|||care
Finding|Finding|Discharge Instructions|7583,7587|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|7583,7587|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Discharge Instructions|7594,7599|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7594,7599|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7594,7599|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7600,7606|false|false|false|||counts
Event|Event|Discharge Instructions|7612,7618|false|false|false|||stable
Finding|Intellectual Product|Discharge Instructions|7612,7618|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|7622,7630|false|false|false|||improved
Finding|Finding|Discharge Instructions|7622,7630|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|Discharge Instructions|7622,7630|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Idea or Concept|Discharge Instructions|7638,7641|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|7638,7641|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|7646,7655|false|false|false|||admission
Procedure|Health Care Activity|Discharge Instructions|7646,7655|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Discharge Instructions|7665,7674|false|false|false|||important
Event|Event|Discharge Instructions|7688,7699|false|false|false|||participate
Event|Activity|Discharge Instructions|7718,7728|false|false|false|C0441655|Activities|activities
Event|Event|Discharge Instructions|7718,7728|false|false|false|||activities
Finding|Finding|Discharge Instructions|7718,7728|false|false|false|C2239122|activities (history)|activities
Event|Event|Discharge Instructions|7747,7752|false|false|false|||bleed
Finding|Pathologic Function|Discharge Instructions|7747,7752|false|false|false|C0019080|Hemorrhage|bleed
Disorder|Disease or Syndrome|Discharge Instructions|7762,7772|false|false|false|C0019069;C0684275|Hemophilia A|hemophilia
Event|Event|Discharge Instructions|7762,7772|false|false|false|||hemophilia
Finding|Pathologic Function|Discharge Instructions|7774,7782|false|false|false|C0019080|Hemorrhage|Bleeding
Event|Event|Discharge Instructions|7825,7829|false|false|false|||life
Finding|Idea or Concept|Discharge Instructions|7825,7829|false|false|false|C0376558|Life|life
Procedure|Diagnostic Procedure|Discharge Instructions|7825,7829|false|false|false|C1522684|Laser-Induced Fluorescence Endoscopy|life
Event|Event|Discharge Instructions|7830,7841|false|false|false|||threatening
Disorder|Disease or Syndrome|Discharge Instructions|7860,7865|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7860,7865|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7860,7865|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7873,7880|false|false|false|||checked
Anatomy|Body Location or Region|Discharge Instructions|7888,7892|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|7888,7892|false|false|false|C1546778||site
Event|Event|Discharge Instructions|7916,7922|false|false|false|||Follow
Finding|Intellectual Product|Discharge Instructions|7945,7951|false|false|false|C2348314|Doctor - Title|doctor
Finding|Idea or Concept|Discharge Instructions|7958,7962|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Intellectual Product|Discharge Instructions|7963,7967|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Activity|Discharge Instructions|7992,7996|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|7992,7996|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|7992,7996|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|7992,8001|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|7992,8001|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|8004,8012|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|8013,8025|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|8013,8025|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|8013,8025|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

