 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|160,169|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|160,169|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|160,169|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|181,190|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|181,190|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|181,190|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|201,205|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|201,205|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|206,215|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|218,227|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|218,227|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|236,251|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|242,251|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|242,251|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|242,251|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|253,260|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|253,272|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|264,272|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|264,272|false|false|false|C0015264|Exertion|exertion
Finding|Classification|SIMPLE_SEGMENT|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|302,311|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|302,311|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|321,328|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|321,328|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|321,328|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|321,328|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|321,331|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|321,347|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|321,347|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|332,339|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|332,339|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|332,347|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|340,347|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|360,367|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|360,370|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|374,377|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|374,377|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|379,382|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|379,382|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|379,382|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|379,382|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|379,382|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|387,390|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|387,390|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|387,390|false|false|false|C1413980|DES gene|DES
Finding|Functional Concept|SIMPLE_SEGMENT|396,404|false|false|false|C0475224|Ischemic|ischemic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|413,421|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|SIMPLE_SEGMENT|413,433|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|422,433|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|422,433|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Organic Chemical|SIMPLE_SEGMENT|442,451|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|442,451|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|442,451|false|false|false|||torsemide
Anatomy|Body Location or Region|SIMPLE_SEGMENT|459,462|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|459,462|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|459,462|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|468,476|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|493,500|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|493,500|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|493,500|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|493,512|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|504,512|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|504,512|false|false|false|C0015264|Exertion|exertion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|514,517|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|514,526|false|false|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|SIMPLE_SEGMENT|518,526|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|518,526|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|518,526|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|SIMPLE_SEGMENT|535,541|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|535,541|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|535,541|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|535,541|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|535,541|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|543,547|false|false|false|||gain
Finding|Body Substance|SIMPLE_SEGMENT|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|571,575|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|583,588|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|583,588|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|583,588|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|583,596|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|Heart Failure
Finding|Functional Concept|SIMPLE_SEGMENT|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Event|Event|SIMPLE_SEGMENT|635,640|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|670,677|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|670,677|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|670,677|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|670,689|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|681,689|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|681,689|false|false|false|C0015264|Exertion|exertion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|694,697|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|694,697|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|694,697|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|SIMPLE_SEGMENT|721,736|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|721,736|false|false|false|C0019993|Hospitalization|hospitalization
Anatomy|Body Location or Region|SIMPLE_SEGMENT|741,744|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|741,744|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|741,744|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|SIMPLE_SEGMENT|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|771,778|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|791,800|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|791,800|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|791,800|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|817,825|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|830,838|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|851,858|false|false|false|||holiday
Event|Event|SIMPLE_SEGMENT|851,858|false|false|false|C0019843|Holidays|holiday
Event|Event|SIMPLE_SEGMENT|863,871|false|false|false|||indulged
Finding|Finding|SIMPLE_SEGMENT|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|SIMPLE_SEGMENT|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|887,891|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|887,891|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|887,891|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|887,891|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|896,905|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|918,925|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|918,925|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|918,925|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|918,937|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|929,937|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|929,937|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|939,945|true|false|false|||Denies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|950,960|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|950,960|true|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|950,960|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|962,975|true|false|false|||noncompliance
Anatomy|Body Location or Region|SIMPLE_SEGMENT|977,982|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|977,982|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|977,987|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|977,987|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|983,987|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|983,987|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|983,987|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|983,987|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|989,1001|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|989,1001|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|1003,1015|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|1003,1015|false|false|false|C0030252|Palpitations|palpitations
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1028,1031|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|1028,1031|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|1028,1031|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|SIMPLE_SEGMENT|1043,1051|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1043,1051|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1043,1051|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1043,1061|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|SIMPLE_SEGMENT|1043,1061|false|false|false|C2024889||exercise tolerance
Event|Event|SIMPLE_SEGMENT|1052,1061|false|false|false|||tolerance
Finding|Finding|SIMPLE_SEGMENT|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|SIMPLE_SEGMENT|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|SIMPLE_SEGMENT|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|SIMPLE_SEGMENT|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Event|Event|SIMPLE_SEGMENT|1063,1069|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|1063,1069|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|1073,1077|false|false|false|||walk
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1082,1086|false|false|false|C0016504|Foot|feet
Event|Event|SIMPLE_SEGMENT|1093,1102|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|1093,1102|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1093,1102|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Body Substance|SIMPLE_SEGMENT|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1129,1134|false|false|false|||found
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1156,1161|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1156,1161|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1163,1172|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|1163,1178|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1173,1178|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1173,1178|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1173,1178|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1199,1207|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|1199,1207|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|1211,1215|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1211,1215|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1211,1215|false|false|false|C0582103|Medical Examination|exam
Finding|Body Substance|SIMPLE_SEGMENT|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1236,1239|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1236,1239|false|false|false|C0039985|Plain chest X-ray|CXR
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|SIMPLE_SEGMENT|1241,1244|false|false|false|||BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|1241,1244|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1241,1244|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|SIMPLE_SEGMENT|1264,1268|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|1280,1285|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1280,1285|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|1280,1285|false|false|false|||Lasix
Finding|Idea or Concept|SIMPLE_SEGMENT|1298,1305|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1306,1312|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1356,1364|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1356,1364|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1356,1364|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1356,1364|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1366,1372|false|false|false|||vitals
Finding|Body Substance|SIMPLE_SEGMENT|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1410,1414|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|1421,1431|false|false|false|||remarkable
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|1436,1442|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|1436,1442|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1436,1442|false|false|false|C0337443|Sodium measurement|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1448,1456|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|SIMPLE_SEGMENT|1448,1456|false|false|false|||Chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|1448,1456|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1448,1456|false|false|false|C0201952|Chloride measurement|Chloride
Drug|Organic Chemical|SIMPLE_SEGMENT|1469,1475|false|false|false|C0074722|sodium bicarbonate|Bicarb
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1469,1475|false|false|false|C0074722|sodium bicarbonate|Bicarb
Event|Event|SIMPLE_SEGMENT|1469,1475|false|false|false|||Bicarb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1480,1483|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1480,1483|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|1480,1483|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1480,1483|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1489,1499|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|1489,1499|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|1489,1499|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|1489,1499|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1489,1499|false|false|false|C0201975|Creatinine measurement|Creatinine
Finding|Body Substance|SIMPLE_SEGMENT|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1517,1519|false|false|false|||CK
Finding|Body Substance|SIMPLE_SEGMENT|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|SIMPLE_SEGMENT|1562,1565|false|false|false|||BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|1562,1565|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1562,1565|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Finding|Body Substance|SIMPLE_SEGMENT|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1594,1597|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1594,1597|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|1594,1597|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1594,1597|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1594,1597|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|SIMPLE_SEGMENT|1603,1606|false|false|false|||Hct
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1603,1606|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1603,1606|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Anatomy|Cell|SIMPLE_SEGMENT|1614,1622|false|false|false|C0005821|Blood Platelets|Platelet
Anatomy|Cell|SIMPLE_SEGMENT|1628,1631|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1637,1647|false|false|false|||Urinalysis
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1637,1647|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|Urinalysis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1648,1653|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|1654,1661|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|1654,1661|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Event|Event|SIMPLE_SEGMENT|1667,1676|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1667,1676|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|1680,1683|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|1680,1683|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1680,1683|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|1685,1692|false|false|false|||notable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1709,1712|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1709,1712|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|1709,1712|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1709,1712|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Social Behavior|SIMPLE_SEGMENT|1725,1733|false|false|false|C0678975|inferiority|inferior
Event|Event|SIMPLE_SEGMENT|1755,1764|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|1755,1764|false|true|false|C0442739||unchanged
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1791,1796|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|1820,1828|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|1835,1841|false|false|false|||coming
Event|Event|SIMPLE_SEGMENT|1850,1852|false|false|false|||ED
Finding|Finding|SIMPLE_SEGMENT|1857,1877|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1862,1869|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1862,1869|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1862,1869|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1862,1869|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1862,1869|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1862,1877|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1870,1877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1881,1893|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|1881,1893|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1898,1906|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|1898,1906|false|false|false|||diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1914,1917|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1914,1917|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|1914,1917|false|false|false|||CVA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1919,1929|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1930,1939|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1940,1946|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1940,1946|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1940,1946|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1958,1961|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1958,1961|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1958,1961|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1958,1961|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1958,1961|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1979,1982|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|1979,1982|false|false|false|||BMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2014,2041|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2025,2033|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2025,2041|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2034,2041|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2034,2041|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2043,2055|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|SIMPLE_SEGMENT|2043,2055|false|false|false|||claudication
Finding|Finding|SIMPLE_SEGMENT|2043,2055|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2070,2078|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|SIMPLE_SEGMENT|2080,2087|false|false|false|||managed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2105,2110|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|2105,2113|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2114,2117|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|2114,2117|false|false|false|||CKD
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2119,2127|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|2119,2127|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|2119,2127|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2141,2145|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|2141,2145|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2146,2156|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2146,2162|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Event|SIMPLE_SEGMENT|2157,2162|false|false|false|||rings
Finding|Functional Concept|SIMPLE_SEGMENT|2165,2171|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2165,2179|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2172,2179|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2172,2179|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2172,2179|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2172,2179|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2185,2191|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2185,2191|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2185,2191|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2185,2191|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2185,2199|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2192,2199|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2192,2199|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2192,2199|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2192,2199|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2201,2207|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2201,2207|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|2208,2212|false|false|false|||died
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2231,2235|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2231,2235|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2231,2235|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2231,2235|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2231,2243|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2236,2243|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2236,2243|false|false|false|||disease
Finding|Idea or Concept|SIMPLE_SEGMENT|2246,2252|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|SIMPLE_SEGMENT|2253,2257|false|false|false|||died
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|2280,2287|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|2288,2293|false|false|false|||cause
Finding|Conceptual Entity|SIMPLE_SEGMENT|2288,2293|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|SIMPLE_SEGMENT|2288,2293|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2305,2308|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2305,2308|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2305,2308|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2305,2308|true|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2305,2308|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2319,2326|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2319,2326|true|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|2328,2333|true|false|false|||death
Finding|Finding|SIMPLE_SEGMENT|2328,2333|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|SIMPLE_SEGMENT|2328,2333|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|SIMPLE_SEGMENT|2328,2333|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|SIMPLE_SEGMENT|2350,2357|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2350,2357|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2350,2357|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2350,2357|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2350,2360|true|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|2350,2367|true|false|false|C0455471|History of malignant neoplasm|history of cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2361,2367|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2361,2367|true|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|2371,2379|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2371,2379|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2371,2379|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2371,2379|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2371,2384|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2371,2384|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2380,2384|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2380,2384|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2380,2384|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2386,2395|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|SIMPLE_SEGMENT|2396,2404|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2396,2404|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2396,2404|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2396,2416|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2396,2416|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|2405,2416|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|2405,2416|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|2405,2416|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|2424,2425|false|false|false|||T
Event|Event|SIMPLE_SEGMENT|2457,2460|false|false|false|||sat
Event|Event|SIMPLE_SEGMENT|2477,2486|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2477,2486|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2487,2493|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|2487,2493|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|2487,2493|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2487,2493|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2487,2493|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|2501,2508|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2501,2508|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2501,2508|false|false|false|C3812897|General medical service|GENERAL
Event|Event|SIMPLE_SEGMENT|2510,2514|false|false|false|||WDWN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2516,2521|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2516,2521|false|false|false|||obese
Event|Event|SIMPLE_SEGMENT|2523,2530|false|false|false|||sitting
Finding|Finding|SIMPLE_SEGMENT|2523,2538|false|false|false|C1280451|Sitting upright|sitting upright
Event|Event|SIMPLE_SEGMENT|2531,2538|false|false|false|||upright
Finding|Intellectual Product|SIMPLE_SEGMENT|2531,2538|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|2531,2538|false|false|false|C1550585|Entity Handling - upright|upright
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2542,2545|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|2542,2545|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2542,2545|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2550,2553|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2550,2553|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2550,2553|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2550,2553|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|2555,2559|false|false|false|||AOx3
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2562,2566|false|false|false|C2713234||Mood
Event|Event|SIMPLE_SEGMENT|2562,2566|false|false|false|||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|2568,2574|false|false|false|||affect
Event|Event|SIMPLE_SEGMENT|2575,2586|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2590,2595|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2597,2601|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2603,2609|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2603,2609|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2603,2609|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2603,2609|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2610,2619|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2610,2619|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2621,2626|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|2621,2626|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|2628,2632|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2634,2645|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2634,2645|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2634,2645|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|2634,2645|true|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|2634,2645|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|2634,2645|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|2634,2645|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|2661,2667|true|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|2661,2667|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|2671,2679|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2671,2679|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2687,2691|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2687,2691|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|2687,2691|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|2687,2691|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2687,2698|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|2692,2698|true|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|2692,2698|true|false|false|C1561514||mucosa
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2700,2704|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2706,2712|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|2706,2712|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|2718,2721|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2718,2721|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2732,2739|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2732,2739|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2741,2744|false|false|false|||PMI
Finding|Finding|SIMPLE_SEGMENT|2741,2744|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|SIMPLE_SEGMENT|2741,2744|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2760,2777|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2772,2777|false|false|false|C0282173|Space (Astronomy)|space
Event|Event|SIMPLE_SEGMENT|2779,2792|false|false|false|||midclavicular
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|2794,2798|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|2794,2798|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|2827,2834|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2827,2834|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|2835,2839|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2840,2847|true|false|false|||gallops
Event|Event|SIMPLE_SEGMENT|2853,2860|true|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|2853,2860|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|2862,2867|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2870,2875|false|false|false|C0024109|Lung|LUNGS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2877,2881|true|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2877,2881|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|2877,2881|true|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|2887,2896|true|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|2887,2896|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2901,2917|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|2901,2921|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2911,2917|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2911,2917|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|2918,2921|true|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|2918,2921|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2918,2921|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|SIMPLE_SEGMENT|2923,2931|true|false|false|||dyspneic
Finding|Finding|SIMPLE_SEGMENT|2923,2931|true|false|false|C0277854|dyspneic|dyspneic
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2940,2943|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|SIMPLE_SEGMENT|2940,2943|false|false|false|C0082420|Endoglin, human|end
Event|Event|SIMPLE_SEGMENT|2940,2943|false|false|false|||end
Finding|Functional Concept|SIMPLE_SEGMENT|2940,2943|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|SIMPLE_SEGMENT|2940,2943|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Event|Event|SIMPLE_SEGMENT|2954,2962|false|false|false|||sentence
Finding|Intellectual Product|SIMPLE_SEGMENT|2954,2962|false|false|false|C0876929|Sentence|sentence
Event|Event|SIMPLE_SEGMENT|2974,2982|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2974,2982|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2990,2996|false|false|false|C0817096|Chest|thorax
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2990,2996|false|false|false|C0153661|Malignant neoplasm of thorax|thorax
Finding|Finding|SIMPLE_SEGMENT|2999,3015|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Event|Event|SIMPLE_SEGMENT|3007,3015|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|3007,3015|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3019,3026|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3019,3026|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3019,3026|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3019,3026|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3028,3032|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3028,3032|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|3034,3038|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|3043,3046|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|3043,3046|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|3050,3060|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3050,3060|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3050,3060|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3064,3075|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3080,3085|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3080,3085|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3080,3085|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3089,3094|false|false|false|C0230444|Shin|shins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3099,3106|true|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|3107,3113|true|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|3107,3113|true|false|false|C0006318|Bruit|bruits
Drug|Food|SIMPLE_SEGMENT|3117,3123|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|3117,3123|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3117,3123|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3117,3123|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3126,3132|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|SIMPLE_SEGMENT|3133,3139|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3133,3139|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3133,3139|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3133,3139|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|3153,3162|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3153,3162|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3153,3162|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|SIMPLE_SEGMENT|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3164,3173|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|SIMPLE_SEGMENT|3174,3182|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3174,3182|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3174,3182|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3174,3194|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3174,3194|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|SIMPLE_SEGMENT|3183,3194|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3183,3194|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|3183,3194|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|3202,3203|false|false|false|||T
Event|Event|SIMPLE_SEGMENT|3235,3238|false|false|false|||sat
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3250,3256|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|3250,3256|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|3250,3256|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|3250,3256|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|3250,3256|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|3263,3270|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3263,3270|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3263,3270|false|false|false|C3812897|General medical service|GENERAL
Event|Event|SIMPLE_SEGMENT|3272,3276|false|false|false|||WDWN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3278,3283|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3278,3283|false|false|false|||obese
Event|Event|SIMPLE_SEGMENT|3285,3292|false|false|false|||sitting
Finding|Finding|SIMPLE_SEGMENT|3285,3300|false|false|false|C1280451|Sitting upright|sitting upright
Event|Event|SIMPLE_SEGMENT|3293,3300|false|false|false|||upright
Finding|Intellectual Product|SIMPLE_SEGMENT|3293,3300|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|3293,3300|false|false|false|C1550585|Entity Handling - upright|upright
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3304,3307|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|3304,3307|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3304,3307|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3312,3315|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3312,3315|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3312,3315|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3312,3315|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|3317,3321|false|false|false|||AOx3
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3324,3328|false|false|false|C2713234||Mood
Event|Event|SIMPLE_SEGMENT|3324,3328|false|false|false|||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|3330,3336|false|false|false|||affect
Event|Event|SIMPLE_SEGMENT|3337,3348|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3352,3357|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3359,3363|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3365,3371|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3365,3371|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3365,3371|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3365,3371|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3372,3381|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3372,3381|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3383,3388|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3383,3388|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|3390,3394|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3396,3407|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3396,3407|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3396,3407|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3396,3407|true|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|3396,3407|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|3396,3407|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|3396,3407|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3423,3429|true|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|3423,3429|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|3433,3441|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3433,3441|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3449,3453|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3449,3453|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|3449,3453|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|3449,3453|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3449,3460|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|3454,3460|true|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3454,3460|true|false|false|C1561514||mucosa
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3462,3466|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3462,3466|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3462,3466|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3468,3474|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|3468,3474|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|3480,3483|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3480,3483|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3494,3501|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3494,3501|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|3503,3506|false|false|false|||PMI
Finding|Finding|SIMPLE_SEGMENT|3503,3506|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|SIMPLE_SEGMENT|3503,3506|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3522,3539|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3534,3539|false|false|false|C0282173|Space (Astronomy)|space
Event|Event|SIMPLE_SEGMENT|3541,3554|false|false|false|||midclavicular
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|3556,3560|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|3556,3560|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|3589,3596|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|3589,3596|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|3597,3601|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|3602,3609|true|false|false|||gallops
Event|Event|SIMPLE_SEGMENT|3615,3622|true|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|3615,3622|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|3624,3629|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3632,3637|false|false|false|C0024109|Lung|LUNGS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3639,3643|true|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3639,3643|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|3639,3643|true|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|3649,3658|true|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|3649,3658|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3663,3679|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|3663,3683|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3673,3679|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|3673,3679|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|3680,3683|true|false|false|||use
Finding|Functional Concept|SIMPLE_SEGMENT|3680,3683|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3680,3683|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Finding|SIMPLE_SEGMENT|3696,3704|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|3705,3710|false|false|false|||trace
Finding|Functional Concept|SIMPLE_SEGMENT|3705,3710|false|false|false|C1883002|Sequence Chromatogram|trace
Finding|Finding|SIMPLE_SEGMENT|3712,3728|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Event|Event|SIMPLE_SEGMENT|3720,3728|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|3720,3728|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3732,3739|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3732,3739|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3732,3739|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3732,3739|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3741,3745|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3741,3745|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|3747,3751|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|3756,3759|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|3756,3759|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|3763,3773|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3763,3773|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3763,3773|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3777,3788|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3798,3805|true|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|3806,3812|true|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|3806,3812|true|false|false|C0006318|Bruit|bruits
Drug|Food|SIMPLE_SEGMENT|3816,3822|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|3816,3822|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3816,3822|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3816,3822|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3825,3831|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|SIMPLE_SEGMENT|3832,3838|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3832,3838|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3832,3838|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3832,3838|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|3852,3861|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3852,3861|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3852,3861|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Procedure|Health Care Activity|SIMPLE_SEGMENT|3883,3892|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3893,3897|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3893,3897|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3910,3915|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3910,3915|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3910,3915|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3916,3919|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3924,3927|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3924,3927|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3924,3927|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3934,3937|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3934,3937|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3934,3937|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3934,3937|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3943,3946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3943,3946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3954,3957|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3954,3957|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3954,3957|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3954,3957|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3954,3957|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3964,3967|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3964,3967|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3964,3967|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3964,3967|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3964,3967|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3964,3967|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3973,3977|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3973,3977|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4006,4009|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4026,4031|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4026,4031|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4026,4031|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4044,4050|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4068,4071|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|4068,4071|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4068,4071|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4170,4175|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4170,4175|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4170,4175|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4180,4183|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4180,4183|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4180,4183|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4205,4210|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4205,4210|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4205,4210|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4211,4214|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|SIMPLE_SEGMENT|4211,4214|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|SIMPLE_SEGMENT|4211,4214|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4224,4227|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4224,4227|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Finding|Gene or Genome|SIMPLE_SEGMENT|4224,4227|false|false|false|C1425698;C4723885|DDX41 gene;DDX41 wt Allele|Abs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4228,4231|false|false|false|C0389252|RET protein, human|Ret
Event|Event|SIMPLE_SEGMENT|4228,4231|false|false|false|||Ret
Finding|Gene or Genome|SIMPLE_SEGMENT|4228,4231|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|SIMPLE_SEGMENT|4228,4231|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4249,4254|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4249,4254|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4249,4254|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4249,4262|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4249,4262|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4249,4262|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4255,4262|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4255,4262|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4255,4262|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4255,4262|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4255,4262|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4255,4262|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|4300,4301|false|false|false|||5
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4313,4317|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4313,4317|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4313,4317|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4343,4348|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4343,4348|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4343,4348|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4349,4354|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4349,4354|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4349,4354|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4349,4354|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4352,4356|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4387,4392|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4387,4392|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4387,4392|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4393,4398|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4393,4398|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4393,4398|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4393,4398|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4396,4400|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4427,4432|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4427,4432|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4427,4432|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4427,4440|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4433,4440|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4433,4440|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4433,4440|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Body Substance|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4462,4471|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4472,4476|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4472,4476|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4495,4500|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4495,4500|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4495,4500|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4501,4504|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4510,4513|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4510,4513|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4510,4513|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4520,4523|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4520,4523|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4520,4523|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4520,4523|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4529,4532|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4529,4532|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4540,4543|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4540,4543|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4540,4543|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4540,4543|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4540,4543|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4547,4550|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4547,4550|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4547,4550|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4547,4550|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4547,4550|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4547,4550|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4556,4560|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4556,4560|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4588,4591|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4608,4613|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4608,4613|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4608,4613|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4630,4635|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4630,4635|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4630,4635|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4630,4643|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4630,4643|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4630,4643|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4636,4643|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4636,4643|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4636,4643|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4636,4643|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4636,4643|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4636,4643|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4690,4694|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4690,4694|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4690,4694|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4719,4724|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4719,4724|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4719,4724|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4719,4732|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4725,4732|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4725,4732|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4725,4732|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4754,4761|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4754,4761|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4754,4761|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|4772,4775|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4772,4775|false|false|false|C0039985|Plain chest X-ray|CXR
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4776,4784|false|false|false|C2926606||FINDINGS
Event|Event|SIMPLE_SEGMENT|4776,4784|false|false|false|||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|4776,4784|false|false|false|C2607943|findings aspects|FINDINGS
Finding|Intellectual Product|SIMPLE_SEGMENT|4796,4800|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4801,4810|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4801,4810|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|4801,4810|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|4801,4816|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4811,4816|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4811,4816|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4811,4816|false|false|false|C0013604|Edema|edema
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|4835,4841|false|false|false|C1514562|Protein Domain|region
Event|Event|SIMPLE_SEGMENT|4835,4841|false|false|false|||region
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4861,4874|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4861,4874|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|4882,4886|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4893,4897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4893,4897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4893,4897|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|4893,4897|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|4893,4897|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|4911,4919|false|false|false|C0332149|Possible|possible
Anatomy|Tissue|SIMPLE_SEGMENT|4936,4943|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4936,4943|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|4936,4953|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|4944,4953|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|4944,4953|false|false|false|C0013687|effusion|effusions
Finding|Finding|SIMPLE_SEGMENT|4956,4964|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|4956,4964|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|4966,4978|false|false|false|||cardiomegaly
Finding|Finding|SIMPLE_SEGMENT|4966,4978|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|SIMPLE_SEGMENT|4988,4992|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|4996,5000|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5004,5014|false|false|false|||tortuosity
Finding|Functional Concept|SIMPLE_SEGMENT|5023,5033|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5023,5048|false|false|false|C1522460;C3163626|Descending thoracic aorta;Thoracic aorta|descending thoracic aorta
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5034,5042|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5034,5042|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5034,5048|false|false|false|C1522460;C4037977|Chest>Aorta.thoracic;Thoracic aorta|thoracic aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5043,5048|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|5043,5048|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Intellectual Product|SIMPLE_SEGMENT|5054,5059|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5060,5067|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|5060,5067|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5068,5081|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|5068,5081|true|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|5068,5081|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|5085,5095|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5085,5095|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5085,5095|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5098,5102|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5103,5112|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5103,5112|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5103,5112|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|5103,5118|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5113,5118|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5113,5118|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5113,5118|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|5137,5141|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5148,5152|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5148,5152|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5148,5152|false|false|false|C0024115|Lung diseases|lung
Event|Event|SIMPLE_SEGMENT|5148,5152|false|false|false|||lung
Finding|Finding|SIMPLE_SEGMENT|5148,5152|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5154,5167|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|5154,5167|false|false|false|||consolidation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5196,5201|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5196,5201|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5196,5201|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|5210,5222|false|false|false|||superimposed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5223,5232|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5223,5232|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5223,5232|false|false|false|C3714514|Infection|infection
Finding|Intellectual Product|SIMPLE_SEGMENT|5237,5242|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5243,5251|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5243,5258|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5243,5258|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|5264,5268|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|5264,5268|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|5269,5272|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|5285,5292|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5285,5295|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|5285,5308|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5296,5308|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5296,5308|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5310,5313|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5310,5313|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|5310,5313|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|5310,5313|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5310,5313|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5318,5321|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|5318,5321|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|5318,5321|false|false|false|C1413980|DES gene|DES
Finding|Functional Concept|SIMPLE_SEGMENT|5328,5336|false|false|false|C0475224|Ischemic|ischemic
Event|Event|SIMPLE_SEGMENT|5337,5339|false|false|false|||MR
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5344,5352|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|SIMPLE_SEGMENT|5344,5364|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5353,5364|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|5353,5364|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5377,5380|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5377,5380|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5377,5380|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|5377,5380|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|5387,5395|false|false|false|||admitted
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5400,5403|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5400,5403|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|5404,5416|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|5404,5416|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|SIMPLE_SEGMENT|5421,5426|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|SIMPLE_SEGMENT|5430,5437|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5430,5437|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5438,5465|false|false|false|C0581377|Decompensated cardiac failure|decompensated heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5452,5457|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5452,5457|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5452,5457|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5452,5465|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|5458,5465|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|5467,5476|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|5485,5492|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|5485,5492|false|false|false|C0542559|contextual factors|setting
Finding|Finding|SIMPLE_SEGMENT|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|5506,5510|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|5506,5510|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|5506,5510|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5506,5510|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|5516,5523|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|5516,5523|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5516,5523|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5516,5535|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|5527,5535|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|5527,5535|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|5537,5546|false|false|false|||decreased
Event|Event|SIMPLE_SEGMENT|5548,5556|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5548,5556|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5548,5556|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5548,5566|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|SIMPLE_SEGMENT|5548,5566|false|false|false|C2024889||exercise tolerance
Event|Event|SIMPLE_SEGMENT|5557,5566|false|false|false|||tolerance
Finding|Finding|SIMPLE_SEGMENT|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|SIMPLE_SEGMENT|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|SIMPLE_SEGMENT|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|SIMPLE_SEGMENT|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5572,5577|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5572,5577|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5572,5577|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|5579,5587|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|5579,5587|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|5591,5595|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|5591,5595|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5591,5595|false|false|false|C0582103|Medical Examination|exam
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|SIMPLE_SEGMENT|5606,5609|false|false|false|||BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|5606,5609|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5606,5609|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5634,5640|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|5634,5640|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|5634,5640|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|5634,5640|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|5634,5640|false|false|false|C1305866|Weighing patient|weight
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5645,5654|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5645,5654|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5645,5654|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5645,5665|false|false|false|C0242073|Pulmonary congestion|pulmonary congestion
Event|Event|SIMPLE_SEGMENT|5655,5665|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|5655,5665|false|false|false|C0700148|Congestion|congestion
Event|Event|SIMPLE_SEGMENT|5669,5672|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5669,5672|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|5681,5691|true|false|false|||discovered
Event|Event|SIMPLE_SEGMENT|5695,5703|true|false|false|||pharmacy
Finding|Intellectual Product|SIMPLE_SEGMENT|5695,5703|true|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|SIMPLE_SEGMENT|5695,5703|true|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|SIMPLE_SEGMENT|5704,5710|true|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|5704,5710|true|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|5704,5710|true|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Body Substance|SIMPLE_SEGMENT|5716,5723|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5716,5723|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5716,5723|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5732,5738|true|false|false|||filled
Drug|Organic Chemical|SIMPLE_SEGMENT|5740,5749|true|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5740,5749|true|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|5740,5749|true|false|false|||torsemide
Finding|Classification|SIMPLE_SEGMENT|5761,5771|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5761,5771|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body System|SIMPLE_SEGMENT|5772,5782|true|false|false|C0007226|Cardiovascular system|Cardiology
Event|Activity|SIMPLE_SEGMENT|5783,5794|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|5783,5794|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|5810,5820|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|5824,5829|false|false|false|||start
Event|Event|SIMPLE_SEGMENT|5830,5836|false|false|false|||taking
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5841,5850|false|false|false|C0041199|Troponin|Troponins
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5841,5850|false|false|false|C0041199|Troponin|Troponins
Event|Event|SIMPLE_SEGMENT|5841,5850|false|false|false|||Troponins
Event|Event|SIMPLE_SEGMENT|5863,5871|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5863,5871|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5863,5871|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5863,5871|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|5876,5885|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5876,5885|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|5895,5901|false|false|false|||placed
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|SIMPLE_SEGMENT|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Event|Event|SIMPLE_SEGMENT|5907,5911|false|false|false|||salt
Drug|Substance|SIMPLE_SEGMENT|5916,5921|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5916,5921|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5916,5921|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|SIMPLE_SEGMENT|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Idea or Concept|SIMPLE_SEGMENT|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Intellectual Product|SIMPLE_SEGMENT|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Procedure|Health Care Activity|SIMPLE_SEGMENT|5923,5938|false|false|false|C0425422|Dietary Restriction|restricted diet
Drug|Food|SIMPLE_SEGMENT|5934,5938|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|5934,5938|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|5934,5938|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5934,5938|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|5948,5956|false|false|false|||diuresed
Drug|Organic Chemical|SIMPLE_SEGMENT|5965,5970|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5965,5970|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|5965,5970|false|false|false|||Lasix
Finding|Intellectual Product|SIMPLE_SEGMENT|5992,5996|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|5997,6009|false|false|false|||transitioned
Drug|Organic Chemical|SIMPLE_SEGMENT|6016,6025|true|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6016,6025|true|false|false|C0076840|torsemide|torsemide
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6043,6049|true|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|6043,6049|true|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|6043,6049|true|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|6043,6049|true|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|6043,6049|true|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|6051,6058|false|false|false|||decline
Anatomy|Cell Component|SIMPLE_SEGMENT|6063,6066|true|false|false|C3850088|Neutrophil Extracellular Traps|net
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6063,6066|true|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6063,6066|true|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Drug|Enzyme|SIMPLE_SEGMENT|6063,6066|true|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Finding|Gene or Genome|SIMPLE_SEGMENT|6063,6066|true|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Finding|Intellectual Product|SIMPLE_SEGMENT|6063,6066|true|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Finding|Receptor|SIMPLE_SEGMENT|6063,6066|true|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Event|Event|SIMPLE_SEGMENT|6067,6075|true|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6067,6075|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6067,6075|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6067,6075|true|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|6067,6089|true|false|false|C0429652|Negative fluid balance|negative fluid balance
Drug|Substance|SIMPLE_SEGMENT|6076,6081|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6076,6081|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6076,6081|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Organism Function|SIMPLE_SEGMENT|6076,6089|true|false|false|C0016284|Fluid Balance|fluid balance
Drug|Organic Chemical|SIMPLE_SEGMENT|6082,6089|true|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6082,6089|true|false|false|C4319618|Balance (substance)|balance
Event|Event|SIMPLE_SEGMENT|6082,6089|true|false|false|||balance
Finding|Finding|SIMPLE_SEGMENT|6082,6089|true|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|SIMPLE_SEGMENT|6082,6089|true|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6082,6089|true|false|false|C2174421|examination of balance|balance
Finding|Idea or Concept|SIMPLE_SEGMENT|6093,6097|true|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|6093,6097|true|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|SIMPLE_SEGMENT|6108,6114|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6108,6114|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6115,6120|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6115,6120|false|false|false|C0042075|Urologic Diseases|renal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6115,6129|false|false|false|C0232804|Renal function|renal function
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6115,6129|false|false|false|C0022662|Kidney Function Tests|renal function
Event|Event|SIMPLE_SEGMENT|6121,6129|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6131,6143|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6131,6143|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Event|Event|SIMPLE_SEGMENT|6131,6143|false|false|false|||Electrolytes
Event|Event|SIMPLE_SEGMENT|6144,6152|false|false|false|||repleted
Finding|Idea or Concept|SIMPLE_SEGMENT|6157,6161|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|6157,6161|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|SIMPLE_SEGMENT|6162,6164|false|false|false|||Mg
Event|Event|SIMPLE_SEGMENT|6185,6194|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6198,6202|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6198,6202|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6198,6202|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6203,6213|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6203,6213|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|SIMPLE_SEGMENT|6203,6213|false|false|false|||carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6221,6224|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6221,6224|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6221,6224|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6221,6224|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6221,6224|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6227,6239|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6227,6239|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6255,6265|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6255,6265|false|false|false|C0065374|lisinopril|lisinopril
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6281,6286|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6281,6286|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6281,6286|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|6288,6296|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6288,6296|false|false|false|C0033095||pressure
Drug|Organic Chemical|SIMPLE_SEGMENT|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|6297,6304|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|SIMPLE_SEGMENT|6309,6318|false|false|false|||increased
Finding|Idea or Concept|SIMPLE_SEGMENT|6319,6323|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6319,6323|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6319,6323|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6324,6334|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6324,6334|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|6324,6334|false|false|false|||nifedipine
Event|Event|SIMPLE_SEGMENT|6335,6337|false|false|false|||CR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6355,6358|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6355,6358|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6355,6358|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6355,6358|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6355,6358|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|6362,6369|false|false|false|||achieve
Finding|Idea or Concept|SIMPLE_SEGMENT|6370,6374|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|6370,6374|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6375,6378|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6375,6378|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6375,6378|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|6375,6378|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|6375,6378|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6375,6378|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|SIMPLE_SEGMENT|6385,6395|false|false|false|||Discharged
Finding|Finding|SIMPLE_SEGMENT|6401,6406|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|6401,6406|false|false|false|C0587267;C3810854|Close;Closed|close
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|6407,6410|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|6407,6410|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|6407,6410|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|6431,6438|false|false|false|||weights
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6431,6438|false|false|false|C3812400|Weights - exercise activity|weights
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6443,6448|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6443,6448|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6443,6448|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|6443,6457|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|6443,6457|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|6443,6457|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|6449,6457|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6449,6457|false|false|false|C0033095||pressure
Drug|Organic Chemical|SIMPLE_SEGMENT|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|6459,6466|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6471,6483|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|6471,6483|false|false|false|||Hypertension
Event|Event|SIMPLE_SEGMENT|6493,6502|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6506,6510|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6506,6510|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6506,6510|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6511,6521|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6511,6521|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|SIMPLE_SEGMENT|6511,6521|false|false|false|||carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6529,6532|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6529,6532|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6529,6532|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6529,6532|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6529,6532|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6535,6547|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6535,6547|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6563,6573|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6563,6573|false|false|false|C0065374|lisinopril|lisinopril
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6589,6594|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6589,6594|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6589,6594|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|6596,6604|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6596,6604|false|false|false|C0033095||pressure
Drug|Organic Chemical|SIMPLE_SEGMENT|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|6605,6612|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|SIMPLE_SEGMENT|6617,6626|false|false|false|||increased
Finding|Idea or Concept|SIMPLE_SEGMENT|6627,6631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6627,6631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6627,6631|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6632,6642|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6632,6642|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|6632,6642|false|false|false|||nifedipine
Event|Event|SIMPLE_SEGMENT|6643,6645|false|false|false|||CR
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6663,6666|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6663,6666|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6663,6666|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6663,6666|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6663,6666|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|6670,6677|false|false|false|||achieve
Finding|Idea or Concept|SIMPLE_SEGMENT|6678,6682|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|6678,6682|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6683,6686|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6683,6686|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6683,6686|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|6683,6686|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|6683,6686|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6683,6686|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6697,6705|false|false|false|C4727483|BRAF Gene Rearrangement|Positive
Finding|Classification|SIMPLE_SEGMENT|6697,6705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|SIMPLE_SEGMENT|6697,6705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Event|Event|SIMPLE_SEGMENT|6706,6707|false|false|false|||U
Finding|Body Substance|SIMPLE_SEGMENT|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6719,6731|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|6719,6731|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|SIMPLE_SEGMENT|6756,6764|false|false|false|||bacteria
Finding|Functional Concept|SIMPLE_SEGMENT|6756,6764|false|false|false|C1510439|bacteria aspects|bacteria
Finding|Finding|SIMPLE_SEGMENT|6784,6796|true|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|Asymptomatic
Event|Event|SIMPLE_SEGMENT|6806,6812|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|6806,6812|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|6813,6820|true|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|6813,6820|true|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|6821,6828|true|false|false|||malaise
Finding|Sign or Symptom|SIMPLE_SEGMENT|6821,6828|true|false|false|C0231218|Malaise|malaise
Finding|Body Substance|SIMPLE_SEGMENT|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6830,6843|false|false|false|C0430404|Urine culture|Urine culture
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6830,6852|false|false|false|C0853721|Culture urine negative|Urine culture negative
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6836,6843|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|6836,6843|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|6836,6843|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|6836,6843|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6836,6843|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6836,6852|false|false|false|C0855652|Culture negative|culture negative
Event|Event|SIMPLE_SEGMENT|6844,6852|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6844,6852|false|false|false|C5237010|Expression Negative|negative
Finding|Functional Concept|SIMPLE_SEGMENT|6857,6861|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6868,6872|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6868,6872|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6868,6872|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|6868,6872|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6868,6886|false|false|false|C0521530|Lung consolidation|lung consolidation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6873,6886|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|6873,6886|false|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|6888,6898|false|false|false|||infiltrate
Finding|Functional Concept|SIMPLE_SEGMENT|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|SIMPLE_SEGMENT|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|SIMPLE_SEGMENT|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Finding|SIMPLE_SEGMENT|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Idea or Concept|SIMPLE_SEGMENT|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Intellectual Product|SIMPLE_SEGMENT|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6903,6912|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|Radiology
Event|Event|SIMPLE_SEGMENT|6913,6917|false|false|false|||read
Finding|Conceptual Entity|SIMPLE_SEGMENT|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Intellectual Product|SIMPLE_SEGMENT|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6913,6917|false|false|false|C4723641|Nucleotide Sequence Read|read
Event|Event|SIMPLE_SEGMENT|6922,6931|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6922,6931|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|6932,6935|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6932,6935|false|false|false|C0039985|Plain chest X-ray|CXR
Drug|Organic Chemical|SIMPLE_SEGMENT|6940,6945|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6940,6945|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|6940,6945|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|6940,6945|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|6947,6953|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|6947,6953|true|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6955,6967|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|6955,6967|true|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|6955,6967|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|6969,6979|false|false|false|||Rereviewed
Finding|Functional Concept|SIMPLE_SEGMENT|6989,6993|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|6989,6993|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|6989,6993|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|6989,6993|true|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Event|Event|SIMPLE_SEGMENT|6994,7005|true|false|false|||radiologist
Finding|Intellectual Product|SIMPLE_SEGMENT|6994,7005|true|false|false|C1549438|Procedure Practitioner Identifier Code Type - Radiologist|radiologist
Event|Event|SIMPLE_SEGMENT|7010,7017|true|false|false|||favored
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7018,7027|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7018,7027|true|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7018,7027|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7018,7033|true|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7028,7033|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|7028,7033|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7028,7033|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|7043,7047|true|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|7052,7058|true|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|SIMPLE_SEGMENT|7059,7066|true|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|7059,7066|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7059,7066|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7070,7073|true|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|7070,7073|true|false|false|||PNA
Event|Event|SIMPLE_SEGMENT|7074,7083|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|7074,7083|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|7074,7083|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|7074,7083|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7074,7083|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|7103,7112|false|false|false|||indicated
Event|Event|SIMPLE_SEGMENT|7114,7123|true|false|false|||Monitored
Finding|Idea or Concept|SIMPLE_SEGMENT|7136,7147|true|false|false|C0750502|Significant|significant
Finding|Intellectual Product|SIMPLE_SEGMENT|7148,7156|true|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Finding|Sign or Symptom|SIMPLE_SEGMENT|7148,7165|true|false|false|C0037088|Signs and Symptoms|clinical findings
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7157,7165|true|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|7157,7165|true|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|7157,7165|true|false|false|C2607943|findings aspects|findings
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7170,7173|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7170,7173|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7170,7173|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|7170,7173|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|7175,7189|false|false|false|||anticoagulated
Drug|Organic Chemical|SIMPLE_SEGMENT|7193,7201|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7193,7201|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|7202,7206|false|false|false|||goal
Finding|Idea or Concept|SIMPLE_SEGMENT|7202,7206|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|7202,7206|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|SIMPLE_SEGMENT|7219,7224|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7219,7224|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7219,7224|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|7229,7237|true|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|7229,7237|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|SIMPLE_SEGMENT|7241,7245|true|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|7241,7245|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|7241,7245|true|false|false|C0582103|Medical Examination|exam
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7253,7256|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|7253,7256|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7253,7256|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7253,7256|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|SIMPLE_SEGMENT|7257,7264|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|7269,7278|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|7282,7286|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7282,7286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7282,7286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7282,7286|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7288,7296|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7288,7296|false|false|false|C0699129|Coumadin|Coumadin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7312,7318|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|7312,7318|false|false|false|||Anemia
Event|Event|SIMPLE_SEGMENT|7323,7328|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7323,7328|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7323,7328|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7332,7340|true|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|SIMPLE_SEGMENT|7332,7340|true|false|false|C0521134|External route|external
Event|Event|SIMPLE_SEGMENT|7341,7345|true|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|7341,7345|true|false|false|C5890125|Loss (adaptation)|loss
Event|Event|SIMPLE_SEGMENT|7360,7367|true|false|false|||denying
Event|Event|SIMPLE_SEGMENT|7373,7379|true|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|7373,7379|true|false|false|C0025222|Melena|melena
Event|Event|SIMPLE_SEGMENT|7393,7399|false|false|false|||anemic
Finding|Finding|SIMPLE_SEGMENT|7393,7399|false|false|false|C0857322|Anemic|anemic
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7405,7413|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|7405,7413|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7405,7413|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|7419,7428|false|false|false|||presented
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7434,7437|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7434,7437|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|7434,7437|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|7434,7437|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7434,7437|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Finding|SIMPLE_SEGMENT|7442,7448|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7442,7448|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7453,7458|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7453,7458|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7453,7466|false|false|false|C0022658|Kidney Diseases|renal disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7459,7466|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7459,7466|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7471,7474|false|false|false|C0002873;C1275685;C4554601;C5960004|Amyloidosis cutis dyschromia;Anemia of chronic disease;Angiokeratoma Corporis Diffusum;Avellino corneal dystrophy|ACD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Organic Chemical|SIMPLE_SEGMENT|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Event|Event|SIMPLE_SEGMENT|7471,7474|false|false|false|||ACD
Finding|Gene or Genome|SIMPLE_SEGMENT|7471,7474|false|false|false|C1538901|ACD gene|ACD
Finding|Finding|SIMPLE_SEGMENT|7483,7495|false|true|false|C0302845|Mean corpuscular volume above reference range|elevated MCV
Disorder|Virus|SIMPLE_SEGMENT|7492,7495|false|true|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|7492,7495|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7492,7495|false|true|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7492,7495|false|true|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7492,7495|false|true|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Event|Event|SIMPLE_SEGMENT|7497,7506|false|false|false|||indicates
Finding|Finding|SIMPLE_SEGMENT|7507,7515|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|7516,7531|false|false|false|||reticulocytosis
Finding|Finding|SIMPLE_SEGMENT|7516,7531|false|true|false|C0206160|Reticulocytosis|reticulocytosis
Finding|Finding|SIMPLE_SEGMENT|7544,7547|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|7544,7547|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|7548,7557|false|false|false|||suspicion
Finding|Mental Process|SIMPLE_SEGMENT|7548,7557|false|false|false|C0242114|Suspicion|suspicion
Event|Event|SIMPLE_SEGMENT|7563,7566|false|false|false|||GIB
Drug|Organic Chemical|SIMPLE_SEGMENT|7570,7578|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7570,7578|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|7570,7578|false|false|false|||Coumadin
Event|Event|SIMPLE_SEGMENT|7583,7592|false|false|false|||continued
Anatomy|Cell|SIMPLE_SEGMENT|7594,7607|false|false|false|C0035286|Reticulocytes|Reticulocytes
Event|Event|SIMPLE_SEGMENT|7636,7643|false|false|false|||arguing
Finding|Intellectual Product|SIMPLE_SEGMENT|7652,7657|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|7658,7662|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|7658,7662|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Cell Component|SIMPLE_SEGMENT|7678,7681|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7678,7681|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|7688,7693|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|7694,7702|false|false|false|||uprising
Event|Event|SIMPLE_SEGMENT|7706,7715|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7706,7715|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7720,7727|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|7720,7727|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7720,7727|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7720,7742|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Finding|Classification|SIMPLE_SEGMENT|7720,7749|false|false|false|C2074731|chronic kidney disease stage|Chronic kidney disease, stage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7728,7734|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7728,7734|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|7728,7734|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7728,7734|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7728,7734|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7728,7742|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7735,7742|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7735,7742|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7744,7749|false|false|false|C1300072|Tumor stage|stage
Event|Event|SIMPLE_SEGMENT|7744,7749|false|false|false|||stage
Finding|Intellectual Product|SIMPLE_SEGMENT|7744,7752|false|false|false|C0441772|Stage level 4|stage IV
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7754,7762|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|7754,7762|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7754,7762|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|SIMPLE_SEGMENT|7768,7774|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7768,7774|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7780,7783|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|7780,7783|false|false|false|||HTN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7806,7817|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7806,7817|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7806,7817|true|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7806,7817|true|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7822,7829|true|false|false|||trended
Finding|Idea or Concept|SIMPLE_SEGMENT|7842,7853|true|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|7854,7860|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|7854,7860|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7854,7860|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|7865,7868|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|7870,7879|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7880,7884|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7880,7884|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7880,7884|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7885,7897|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7885,7897|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|7885,7897|false|false|false|||atorvastatin
Event|Event|SIMPLE_SEGMENT|7909,7913|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7909,7913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7909,7913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7909,7913|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7934,7944|false|false|false|||maintained
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Hormone|SIMPLE_SEGMENT|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|7955,7958|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Event|Event|SIMPLE_SEGMENT|7955,7958|false|false|false|||ISS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Event|Event|SIMPLE_SEGMENT|7973,7976|false|false|false|||qHS
Finding|Idea or Concept|SIMPLE_SEGMENT|7982,7986|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7987,8003|false|false|false|C5392125|Glycemic Control|glycemic control
Drug|Organic Chemical|SIMPLE_SEGMENT|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|7996,8003|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|8006,8018|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8045,8048|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8045,8048|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|8045,8048|false|false|false|||CHF
Event|Event|SIMPLE_SEGMENT|8050,8058|false|false|false|||diuresed
Drug|Organic Chemical|SIMPLE_SEGMENT|8067,8072|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8067,8072|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8067,8072|false|false|false|||lasix
Event|Event|SIMPLE_SEGMENT|8074,8086|false|false|false|||transitioned
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8093,8102|false|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|8093,8102|false|false|false|||diuretics
Event|Event|SIMPLE_SEGMENT|8105,8115|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|8116,8120|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8116,8120|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8116,8120|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8116,8120|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8132,8141|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8132,8141|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|8132,8141|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|8146,8150|false|false|false|||take
Event|Event|SIMPLE_SEGMENT|8165,8169|false|false|false|||take
Procedure|Health Care Activity|SIMPLE_SEGMENT|8165,8169|false|false|false|C1515187|Take|take
Drug|Food|SIMPLE_SEGMENT|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Immunologic Factor|SIMPLE_SEGMENT|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Organic Chemical|SIMPLE_SEGMENT|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Event|Event|SIMPLE_SEGMENT|8173,8179|false|false|false|||banana
Event|Event|SIMPLE_SEGMENT|8184,8194|false|false|false|||complained
Finding|Idea or Concept|SIMPLE_SEGMENT|8217,8227|false|false|false|C1548386|Document Completion - incomplete|incomplete
Event|Event|SIMPLE_SEGMENT|8228,8235|false|false|false|||hearing
Finding|Finding|SIMPLE_SEGMENT|8228,8235|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|8228,8235|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Event|Event|SIMPLE_SEGMENT|8237,8241|true|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|8237,8241|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Idea or Concept|SIMPLE_SEGMENT|8245,8248|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8245,8248|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|8252,8261|true|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8252,8261|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8252,8261|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8252,8261|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8252,8261|true|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|8271,8275|true|false|false|||felt
Drug|Organic Chemical|SIMPLE_SEGMENT|8282,8289|true|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|8282,8289|true|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|8282,8289|true|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|8282,8289|true|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8294,8303|true|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|8294,8303|true|false|false|||diuretics
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8319,8322|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|8319,8322|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|8324,8333|false|false|false|||increased
Drug|Organic Chemical|SIMPLE_SEGMENT|8334,8344|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8334,8344|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|8334,8344|false|false|false|||nifedipine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8356,8359|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8356,8359|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8356,8359|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8356,8359|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8356,8359|false|false|false|C1332410|BID gene|BID
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8375,8379|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Event|Event|SIMPLE_SEGMENT|8389,8390|false|false|false|||f
Finding|Idea or Concept|SIMPLE_SEGMENT|8396,8400|false|false|false|C1552851|next - HtmlLinkType|next
Event|Activity|SIMPLE_SEGMENT|8401,8413|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|8401,8413|false|false|false|||appointments
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8415,8421|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|8415,8421|false|false|false|||Anemia
Event|Event|SIMPLE_SEGMENT|8438,8445|false|false|false|||workups
Event|Event|SIMPLE_SEGMENT|8446,8453|false|false|false|||showing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8454,8457|false|false|false|C0002873;C1275685;C4554601;C5960004|Amyloidosis cutis dyschromia;Anemia of chronic disease;Angiokeratoma Corporis Diffusum;Avellino corneal dystrophy|ACD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Organic Chemical|SIMPLE_SEGMENT|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Event|Event|SIMPLE_SEGMENT|8454,8457|false|false|false|||ACD
Finding|Gene or Genome|SIMPLE_SEGMENT|8454,8457|false|false|false|C1538901|ACD gene|ACD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8459,8462|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8459,8462|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|8459,8462|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|8459,8462|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8459,8462|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|SIMPLE_SEGMENT|8466,8472|false|false|false|||during
Event|Event|SIMPLE_SEGMENT|8474,8483|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8474,8483|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8490,8493|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8490,8493|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8490,8493|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|8490,8493|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|8498,8507|false|false|false|||continued
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8508,8519|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8511,8519|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|8511,8519|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8511,8519|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|8511,8519|false|false|false|||warfarin
Event|Event|SIMPLE_SEGMENT|8526,8530|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|8531,8540|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8531,8540|false|false|false|C0549178|Continuous|continued
Event|Activity|SIMPLE_SEGMENT|8542,8552|false|false|false|C1283169||monitoring
Event|Event|SIMPLE_SEGMENT|8542,8552|false|false|false|||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|8542,8552|false|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|SIMPLE_SEGMENT|8557,8564|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|8565,8569|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8565,8569|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8565,8569|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8565,8569|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|8582,8590|false|false|false|C4288901|In-House|in-house
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Hormone|SIMPLE_SEGMENT|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Event|Event|SIMPLE_SEGMENT|8603,8609|false|false|false|||aspart
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Event|Event|SIMPLE_SEGMENT|8610,8618|false|false|false|||glargine
Event|Event|SIMPLE_SEGMENT|8620,8630|false|false|false|||discharged
Finding|Idea or Concept|SIMPLE_SEGMENT|8634,8638|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8634,8638|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8634,8638|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|8639,8646|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|8639,8646|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8639,8646|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Body Substance|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8648,8657|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8658,8664|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|8658,8664|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|8658,8664|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|8658,8664|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|8658,8664|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8671,8680|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8691,8702|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8691,8702|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8691,8702|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8691,8702|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8691,8715|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8706,8715|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8706,8715|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8734,8744|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8734,8744|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8734,8749|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8745,8749|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8745,8749|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8753,8761|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|8766,8774|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|8766,8774|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8766,8774|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8779,8792|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8779,8792|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8779,8792|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8779,8792|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|8811,8814|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8815,8819|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8815,8819|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8815,8819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8815,8819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|8823,8828|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|8823,8828|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|8823,8828|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|SIMPLE_SEGMENT|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8860,8872|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8860,8872|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|8882,8885|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|8890,8900|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8890,8900|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8912,8915|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8912,8915|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8912,8915|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8912,8915|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8912,8915|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8920,8928|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8920,8928|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|8920,8928|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|8920,8935|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8920,8935|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|8929,8935|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8929,8935|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8929,8935|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8946,8949|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8946,8949|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8946,8949|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8946,8949|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8946,8949|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8954,8964|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8954,8964|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|SIMPLE_SEGMENT|8979,8995|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8979,8995|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8991,8995|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8991,8995|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8991,8995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8991,8995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9000,9010|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9000,9010|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|9030,9043|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9046,9049|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9046,9049|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|9063,9073|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9063,9073|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|SIMPLE_SEGMENT|9063,9073|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9086,9089|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9086,9089|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9086,9089|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9086,9089|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9086,9089|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9095,9108|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9095,9108|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|9095,9108|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|9128,9131|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9132,9137|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9132,9137|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9132,9142|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9132,9142|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9138,9142|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9138,9142|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9138,9142|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9138,9142|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9148,9160|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9148,9160|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9180,9192|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|9180,9192|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|9180,9192|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|9180,9199|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9180,9199|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9193,9199|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|9193,9199|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|SIMPLE_SEGMENT|9193,9199|false|false|false|||Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|9219,9224|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9219,9224|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9235,9238|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9235,9238|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9235,9238|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9235,9238|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9235,9238|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|9239,9251|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9239,9251|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9257,9266|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9265,9266|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|9271,9275|false|false|false|||UNIT
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9320,9331|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9320,9331|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|SIMPLE_SEGMENT|9354,9357|false|false|false|||DAY
Finding|Idea or Concept|SIMPLE_SEGMENT|9354,9357|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|SIMPLE_SEGMENT|9354,9357|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|SIMPLE_SEGMENT|9363,9372|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9363,9372|false|false|false|C0076840|torsemide|Torsemide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|SIMPLE_SEGMENT|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|SIMPLE_SEGMENT|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9408,9415|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9408,9415|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9408,9415|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|SIMPLE_SEGMENT|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9416,9419|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9416,9419|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|SIMPLE_SEGMENT|9416,9419|false|false|false|||NPH
Event|Event|SIMPLE_SEGMENT|9460,9472|false|false|false|||subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|9460,9472|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Event|Event|SIMPLE_SEGMENT|9487,9493|false|false|false|||dinner
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9487,9493|false|false|false|C4048877|Dinner|dinner
Event|Event|SIMPLE_SEGMENT|9498,9507|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9498,9507|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9498,9519|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9508,9519|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9508,9519|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9508,9519|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9508,9519|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|SIMPLE_SEGMENT|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Event|Event|SIMPLE_SEGMENT|9524,9531|false|false|false|||HumuLIN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|SIMPLE_SEGMENT|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9539,9546|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9539,9546|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9539,9546|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|SIMPLE_SEGMENT|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9547,9550|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9547,9550|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|SIMPLE_SEGMENT|9547,9550|false|false|false|||NPH
Event|Event|SIMPLE_SEGMENT|9591,9603|false|false|false|||subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|9591,9603|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Event|Event|SIMPLE_SEGMENT|9618,9624|false|false|false|||dinner
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9618,9624|false|false|false|C4048877|Dinner|dinner
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9658,9667|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9666,9667|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|9672,9676|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|9690,9703|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9690,9703|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|9690,9703|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9690,9703|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|9722,9725|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9726,9730|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9726,9730|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9726,9730|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9726,9730|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9734,9739|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|9734,9739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9734,9739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|SIMPLE_SEGMENT|9744,9755|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9744,9755|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|SIMPLE_SEGMENT|9778,9781|false|false|false|||DAY
Finding|Idea or Concept|SIMPLE_SEGMENT|9778,9781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|SIMPLE_SEGMENT|9778,9781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|SIMPLE_SEGMENT|9786,9793|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9786,9793|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9813,9825|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9813,9825|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|9835,9838|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|9843,9851|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9843,9851|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|9843,9851|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|9843,9858|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9843,9858|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|9852,9858|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|9852,9858|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9852,9858|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9869,9872|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9869,9872|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9869,9872|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9869,9872|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9869,9872|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9877,9887|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9877,9887|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|SIMPLE_SEGMENT|9902,9918|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9902,9918|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9914,9918|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9914,9918|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9914,9918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9914,9918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9924,9934|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9924,9934|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|9955,9968|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9971,9974|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9971,9974|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|9989,10002|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9989,10002|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|9989,10002|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|10022,10025|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10026,10031|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|10026,10031|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10026,10036|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10026,10036|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10032,10036|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10032,10036|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10032,10036|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10032,10036|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10042,10054|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10042,10054|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|10042,10054|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|10042,10061|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10042,10061|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10055,10061|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|10055,10061|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|10081,10086|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10081,10086|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10097,10100|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10097,10100|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10097,10100|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10097,10100|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10097,10100|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|10101,10113|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|10101,10113|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|10119,10128|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10119,10128|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|SIMPLE_SEGMENT|10149,10158|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10149,10158|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|10149,10158|false|false|false|||torsemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10167,10173|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10177,10185|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|10186,10190|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10208,10214|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10215,10222|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10215,10222|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|10230,10242|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10230,10242|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|10262,10272|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10262,10272|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10282,10285|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10282,10285|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10282,10285|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10282,10285|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10282,10285|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10291,10301|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10291,10301|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|SIMPLE_SEGMENT|10291,10301|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10314,10317|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10314,10317|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10314,10317|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|10314,10317|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|10314,10317|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|10323,10333|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10323,10333|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|10323,10333|false|false|false|||nifedipine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10342,10349|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10342,10349|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10342,10349|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|10353,10361|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10356,10361|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10356,10361|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|10374,10378|false|false|false|||Disp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10386,10393|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|10386,10393|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10386,10393|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|10394,10401|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10394,10401|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|10408,10417|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10408,10417|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10408,10429|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10408,10429|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10418,10429|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10418,10429|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10418,10429|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|10431,10435|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|10431,10435|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|10431,10435|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10431,10435|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|10441,10448|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|10441,10448|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|10451,10459|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|10451,10459|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|10467,10476|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10467,10476|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10467,10486|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10477,10486|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10477,10486|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10477,10486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10477,10486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10477,10486|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|10496,10505|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10496,10505|false|false|false|C0011900|Diagnosis|Diagnoses
Finding|Intellectual Product|SIMPLE_SEGMENT|10507,10512|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|SIMPLE_SEGMENT|10516,10523|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10516,10523|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10538,10562|false|false|false|C0018802|Congestive heart failure|congestive Heart Failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10549,10554|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10549,10554|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|10549,10554|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10549,10562|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|Heart Failure
Event|Event|SIMPLE_SEGMENT|10555,10562|false|false|false|||Failure
Finding|Functional Concept|SIMPLE_SEGMENT|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10563,10575|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|10563,10575|false|false|false|||Hypertension
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10577,10586|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|10577,10586|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|10577,10586|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|SIMPLE_SEGMENT|10587,10596|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10587,10596|false|false|false|C0011900|Diagnosis|Diagnoses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10598,10604|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|10598,10604|false|false|false|||Anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10605,10613|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10605,10622|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Event|Event|SIMPLE_SEGMENT|10614,10622|false|false|false|||mellitus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10629,10633|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10629,10638|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10629,10649|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10634,10638|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|10634,10649|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|10639,10649|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|10639,10649|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Intellectual Product|SIMPLE_SEGMENT|10650,10657|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|10650,10657|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10650,10672|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10658,10664|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10658,10664|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Event|Event|SIMPLE_SEGMENT|10658,10664|false|false|false|||Kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|10658,10664|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10658,10664|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10658,10664|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10658,10672|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10665,10672|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|10665,10672|false|false|false|||Disease
Event|Event|SIMPLE_SEGMENT|10676,10685|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10676,10685|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10676,10685|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10676,10685|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10676,10685|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10686,10695|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10686,10695|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10686,10695|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10686,10695|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10697,10703|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10697,10710|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10697,10710|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10704,10710|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10704,10710|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10712,10717|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10712,10717|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10722,10730|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10722,10730|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10732,10737|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10732,10754|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10732,10754|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10741,10754|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10741,10754|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10741,10754|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10756,10761|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10756,10761|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10756,10761|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10756,10761|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10766,10777|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10766,10777|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10779,10787|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10779,10787|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10779,10787|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10788,10794|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10788,10794|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10788,10794|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10796,10806|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|10796,10806|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|10809,10820|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|10809,10820|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|10809,10820|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|10825,10834|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10825,10834|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10825,10834|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10825,10834|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10825,10834|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10825,10847|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10825,10847|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|10825,10847|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10835,10847|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10835,10847|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10835,10847|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|10870,10878|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|10890,10899|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10890,10899|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10890,10899|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10890,10899|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10890,10899|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|10908,10918|false|false|false|||congestive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10920,10925|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10920,10925|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|10920,10925|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10920,10933|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|10926,10933|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10938,10950|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|10938,10950|false|false|false|||hypertension
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10970,10979|false|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|10970,10979|false|false|false|||diuretics
Event|Event|SIMPLE_SEGMENT|10986,10997|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|10986,10997|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|11006,11014|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|11006,11014|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|11006,11014|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|11016,11020|false|false|false|||labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11016,11020|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|11025,11029|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|11025,11029|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|11025,11029|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|11034,11043|false|false|false|||increased
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11057,11062|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|11057,11062|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|11057,11062|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|11057,11071|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|11057,11071|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|11057,11071|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|11063,11071|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11063,11071|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11072,11083|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11072,11083|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|11072,11083|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11072,11083|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|11088,11097|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|11109,11113|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11109,11113|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11109,11113|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11109,11113|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11115,11124|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|SIMPLE_SEGMENT|11115,11124|false|false|false|||medicines
Event|Event|SIMPLE_SEGMENT|11137,11145|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11137,11145|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11137,11145|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11153,11157|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11153,11157|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11153,11157|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11153,11157|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11153,11160|false|false|false|C1555558|care of - AddressPartType|care of
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11186,11190|false|false|false|C3273412|NCK-Interacting Protein with SH3 Domain|wish
Event|Event|SIMPLE_SEGMENT|11186,11190|false|false|false|||wish
Finding|Gene or Genome|SIMPLE_SEGMENT|11186,11190|false|false|false|C1423524;C3273411|NCKIPSD gene;NCKIPSD wt Allele|wish
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11204,11208|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|11204,11208|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|11204,11208|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|11229,11237|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11238,11250|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11238,11250|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11238,11250|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

