CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Hypertensive disease|Disorder|false|false||HTNnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Fever|Finding|false|false||feversnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Usual|Modifier|false|false||usualnull|personal health|Finding|false|false||state of healthnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Health|Finding|false|false||healthnull|Evening|Time|false|false||eveningnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Robitussin|Drug|false|false||robitussin
null|Robitussin|Drug|false|false||robitussinnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Morning|Time|false|false||morningnull|Malaise|Finding|false|false||general malaisenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||generalnull|General medical service|Procedure|false|false||generalnull|Generalized|Modifier|false|false||generalnull|Malaise|Finding|false|false||malaisenull|Nasal congestion (finding)|Finding|false|false|C0028429|nasal congestionnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C0027424;C4520890;C1522019;C1272939;C0721966|nasalnull|Congestion|Finding|false|false||congestionnull|Productive Cough|Finding|false|false||productive coughnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Episode of|Time|false|false||episodesnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Vomiting|Finding|false|false||vomitingnull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Fever|Finding|true|false||feversnull|Chills|Finding|false|false||chillsnull|Sweating|Finding|true|false||sweats
null|Sweat|Finding|true|false||sweatsnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Pack|Drug|false|false||packnull|Pack (physical object)|Device|false|false||pack
null|Pack unit|Device|false|false||packnull|Packing (action)|Event|false|false||packnull|Package Dosing Unit|LabModifier|false|false||packnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Coughing|Finding|false|false||coughingnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Abdomen|Anatomy|false|false|C2003888;C0941288;C0741025;C0153662|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726;C0000726;C0446470|abdomennull|Abdomen problem|Finding|false|false|C0000726;C0446470;C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288;C0741025|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288;C0741025|abdomennull|Surface region of lower chest|Anatomy|false|false|C0741025;C0941288;C0153662;C2003888|lower chestnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C0741025|lowernull|Lower (action)|Event|false|false|C0000726;C1548802;C0446470|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Chest problem|Finding|false|false|C1527391;C0817096;C0446470;C0000726;C0230168;C0000726;C1548802|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417|jointnull|null|Anatomy|false|false|C0575044;C0231528|joint
null|Joints|Anatomy|false|false|C0575044;C0231528|joint
null|Articular system|Anatomy|false|false|C0575044;C0231528|jointnull|Joint Device|Device|false|false||jointnull|Myalgia|Finding|false|false|C4083049;C0026845;C0392905;C1269611;C0022417|muscle painnull|Muscle (organ)|Anatomy|false|false|C1549543;C0030193;C0231528|muscle
null|Muscle Tissue|Anatomy|false|false|C1549543;C0030193;C0231528|musclenull|Administration Method - Pain|Finding|false|false|C4083049;C0026845|pain
null|Pain|Finding|false|false|C4083049;C0026845|painnull|null|Attribute|false|false||painnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Hypoxia|Finding|false|false||hypoxicnull|Influenza virus vaccine|Drug|false|false||flu vaccine
null|Influenza virus vaccine|Drug|false|false||flu vaccinenull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|Vaccine [APC]|Drug|false|false||vaccine
null|Vaccines|Drug|false|false||vaccine
null|Vaccines|Drug|false|false||vaccine
null|Vaccines|Drug|false|false||vaccinenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Pneumovax|Drug|false|false||pneumovax
null|Pneumovax|Drug|false|false||pneumovaxnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Wheezing|Finding|false|false||wheezynull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Apyrexial|Finding|false|false||afebrilenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Wheezing|Finding|false|false||wheezesnull|Peak flow|Finding|false|false||peak flownull|Peak level|Modifier|false|false||peaknull|Flow|Phenomenon|false|false||flownull|BaseLine dental cement|Drug|true|false||baselinenull|baseline - TableCellVerticalAlign|Finding|true|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Full|Modifier|false|false||fullnull|Sentence|Finding|false|false||sentencesnull|Use of accessory muscles|Finding|true|false|C4083049;C0026845|accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false|C4083049;C0026845|accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false|C1947944;C0042153;C0457083;C0158784;C1821466|muscle
null|Muscle Tissue|Anatomy|false|false|C1947944;C0042153;C0457083;C0158784;C1821466|musclenull|Use - dosing instruction imperative|Finding|false|false|C4083049;C0026845|use
null|utilization qualifier|Finding|false|false|C4083049;C0026845|use
null|Usage|Finding|false|false|C4083049;C0026845|usenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Influenza|Disorder|false|false||Flunull|ZMYND10 wt Allele|Finding|false|false||Flunull|Fluorescence Units|LabModifier|false|false||Flunull|Toxicology screen, general (procedure)|Procedure|false|false||screen
null|Disease Screening|Procedure|false|false||screen
null|Screening for cancer|Procedure|false|false||screen
null|Screening procedure|Procedure|false|false||screennull|Screen Device|Device|false|false||screennull|Plain chest X-ray|Procedure|false|false||CXRnull|null|Modifier|false|false||unremarkablenull|null|Time|false|false||priornull|Nebulizer solution|Drug|false|false||nebsnull|prednylidene|Drug|false|false||pred
null|prednisone|Drug|false|false||pred
null|prednisone|Drug|false|false||pred
null|prednisone|Drug|false|false||pred
null|prednylidene|Drug|false|false||prednull|Asthma|Disorder|false|false||ASTHMAnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Headache|Finding|false|false||HEADACHEnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Atypical chest pain|Finding|false|false|C1527391;C0817096|ATYPICAL CHEST PAINnull|atypia morphology|Finding|false|false|C1527391;C0817096|ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Chest Pain|Finding|false|false|C1527391;C0817096|CHEST PAINnull|null|Attribute|false|false|C1527391;C0817096|CHEST PAINnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C2598155;C0741302;C1549543;C0030193;C0741025;C0262384;C0008031;C2926613|CHEST
null|Anterior thoracic region|Anatomy|false|false|C2598155;C0741302;C1549543;C0030193;C0741025;C0262384;C0008031;C2926613|CHESTnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|PAIN
null|Pain|Finding|false|false|C1527391;C0817096|PAINnull|null|Attribute|false|false|C1527391;C0817096|PAINnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Standard chest X-ray abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL CHEST XRAYnull|chest abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL CHESTnull|Observation Interpretation - Abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL
null|Abnormal|Finding|false|false|C1527391;C0817096|ABNORMALnull|Plain chest X-ray|Procedure|false|false|C1527391;C0817096|CHEST XRAYnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0741025;C0436503;C1550458;C0205161;C0043309;C0043299;C0742257;C0039985|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0436503;C1550458;C0205161;C0043309;C0043299;C0742257;C0039985|CHESTnull|Diagnostic radiologic examination|Procedure|false|false|C1527391;C0817096|XRAYnull|Roentgen Rays|Phenomenon|false|false|C1527391;C0817096|XRAYnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|On admission|Time|false|false||On Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429;C1550232|nasal
null|Nasal (intended site)|Finding|false|false|C0028429;C1550232|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966;C1550622;C1546577|nasalnull|Specimen Type - Cannula|Finding|false|false|C1550232;C0028429|cannula
null|null|Finding|false|false|C1550232;C0028429|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577;C4520890;C1522019|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Respiratory distress|Finding|true|false||respiratory distressnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Supple neck|Finding|false|false|C0027530;C3159206|neck supplenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C2230237;C0332254|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C2230237;C0332254|necknull|Supple|Finding|false|false|C0027530;C3159206|supplenull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Pulmonary ventilator management|Procedure|false|false||Pulmnull|cetrimonium bromide|Drug|false|false||CTABnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Inspiration (function)|Finding|false|false||inspiratorynull|Exertion|Finding|false|false||effortnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Prolonged|Time|false|false||prolongednull|Expiration, Respiratory|Finding|false|false||expiratorynull|Phase|Time|false|false||phasenull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Neg - answer|Finding|false|false||negnull|Negative - qualifier|Modifier|false|false||negnull|LRRC4B gene|Finding|false|false||HSMnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|PDSS1 gene|Finding|false|false||DPsnull|Disintegration per Second|LabModifier|false|false||DPsnull|PTS protein, human|Drug|false|false||PTs
null|4-toluenesulfonamide|Drug|false|false||PTs
null|4-toluenesulfonamide|Drug|false|false||PTs
null|PTS protein, human|Drug|false|false||PTsnull|PTS gene|Finding|false|false||PTs
null|Patient Tracking System|Finding|false|false||PTsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skinnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|Central Nervous System|Anatomy|false|false||CNsnull|Clinical Nurse Specialists|Subject|false|false||CNsnull|Certified Nurse Specialist|Title|false|false||CNsnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||CNsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C1550232;C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C1550232;C0028429|nasalnull|null|Anatomy|false|false|C1550622;C1546577;C1272939;C0721966;C4520890;C1522019|nasalnull|Specimen Type - Cannula|Finding|false|false|C0028429;C1550232|cannula
null|null|Finding|false|false|C0028429;C1550232|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577;C4520890;C1522019|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Respiratory distress|Finding|true|false||respiratory distressnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Supple neck|Finding|false|false|C0027530;C3159206|neck supplenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C2230237;C0812434;C0684335;C0332254|neck
null|Neck|Anatomy|false|false|C2230237;C0812434;C0684335;C0332254|necknull|Supple|Finding|false|false|C0027530;C3159206|supplenull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Pulmonary ventilator management|Procedure|false|false||Pulmnull|cetrimonium bromide|Drug|false|false||CTABnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Inspiration (function)|Finding|false|false||inspiratorynull|Exertion|Finding|false|false||effortnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Prolonged|Time|false|false||prolongednull|Expiration, Respiratory|Finding|false|false||expiratorynull|Phase|Time|false|false||phasenull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Neg - answer|Finding|false|false||negnull|Negative - qualifier|Modifier|false|false||negnull|LRRC4B gene|Finding|false|false||HSMnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|PDSS1 gene|Finding|false|false||DPsnull|Disintegration per Second|LabModifier|false|false||DPsnull|PTS protein, human|Drug|false|false||PTs
null|4-toluenesulfonamide|Drug|false|false||PTs
null|4-toluenesulfonamide|Drug|false|false||PTs
null|PTS protein, human|Drug|false|false||PTsnull|PTS gene|Finding|false|false||PTs
null|Patient Tracking System|Finding|false|false||PTsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skinnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|Central Nervous System|Anatomy|false|false||CNsnull|Clinical Nurse Specialists|Subject|false|false||CNsnull|Certified Nurse Specialist|Title|false|false||CNsnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||CNsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right lateral incisor mesial prosthesis|Device|false|false||26PMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right lateral incisor mesial prosthesis|Device|false|false||26PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Micro (prefix)|Finding|false|false||MICRO
null|Microbiology - Laboratory Class|Finding|false|false||MICROnull|Microbiology procedure|Procedure|false|false||MICROnull|Unit Of Measure Prefix - micro|LabModifier|false|false||MICROnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Direct - PostalAddressUse|Finding|false|false||DIRECT
null|direct address|Finding|false|false||DIRECTnull|Direct type of relationship|Modifier|false|false||DIRECT
null|Direct (qualifier)|Modifier|false|false||DIRECTnull|influenza A|Disorder|false|false||INFLUENZA Anull|Influenza virus vaccine|Drug|false|false||INFLUENZA
null|Influenza virus vaccine|Drug|false|false||INFLUENZAnull|Influenza|Disorder|false|false||INFLUENZAnull|Blood group antigen A|Drug|false|false||A ANTIGENnull|Antigen test|Procedure|false|false|C4318744|ANTIGEN TESTnull|Antigens|Drug|false|false||ANTIGENnull|Tests (qualifier value)|Finding|false|false|C4318744|TEST
null|Testing|Finding|false|false|C4318744|TESTnull|Laboratory Procedures|Procedure|false|false|C4318744|TESTnull|Test - temporal region|Anatomy|false|false|C0456984;C1546485;C0022885;C0729856;C0039593;C0392366|TESTnull|Test Result|Lab|false|false|C4318744|TESTnull|Test Dosing Unit|LabModifier|false|false||TESTnull|Diagnosis Type - Final|Finding|false|false|C4318744|Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Positive|Finding|false|false||POSITIVE FORnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|influenza A|Disorder|false|false||INFLUENZA Anull|Influenza virus vaccine|Drug|false|false||INFLUENZA
null|Influenza virus vaccine|Drug|false|false||INFLUENZAnull|Influenza|Disorder|false|false||INFLUENZAnull|Antigens, Viral|Drug|false|false||VIRAL ANTIGENnull|Viral|Finding|false|false||VIRALnull|Antigens|Drug|false|false||ANTIGENnull|Authorization Mode - Phone|Finding|false|false||PHONE
null|Visit User Code - Phone|Finding|false|false||PHONE
null|Telephone Number|Finding|false|false||PHONE
null|MDFAttributeType - Phone|Finding|false|false||PHONEnull|Telephone|Device|false|false||PHONEnull|Person location type - Phone|Modifier|false|false||PHONEnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|CHEST PATHOLOGY|Disorder|true|false|C1527391;C0817096|chest pathologynull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0919386;C0742323;C0741025;C0205469;C0677042|chest
null|Anterior thoracic region|Anatomy|false|false|C0919386;C0742323;C0741025;C0205469;C0677042|chestnull|Pathology processes|Finding|false|false|C1527391;C0817096|pathology
null|Pathological aspects|Finding|false|false|C1527391;C0817096|pathologynull|Pathology procedure|Procedure|false|false|C1527391;C0817096|pathologynull|Pathology|Title|false|false||pathologynull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0032226|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Scar Tissue|Finding|false|false||scar
null|Cicatrix|Finding|false|false||scar
null|RPS4X gene|Finding|false|false||scarnull|Flattened|Finding|false|false|C1269845|Flatteningnull|Structure of hemidiaphragm|Anatomy|false|false|C0016203;C0332290|hemidiaphragmsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C1269845|consistentnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Recent|Time|false|false||recentnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Fever|Finding|false|false||feversnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Pleuritic pain|Finding|false|false||pleuritic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|influenza A|Disorder|false|false||influenza Anull|Influenza virus vaccine|Drug|false|false||influenza
null|Influenza virus vaccine|Drug|false|false||influenzanull|Influenza|Disorder|false|false||influenzanull|Fever|Finding|false|false||Feversnull|Malaise|Finding|false|false||malaisenull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Virus Diseases|Disorder|false|false||viral infectionnull|Viral|Finding|false|false||viralnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Respiratory secretion precautions|Procedure|false|false||droplet precautionsnull|Precaution|Finding|false|false||precautionsnull|Concern|Finding|false|false||concernnull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|oseltamivir|Drug|false|false||Oseltamivir
null|oseltamivir|Drug|false|false||Oseltamivirnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Nasopharyngeal swab (specimen)|Finding|false|false|C0027442|nasopharyngeal swabnull|nasopharyngeal swab (lab test)|Procedure|false|false|C0027442|nasopharyngeal swab
null|Nasal Swab Test|Procedure|false|false|C0027442|nasopharyngeal swabnull|Nasopharyngeal swab (physical object)|Device|false|false||nasopharyngeal swabnull|Nasopharynx|Anatomy|false|false|C0444192;C0563454;C4318939;C2266655|nasopharyngealnull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false|C0027442|swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Influenza virus vaccine|Drug|false|false||influenza
null|Influenza virus vaccine|Drug|false|false||influenzanull|Influenza|Disorder|false|false||influenzanull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|oseltamivir|Drug|false|false||oseltamivir
null|oseltamivir|Drug|false|false||oseltamivirnull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Sputum production|Finding|false|false||sputum productionnull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Production Processing ID|Finding|false|false||productionnull|production|Event|false|false||productionnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Daily|Time|false|false||Dailynull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycinnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429;C1550232|nasal
null|Nasal (intended site)|Finding|false|false|C0028429;C1550232|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966;C1550622;C1546577|nasalnull|Specimen Type - Cannula|Finding|false|false|C0028429;C1550232|cannula
null|null|Finding|false|false|C0028429;C1550232|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577;C4520890;C1522019|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Rest|Finding|false|false||restingnull|Initially|Time|false|false||initiallynull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Daily|Time|false|false||Dailynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|null|Procedure|false|false||tapernull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|More|LabModifier|false|false||morenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Asthma|Disorder|false|false||ASTHMAnull|Wheezing|Finding|false|false||wheezingnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Asthma|Disorder|false|false||asthmanull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizernull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Respiratory Status|Finding|false|false||Respiratory statusnull|null|Attribute|false|false||Respiratory statusnull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Hypertensive (finding)|Finding|false|false||hypertensivenull|Continuous|Finding|false|false||continuenull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Morning|Time|false|false||in the morningnull|Morning|Time|false|false||morningnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Every twenty four hours|Time|false|false||Q24Hnull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|Daily|Time|false|false||DAILYnull|Imdur|Drug|false|false||IMDUR
null|Imdur|Drug|false|false||IMDURnull|Daily|Time|false|false||DAILYnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Current (present time)|Time|false|false||Currentlynull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Daily|Time|false|false||Dailynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Recent|Time|false|false||recentlynull|Single vessel disease|Disorder|false|false||single vessel diseasenull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Daily|Time|false|false||DAILYnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|year|Time|false|false||yearsnull|Patient need for (contextual qualifier)|Finding|false|false||need fornull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|Nicotine Transdermal Patch|Drug|false|false||nicotine patchnull|nicotine|Drug|false|false||nicotine
null|nicotine|Drug|false|false||nicotinenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Gum as an ingredient|Drug|false|false|C0017562|gum
null|Gum Dose Form|Drug|false|false|C0017562|gumnull|OTULIN wt Allele|Finding|false|false|C0017562|gum
null|OTULIN gene|Finding|false|false|C0017562|gumnull|Gingiva|Anatomy|false|false|C0812395;C1378701;C5444202;C1825233|gumnull|Gum - unit of product usage|LabModifier|false|false||gum
null|Gum Dosing Unit|LabModifier|false|false||gumnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||Dailynull|B-Complex|Drug|false|false||B complex
null|B-Complex|Drug|false|false||B complex
null|B-Complex|Drug|false|false||B complexnull|complex (molecular entity)|Drug|false|false||complexnull|Complex|Modifier|false|false||complexnull|Vitamin C Drug Class|Drug|false|false||vitamin C
null|ascorbic acid|Drug|false|false||vitamin C
null|ascorbic acid|Drug|false|false||vitamin C
null|ascorbic acid|Drug|false|false||vitamin C
null|Vitamin C Vitamins|Drug|false|false||vitamin C
null|Vitamin C Vitamins|Drug|false|false||vitamin C
null|Vitamin C [EPC]|Drug|false|false||vitamin C
null|Vitamin C Drug Class|Drug|false|false||vitamin Cnull|Ascorbic acid measurement|Procedure|false|false||vitamin Cnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acidnull|Folic acid measurement|Procedure|false|false||folic acidnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|cinacalcet|Drug|false|false||cinacalcet
null|cinacalcet|Drug|false|false||cinacalcetnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|metoprolol succinate|Drug|false|false||metoprolol succinate
null|metoprolol succinate|Drug|false|false||metoprolol succinatenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|succinate|Drug|false|false||succinate
null|Succinates|Drug|false|false||succinatenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|doxazosin|Drug|false|false||doxazosin
null|doxazosin|Drug|false|false||doxazosinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|sevelamer hydrochloride|Drug|false|false||sevelamer HCl
null|sevelamer hydrochloride|Drug|false|false||sevelamer HClnull|sevelamer|Drug|false|false||sevelamer
null|sevelamer|Drug|false|false||sevelamernull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Meal (occasion for eating)|Finding|false|false||MEALSnull|With meals|Time|false|false||MEALSnull|3 times|Finding|false|false||3 TIMESnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||TIMESnull|Time|Time|false|false||TIMESnull|Times|LabModifier|false|false||TIMESnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|With meals|Time|false|false||WITH MEALSnull|Meal (occasion for eating)|Finding|false|false||MEALSnull|With meals|Time|false|false||MEALSnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|clonazepam|Drug|false|false||clonazepam
null|clonazepam|Drug|false|false||clonazepamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|Inhalers, Aerosol|Device|false|false||Aerosol Inhalernull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Hour|Time|false|false||hoursnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every twenty four hours|Time|false|false||Q24Hnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|24 Hours|Time|false|false||24 hoursnull|Hour|Time|false|false||hoursnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1332410;C4546282|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1332410;C4546282|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0524463;C1325531|BIDnull|BID gene|Finding|false|false|C0524463;C1325531|BIDnull|Twice a day|Time|false|false||BIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabnull|Tablet Dosing Unit|LabModifier|false|false||tabnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|diltiazem hydrochloride|Drug|false|false||diltiazem HCl
null|diltiazem hydrochloride|Drug|false|false||diltiazem HClnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false|C0524463;C1325531|HClnull|Extended Release Oral Capsule|Drug|false|false|C0524463;C1325531|Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0231448;C5781021;C0023443;C0991505;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0231448;C5781021;C0023443;C0991505;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false|C0524463;C1325531|Extended
null|Extension|Finding|false|false|C0524463;C1325531|Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Extended Release Oral Capsule|Drug|false|false|C0524463;C1325531|Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C0231448;C5781021;C1283071;C0391871;C0006935;C0991505|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C0231448;C5781021;C1283071;C0391871;C0006935;C0991505|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false|C0524463;C1325531|Extended
null|Extension|Finding|false|false|C0524463;C1325531|Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false|C0028429|Spraynull|Spray (action)|Event|false|false|C0028429|Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C2003858;C4521772;C4520890;C1522019;C1272939;C0721966|Nasalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C1550509;C0993608;C0034789|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329;C1556138|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C4035627;C4546282;C0993608;C0004048;C0205535;C1550509;C1561538;C1561539;C1332410|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false|C1556138|Inhalation
null|Inspiration (function)|Finding|false|false|C1556138|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C1556138|BIDnull|BID gene|Finding|false|false|C1556138|BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false|C1556138|2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false|C1556138|day
null|Precision - day|Finding|false|false|C1556138|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|hydrochlorothiazide|Drug|false|false||hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||hydrochlorothiazidenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|isosorbide mononitrate|Drug|false|false||isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||isosorbide mononitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|montelukast|Drug|false|false||montelukast
null|montelukast|Drug|false|false||montelukastnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|tiotropium bromide|Drug|false|false||tiotropium bromide
null|tiotropium bromide|Drug|false|false||tiotropium bromidenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false|C0524463;C1325531|bromidenull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C0202341;C0004048;C0205535|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C0202341;C0004048;C0205535|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Inhalation Devices|Device|false|false||Inhalation Devicenull|Inhalation Route of Administration|Finding|false|false|C0524463;C1325531|Inhalation
null|Inspiration (function)|Finding|false|false|C0524463;C1325531|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|calcium carbonate|Drug|false|false||calcium carbonate
null|calcium carbonate|Drug|false|false||calcium carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|carbonate ion|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonatenull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Multivitamin tablet|Drug|false|false||multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|oxygen|Drug|false|false||Oxygen
null|oxygen|Drug|false|false||Oxygen
null|oxygen|Drug|false|false||Oxygennull|Oxygen Therapy Care|Procedure|false|false||Oxygennull|Oxygen Equipment Location|Modifier|false|false||Oxygennull|Home oxygen supply|Finding|false|false||Home Oxygennull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|oxygen|Drug|false|false||Oxygen
null|oxygen|Drug|false|false||Oxygen
null|oxygen|Drug|false|false||Oxygennull|Oxygen Therapy Care|Procedure|false|false||Oxygennull|Oxygen Equipment Location|Modifier|false|false||Oxygennull|Continuous|Finding|false|false||Continuousnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429;C1550232|nasal
null|Nasal (intended site)|Finding|false|false|C0028429;C1550232|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966|nasalnull|Specimen Type - Cannula|Finding|false|false|C1550232|cannula
null|null|Finding|false|false|C1550232|cannulanull|Body Parts - Cannula|Anatomy|false|false|C1550622;C1546577;C4520890;C1522019|cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|Participation Type - device|Finding|false|false||devicenull|Medical Devices|Device|false|false||device
null|Devices|Device|false|false||devicenull|Kind of quantity - Device|LabModifier|false|false||devicenull|portability|Modifier|false|false||portabilitynull|Physiologic pulse|Finding|false|false||Pulsenull|Pulse taking|Procedure|false|false||Pulsenull|Pulse Rate|Attribute|false|false||Pulsenull|Pulse phenomenon|Phenomenon|false|false||Pulsenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|portability|Modifier|false|false||portabilitynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Influenza virus vaccine|Drug|false|false||Influenza
null|Influenza virus vaccine|Drug|false|false||Influenzanull|Influenza|Disorder|false|false||Influenzanull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|Secondary diagnosis|Finding|false|false||Secondary Diagnosisnull|null|Attribute|false|false||Secondary Diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Asthma|Disorder|false|false||ASTHMAnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Headache|Finding|false|false||HEADACHEnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Atypical chest pain|Finding|false|false|C1527391;C0817096|ATYPICAL CHEST PAINnull|atypia morphology|Finding|false|false|C1527391;C0817096|ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Chest Pain|Finding|false|false|C1527391;C0817096|CHEST PAINnull|null|Attribute|false|false|C1527391;C0817096|CHEST PAINnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C1549543;C0030193;C0262384;C0008031;C0741302;C2926613;C2598155;C0741025|CHEST
null|Anterior thoracic region|Anatomy|false|false|C1549543;C0030193;C0262384;C0008031;C0741302;C2926613;C2598155;C0741025|CHESTnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|PAIN
null|Pain|Finding|false|false|C1527391;C0817096|PAINnull|null|Attribute|false|false|C1527391;C0817096|PAINnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Standard chest X-ray abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL CHEST XRAYnull|chest abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL CHESTnull|Observation Interpretation - Abnormal|Finding|false|false|C1527391;C0817096|ABNORMAL
null|Abnormal|Finding|false|false|C1527391;C0817096|ABNORMALnull|Plain chest X-ray|Procedure|false|false|C1527391;C0817096|CHEST XRAYnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0043299;C0436503;C0039985;C0043309;C0742257;C0741025;C1550458;C0205161|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0043299;C0436503;C0039985;C0043309;C0742257;C0741025;C1550458;C0205161|CHESTnull|Diagnostic radiologic examination|Procedure|false|false|C1527391;C0817096|XRAYnull|Roentgen Rays|Phenomenon|false|false|C1527391;C0817096|XRAYnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Similarity|Modifier|false|false||similarnull|Common Cold|Disorder|false|false||common coldnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||cold
null|Cold brand of chlorpheniramine-phenylpropanolamine|Drug|false|false||coldnull|Common Cold|Disorder|false|false||cold
null|Chronic Obstructive Airway Disease|Disorder|false|false||coldnull|Cold Sensation|Finding|false|false||coldnull|Cold Therapy|Procedure|false|false||coldnull|Cold Temperature|Phenomenon|false|false||coldnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Respiratory Status|Finding|false|false||respiratory statusnull|null|Attribute|false|false||respiratory statusnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|COPD exacerbation|Disorder|false|false||COPD exacerbationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Exacerbation|Finding|false|false||exacerbationnull|High dose|LabModifier|false|false||high dosenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Steroids|Drug|false|false||steroids
null|Steroids|Drug|false|false||steroidsnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Tamiflu|Drug|false|false||tamiflu
null|Tamiflu|Drug|false|false||tamiflunull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Oxygen Therapy Care|Procedure|false|false||on oxygennull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Inflammation|Finding|false|false||inflammationnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|prednisone|Drug|false|false||Prednisone
null|prednisone|Drug|false|false||Prednisone
null|prednisone|Drug|false|false||Prednisonenull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|Daily|Time|false|false||day
null|day|Time|false|false||daynull|Daily|Time|false|false||Dailynull|day|Time|false|false||daysnull|Daily|Time|false|false||Dailynull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Daily|Time|false|false||Dailynull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then stop|Finding|false|false||then stopnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycinnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Daily|Time|false|false||Dailynull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|Daily|Time|false|false||day
null|day|Time|false|false||daynull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Tamiflu|Drug|false|false||Tamiflu
null|Tamiflu|Drug|false|false||Tamiflunull|Twice (Numerical Qualifier)|LabModifier|false|false||two timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|day|Time|false|false||daysnull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions