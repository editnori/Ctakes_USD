 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
MEDICINE|158,166
<EOL>|166,167
<EOL>|168,169
Allergies|169,178
:|178,179
<EOL>|180,181
No|181,183
Known|184,189
Allergies|190,199
/|200,201
Adverse|202,209
Drug|210,214
Reactions|215,224
<EOL>|224,225
<EOL>|226,227
Attending|227,236
:|236,237
_|238,239
_|239,240
_|240,241
.|241,242
<EOL>|242,243
<EOL>|244,245
Chief|245,250
Complaint|251,260
:|260,261
<EOL>|261,262
fever|262,267
<EOL>|267,268
<EOL>|269,270
Major|270,275
Surgical|276,284
or|285,287
Invasive|288,296
Procedure|297,306
:|306,307
<EOL>|307,308
none|308,312
<EOL>|312,313
<EOL>|313,314
<EOL>|315,316
History|316,323
of|324,326
Present|327,334
Illness|335,342
:|342,343
<EOL>|343,344
_|344,345
_|345,346
_|346,347
with|348,352
history|353,360
of|361,363
morbid|364,370
obesity|371,378
,|378,379
coronary|380,388
artery|389,395
disease|396,403
,|403,404
<EOL>|405,406
presenting|406,416
today|417,422
with|423,427
cough|428,433
productive|434,444
of|445,447
brown|448,453
sputum|454,460
and|461,464
<EOL>|465,466
fevers|466,472
up|473,475
to|476,478
103.2|479,484
for|485,488
last|489,493
2|494,495
days|496,500
.|500,501
Also|502,506
endorses|507,515
chills|516,522
.|522,523
<EOL>|524,525
Husband|525,532
with|533,537
similar|538,545
symptoms|546,554
2d|555,557
prior|558,563
,|563,564
now|565,568
improving|569,578
without|579,586
<EOL>|587,588
antibiotics|588,599
.|599,600
Denies|601,607
any|608,611
chest|612,617
pain|618,622
but|623,626
states|627,633
that|634,638
he|639,641
she|642,645
has|646,649
<EOL>|650,651
been|651,655
more|656,660
short|661,666
of|667,669
breath|670,676
.|676,677
<EOL>|679,680
<EOL>|681,682
In|682,684
the|685,688
ED|689,691
,|691,692
initial|693,700
VS|701,703
:|703,704
101.3|705,710
97|711,713
168|714,717
/|717,718
58|718,720
18|721,723
93|724,726
%|726,727
ra|728,730
.|730,731
CXR|732,735
showed|736,742
b|743,744
/|744,745
l|745,746
<EOL>|747,748
perihilar|748,757
prominence|758,768
but|769,772
no|773,775
evidence|776,784
of|785,787
CHF|788,791
or|792,794
pneumonia|795,804
.|804,805
CT|806,808
A|809,810
/|810,811
P|811,812
<EOL>|813,814
showed|814,820
no|821,823
acute|824,829
abdominal|830,839
process|840,847
.|847,848
Labs|849,853
notable|854,861
for|862,865
WBC|866,869
7.2|870,873
with|874,878
<EOL>|879,880
81|880,882
%|882,883
N|883,884
,|884,885
TroT|886,890
<|891,892
.01|892,895
x1|896,898
,|898,899
lactate|900,907
2|908,909
,|909,910
UA|911,913
with|914,918
trace|919,924
leuks|925,930
.|930,931
Given|932,937
<EOL>|938,939
clinical|939,947
picture|948,955
and|956,959
fever|960,965
,|965,966
patient|967,974
was|975,978
treated|979,986
for|987,990
presumptive|991,1002
<EOL>|1003,1004
PNA|1004,1007
with|1008,1012
Levofloxacin|1013,1025
750mg|1026,1031
IV|1032,1034
.|1034,1035
She|1036,1039
was|1040,1043
also|1044,1048
given|1049,1054
Ativan|1055,1061
2mg|1062,1065
<EOL>|1066,1067
PO|1067,1069
,|1069,1070
Tylenol|1071,1078
2g|1079,1081
,|1081,1082
Zofran|1083,1089
4mg|1090,1093
.|1093,1094
SpO2|1095,1099
dropped|1100,1107
to|1108,1110
91|1111,1113
&|1113,1114
with|1115,1119
ambulation|1120,1130
.|1130,1131
<EOL>|1132,1133
Pt.|1133,1136
initially|1137,1146
wanted|1147,1153
to|1154,1156
leave|1157,1162
,|1162,1163
but|1164,1167
was|1168,1171
convinced|1172,1181
to|1182,1184
stay|1185,1189
.|1189,1190
VS|1191,1193
at|1194,1196
<EOL>|1197,1198
transfer|1198,1206
:|1206,1207
100.3|1208,1213
98|1214,1216
18|1217,1219
127|1220,1223
/|1223,1224
71|1224,1226
95|1227,1229
%|1229,1230
ra|1230,1232
.|1232,1233
<EOL>|1235,1236
.|1236,1237
<EOL>|1239,1240
Currently|1240,1249
,|1249,1250
she|1251,1254
is|1255,1257
tired|1258,1263
but|1264,1267
denies|1268,1274
F|1275,1276
/|1276,1277
C|1277,1278
/|1278,1279
SOB|1279,1282
.|1282,1283
<EOL>|1285,1286
.|1286,1287
<EOL>|1289,1290
ROS|1290,1293
:|1293,1294
As|1295,1297
per|1298,1301
HPI|1302,1305
<EOL>|1307,1308
<EOL>|1308,1309
<EOL>|1310,1311
Past|1311,1315
Medical|1316,1323
History|1324,1331
:|1331,1332
<EOL>|1332,1333
MYOCARDIAL|1333,1343
INFARCT|1344,1351
-|1352,1353
INFEROPOSTERIOR|1354,1369
<EOL>|1371,1372
HYPERCHOLESTEROLEMIA|1372,1392
<EOL>|1394,1395
DM|1395,1397
(|1398,1399
diabetes|1399,1407
mellitus|1408,1416
)|1416,1417
,|1417,1418
type|1419,1423
2|1424,1425
,|1425,1426
uncontrolled|1427,1439
<EOL>|1441,1442
HYPERTENSION|1442,1454
-|1455,1456
ESSENTIAL|1457,1466
,|1466,1467
UNSPEC|1468,1474
<EOL>|1476,1477
Anemia|1477,1483
<EOL>|1485,1486
Thyroid|1486,1493
nodule|1494,1500
<EOL>|1502,1503
Asymptomatic|1503,1515
carotid|1516,1523
artery|1524,1530
stenosis|1531,1539
<EOL>|1541,1542
OBESITY|1542,1549
-|1550,1551
MORBID|1552,1558
<EOL>|1560,1561
ESOPHAGEAL|1561,1571
REFLUX|1572,1578
<EOL>|1580,1581
HYPOTHYROIDISM|1581,1595
,|1595,1596
UNSPEC|1597,1603
<EOL>|1605,1606
ANXIETY|1606,1613
STATES|1614,1620
,|1620,1621
UNSPEC|1622,1628
<EOL>|1630,1631
DERMATITIS|1631,1641
-|1642,1643
ECZEMATOUS|1644,1654
<EOL>|1656,1657
HEADACHE|1657,1665
<EOL>|1667,1668
COLONIC|1668,1675
ADENOMA|1676,1683
<EOL>|1685,1686
DISC|1686,1690
DISEASE|1691,1698
-|1699,1700
LUMBAR|1701,1707
<EOL>|1709,1710
Ovarian|1710,1717
Retention|1718,1727
Cyst|1728,1732
<EOL>|1734,1735
.|1735,1736
<EOL>|1738,1739
<EOL>|1739,1740
<EOL>|1741,1742
Social|1742,1748
History|1749,1756
:|1756,1757
<EOL>|1757,1758
_|1758,1759
_|1759,1760
_|1760,1761
<EOL>|1761,1762
Family|1762,1768
History|1769,1776
:|1776,1777
<EOL>|1777,1778
Non|1778,1781
contributory|1782,1794
<EOL>|1795,1796
<EOL>|1797,1798
Physical|1798,1806
Exam|1807,1811
:|1811,1812
<EOL>|1812,1813
Physical|1813,1821
Exam|1822,1826
on|1827,1829
Admission|1830,1839
:|1839,1840
<EOL>|1840,1841
VS|1841,1843
-|1844,1845
Temp|1846,1850
98.3|1851,1855
F|1855,1856
,|1856,1857
BP|1858,1860
141|1861,1864
/|1864,1865
61|1865,1867
,|1867,1868
HR|1869,1871
101|1872,1875
,|1875,1876
R|1877,1878
20|1879,1881
,|1881,1882
O2|1883,1885
-|1885,1886
sat|1886,1889
93|1890,1892
%|1892,1893
RA|1894,1896
<EOL>|1898,1899
GENERAL|1899,1906
-|1907,1908
morbidly|1909,1917
obese|1918,1923
female|1924,1930
in|1931,1933
NAD|1934,1937
,|1937,1938
comfortable|1939,1950
,|1950,1951
appropriate|1952,1963
<EOL>|1964,1965
<EOL>|1966,1967
HEENT|1967,1972
-|1973,1974
NC|1975,1977
/|1977,1978
AT|1978,1980
,|1980,1981
PERRLA|1982,1988
,|1988,1989
EOMI|1990,1994
,|1994,1995
sclerae|1996,2003
anicteric|2004,2013
,|2013,2014
MM|2015,2017
slightly|2018,2026
dry|2027,2030
,|2030,2031
<EOL>|2032,2033
OP|2033,2035
clear|2036,2041
<EOL>|2043,2044
NECK|2044,2048
-|2049,2050
supple|2051,2057
,|2057,2058
no|2059,2061
thyromegaly|2062,2073
,|2073,2074
no|2075,2077
JVD|2078,2081
,|2081,2082
no|2083,2085
carotid|2086,2093
bruits|2094,2100
<EOL>|2102,2103
LUNGS|2103,2108
-|2109,2110
very|2111,2115
distant|2116,2123
breath|2124,2130
sounds|2131,2137
,|2137,2138
scattered|2139,2148
exp|2149,2152
wheezes|2153,2160
,|2160,2161
no|2162,2164
<EOL>|2165,2166
crackles|2166,2174
,|2174,2175
resp|2176,2180
unlabored|2181,2190
,|2190,2191
no|2192,2194
accessory|2195,2204
muscle|2205,2211
use|2212,2215
<EOL>|2217,2218
HEART|2218,2223
-|2224,2225
RRR|2226,2229
,|2229,2230
no|2231,2233
MRG|2234,2237
,|2237,2238
nl|2239,2241
S1|2242,2244
-|2244,2245
S2|2245,2247
<EOL>|2249,2250
ABDOMEN|2250,2257
-|2258,2259
NABS|2260,2264
,|2264,2265
obese|2266,2271
,|2271,2272
soft|2273,2277
/|2277,2278
NT|2278,2280
/|2280,2281
ND|2281,2283
,|2283,2284
no|2285,2287
masses|2288,2294
or|2295,2297
HSM|2298,2301
,|2301,2302
no|2303,2305
<EOL>|2306,2307
rebound|2307,2314
/|2314,2315
guarding|2315,2323
<EOL>|2325,2326
EXTREMITIES|2326,2337
-|2338,2339
WWP|2340,2343
,|2343,2344
no|2345,2347
c|2348,2349
/|2349,2350
c|2350,2351
/|2351,2352
e|2352,2353
,|2353,2354
2|2355,2356
+|2356,2357
peripheral|2358,2368
pulses|2369,2375
(|2376,2377
radials|2377,2384
,|2384,2385
DPs|2386,2389
)|2389,2390
<EOL>|2391,2392
<EOL>|2393,2394
SKIN|2394,2398
-|2399,2400
no|2401,2403
rashes|2404,2410
or|2411,2413
lesions|2414,2421
<EOL>|2423,2424
NEURO|2424,2429
-|2430,2431
awake|2432,2437
,|2437,2438
A|2439,2440
&|2440,2441
Ox3|2441,2444
<EOL>|2445,2446
.|2446,2447
<EOL>|2447,2448
Physical|2448,2456
Exam|2457,2461
on|2462,2464
Discharge|2465,2474
:|2474,2475
<EOL>|2475,2476
VS|2476,2478
-|2479,2480
Tm|2481,2483
100.3|2484,2489
Tc|2490,2492
98.6|2493,2497
BP|2498,2500
137|2501,2504
/|2504,2505
46|2505,2507
HR|2508,2510
R|2512,2513
20|2514,2516
O2|2517,2519
-|2519,2520
sat|2520,2523
94|2524,2526
%|2526,2527
RA|2528,2530
<EOL>|2532,2533
GENERAL|2533,2540
-|2541,2542
morbidly|2543,2551
obese|2552,2557
female|2558,2564
in|2565,2567
NAD|2568,2571
,|2571,2572
comfortable|2573,2584
,|2584,2585
appropriate|2586,2597
<EOL>|2598,2599
<EOL>|2600,2601
HEENT|2601,2606
-|2607,2608
NC|2609,2611
/|2611,2612
AT|2612,2614
,|2614,2615
PERRLA|2616,2622
,|2622,2623
EOMI|2624,2628
,|2628,2629
sclerae|2630,2637
anicteric|2638,2647
,|2647,2648
MM|2649,2651
slightly|2652,2660
dry|2661,2664
,|2664,2665
<EOL>|2666,2667
OP|2667,2669
clear|2670,2675
<EOL>|2677,2678
NECK|2678,2682
-|2683,2684
supple|2685,2691
,|2691,2692
no|2693,2695
thyromegaly|2696,2707
,|2707,2708
no|2709,2711
JVD|2712,2715
,|2715,2716
no|2717,2719
carotid|2720,2727
bruits|2728,2734
<EOL>|2736,2737
LUNGS|2737,2742
-|2743,2744
very|2745,2749
distant|2750,2757
breath|2758,2764
sounds|2765,2771
,|2771,2772
few|2773,2776
scattered|2777,2786
exp|2787,2790
wheezes|2791,2798
,|2798,2799
<EOL>|2800,2801
no|2801,2803
crackles|2804,2812
,|2812,2813
resp|2814,2818
unlabored|2819,2828
,|2828,2829
no|2830,2832
accessory|2833,2842
muscle|2843,2849
use|2850,2853
<EOL>|2855,2856
HEART|2856,2861
-|2862,2863
RRR|2864,2867
,|2867,2868
no|2869,2871
MRG|2872,2875
,|2875,2876
nl|2877,2879
S1|2880,2882
-|2882,2883
S2|2883,2885
<EOL>|2887,2888
ABDOMEN|2888,2895
-|2896,2897
NABS|2898,2902
,|2902,2903
obese|2904,2909
,|2909,2910
soft|2911,2915
/|2915,2916
NT|2916,2918
/|2918,2919
ND|2919,2921
,|2921,2922
no|2923,2925
masses|2926,2932
or|2933,2935
HSM|2936,2939
,|2939,2940
no|2941,2943
<EOL>|2944,2945
rebound|2945,2952
/|2952,2953
guarding|2953,2961
<EOL>|2963,2964
EXTREMITIES|2964,2975
-|2976,2977
WWP|2978,2981
,|2981,2982
no|2983,2985
c|2986,2987
/|2987,2988
c|2988,2989
/|2989,2990
e|2990,2991
,|2991,2992
2|2993,2994
+|2994,2995
peripheral|2996,3006
pulses|3007,3013
(|3014,3015
radials|3015,3022
,|3022,3023
DPs|3024,3027
)|3027,3028
<EOL>|3029,3030
<EOL>|3031,3032
SKIN|3032,3036
-|3037,3038
no|3039,3041
rashes|3042,3048
or|3049,3051
lesions|3052,3059
<EOL>|3061,3062
NEURO|3062,3067
-|3068,3069
awake|3070,3075
,|3075,3076
A|3077,3078
&|3078,3079
Ox3|3079,3082
<EOL>|3084,3085
<EOL>|3085,3086
<EOL>|3087,3088
Pertinent|3088,3097
Results|3098,3105
:|3105,3106
<EOL>|3106,3107
Labs|3107,3111
on|3112,3114
Admission|3115,3124
:|3124,3125
<EOL>|3125,3126
<EOL>|3126,3127
_|3127,3128
_|3128,3129
_|3129,3130
10|3131,3133
:|3133,3134
00PM|3134,3138
WBC|3141,3144
-|3144,3145
7.2|3145,3148
RBC|3149,3152
-|3152,3153
4|3153,3154
.|3154,3155
11|3155,3157
*|3157,3158
HGB|3159,3162
-|3162,3163
11|3163,3165
.|3165,3166
5|3166,3167
*|3167,3168
HCT|3169,3172
-|3172,3173
35|3173,3175
.|3175,3176
4|3176,3177
*|3177,3178
MCV|3179,3182
-|3182,3183
86|3183,3185
<EOL>|3186,3187
MCH|3187,3190
-|3190,3191
27.8|3191,3195
MCHC|3196,3200
-|3200,3201
32.3|3201,3205
RDW|3206,3209
-|3209,3210
15.5|3210,3214
<EOL>|3214,3215
_|3215,3216
_|3216,3217
_|3217,3218
10|3219,3221
:|3221,3222
00PM|3222,3226
NEUTS|3229,3234
-|3234,3235
81|3235,3237
.|3237,3238
1|3238,3239
*|3239,3240
LYMPHS|3241,3247
-|3247,3248
10|3248,3250
.|3250,3251
8|3251,3252
*|3252,3253
MONOS|3254,3259
-|3259,3260
6.9|3260,3263
EOS|3264,3267
-|3267,3268
0.8|3268,3271
<EOL>|3272,3273
BASOS|3273,3278
-|3278,3279
0.4|3279,3282
<EOL>|3282,3283
_|3283,3284
_|3284,3285
_|3285,3286
10|3287,3289
:|3289,3290
00PM|3290,3294
cTropnT|3297,3304
-|3304,3305
<|3305,3306
0|3306,3307
.|3307,3308
01|3308,3310
<EOL>|3310,3311
_|3311,3312
_|3312,3313
_|3313,3314
10|3315,3317
:|3317,3318
00PM|3318,3322
LIPASE|3325,3331
-|3331,3332
21|3332,3334
<EOL>|3334,3335
_|3335,3336
_|3336,3337
_|3337,3338
10|3339,3341
:|3341,3342
00PM|3342,3346
ALT|3349,3352
(|3352,3353
SGPT|3353,3357
)|3357,3358
-|3358,3359
54|3359,3361
*|3361,3362
AST|3363,3366
(|3366,3367
SGOT|3367,3371
)|3371,3372
-|3372,3373
50|3373,3375
*|3375,3376
ALK|3377,3380
PHOS|3381,3385
-|3385,3386
64|3386,3388
TOT|3389,3392
<EOL>|3393,3394
BILI|3394,3398
-|3398,3399
0.4|3399,3402
<EOL>|3402,3403
_|3403,3404
_|3404,3405
_|3405,3406
10|3407,3409
:|3409,3410
00PM|3410,3414
GLUCOSE|3417,3424
-|3424,3425
119|3425,3428
*|3428,3429
UREA|3430,3434
N|3435,3436
-|3436,3437
14|3437,3439
CREAT|3440,3445
-|3445,3446
0.7|3446,3449
SODIUM|3450,3456
-|3456,3457
136|3457,3460
<EOL>|3461,3462
POTASSIUM|3462,3471
-|3471,3472
3.9|3472,3475
CHLORIDE|3476,3484
-|3484,3485
98|3485,3487
TOTAL|3488,3493
CO2|3494,3497
-|3497,3498
28|3498,3500
ANION|3501,3506
GAP|3507,3510
-|3510,3511
14|3511,3513
<EOL>|3513,3514
_|3514,3515
_|3515,3516
_|3516,3517
10|3518,3520
:|3520,3521
11PM|3521,3525
LACTATE|3528,3535
-|3535,3536
2.0|3536,3539
<EOL>|3539,3540
_|3540,3541
_|3541,3542
_|3542,3543
10|3544,3546
:|3546,3547
47PM|3547,3551
URINE|3552,3557
COLOR|3559,3564
-|3564,3565
Yellow|3565,3571
APPEAR|3572,3578
-|3578,3579
Clear|3579,3584
SP|3585,3587
_|3588,3589
_|3589,3590
_|3590,3591
<EOL>|3591,3592
_|3592,3593
_|3593,3594
_|3594,3595
10|3596,3598
:|3598,3599
47PM|3599,3603
URINE|3604,3609
BLOOD|3611,3616
-|3616,3617
NEG|3617,3620
NITRITE|3621,3628
-|3628,3629
NEG|3629,3632
PROTEIN|3633,3640
-|3640,3641
NEG|3641,3644
<EOL>|3645,3646
GLUCOSE|3646,3653
-|3653,3654
NEG|3654,3657
KETONE|3658,3664
-|3664,3665
NEG|3665,3668
BILIRUBIN|3669,3678
-|3678,3679
NEG|3679,3682
UROBILNGN|3683,3692
-|3692,3693
NEG|3693,3696
PH|3697,3699
-|3699,3700
5.5|3700,3703
<EOL>|3704,3705
LEUK|3705,3709
-|3709,3710
TR|3710,3712
<EOL>|3712,3713
_|3713,3714
_|3714,3715
_|3715,3716
10|3717,3719
:|3719,3720
47PM|3720,3724
URINE|3725,3730
RBC|3732,3735
-|3735,3736
<|3736,3737
1|3737,3738
WBC|3739,3742
-|3742,3743
4|3743,3744
BACTERIA|3745,3753
-|3753,3754
NONE|3754,3758
YEAST|3759,3764
-|3764,3765
NONE|3765,3769
<EOL>|3770,3771
EPI|3771,3774
-|3774,3775
1|3775,3776
<EOL>|3776,3777
_|3777,3778
_|3778,3779
_|3779,3780
10|3781,3783
:|3783,3784
47PM|3784,3788
URINE|3789,3794
MUCOUS|3796,3802
-|3802,3803
RARE|3803,3807
<EOL>|3807,3808
<EOL>|3808,3809
Imaging|3809,3816
:|3816,3817
<EOL>|3817,3818
<EOL>|3818,3819
CXR|3819,3822
_|3823,3824
_|3824,3825
_|3825,3826
:|3826,3827
<EOL>|3827,3828
IMPRESSION|3828,3838
:|3838,3839
Mild|3841,3845
perihilar|3846,3855
prominence|3856,3866
,|3866,3867
suspected|3868,3877
to|3878,3880
represent|3881,3890
<EOL>|3891,3892
mildly|3892,3898
prominent|3899,3908
pulmonary|3909,3918
vessels|3919,3926
without|3927,3934
definite|3935,3943
pneumonia|3944,3953
.|3953,3954
<EOL>|3956,3957
Streaky|3957,3964
left|3965,3969
basilar|3970,3977
opacification|3978,3991
seen|3992,3996
only|3997,4001
on|4002,4004
the|4005,4008
frontal|4009,4016
view|4017,4021
<EOL>|4022,4023
is|4023,4025
probably|4026,4034
due|4035,4038
to|4039,4041
minor|4042,4047
atelectasis|4048,4059
or|4060,4062
scarring|4063,4071
.|4071,4072
<EOL>|4073,4074
.|4074,4075
<EOL>|4077,4078
CT|4078,4080
A|4081,4082
/|4082,4083
P|4083,4084
_|4085,4086
_|4086,4087
_|4087,4088
:|4088,4089
<EOL>|4090,4091
1|4091,4092
.|4092,4093
No|4095,4097
acute|4098,4103
intra-abdominal|4104,4119
pathology|4120,4129
.|4129,4130
There|4131,4136
is|4137,4139
diverticulosis|4140,4154
<EOL>|4155,4156
and|4156,4159
sequelae|4160,4168
of|4169,4171
prior|4172,4177
inflammation|4178,4190
,|4190,4191
but|4192,4195
no|4196,4198
active|4199,4205
<EOL>|4206,4207
diverticulitis|4207,4221
.|4221,4222
<EOL>|4223,4224
2.|4224,4226
3|4228,4229
-|4229,4230
mm|4230,4232
nodule|4233,4239
seen|4240,4244
along|4245,4250
the|4251,4254
right|4255,4260
major|4261,4266
fissure|4267,4274
and|4275,4278
right|4279,4284
<EOL>|4285,4286
lower|4286,4291
lobe|4292,4296
.|4296,4297
According|4299,4308
to|4309,4311
_|4312,4313
_|4313,4314
_|4314,4315
guidelines|4316,4326
,|4326,4327
in|4328,4330
the|4331,4334
absence|4335,4342
<EOL>|4343,4344
of|4344,4346
risk|4347,4351
factors|4352,4359
,|4359,4360
no|4361,4363
further|4364,4371
followup|4372,4380
is|4381,4383
needed|4384,4390
.|4390,4391
If|4393,4395
patient|4396,4403
has|4404,4407
<EOL>|4408,4409
risk|4409,4413
factors|4414,4421
such|4422,4426
as|4427,4429
smoking|4430,4437
,|4437,4438
followup|4439,4447
chest|4448,4453
CT|4454,4456
at|4457,4459
12|4460,4462
months|4463,4469
is|4470,4472
<EOL>|4473,4474
recommended|4474,4485
to|4486,4488
document|4489,4497
stability|4498,4507
.|4507,4508
<EOL>|4509,4510
<EOL>|4510,4511
CXR|4511,4514
_|4515,4516
_|4516,4517
_|4517,4518
:|4518,4519
<EOL>|4519,4520
There|4520,4525
are|4526,4529
low|4530,4533
lung|4534,4538
volumes|4539,4546
with|4547,4551
an|4552,4554
appearance|4555,4565
of|4566,4568
bronchovascular|4569,4584
<EOL>|4585,4586
crowding|4586,4594
.|4594,4595
Despite|4597,4604
this|4605,4609
,|4609,4610
there|4611,4616
is|4617,4619
likely|4620,4626
mild|4627,4631
vascular|4632,4640
<EOL>|4641,4642
congestion|4642,4652
and|4653,4656
edema|4657,4662
.|4662,4663
No|4665,4667
focal|4668,4673
consolidation|4674,4687
is|4688,4690
seen|4691,4695
with|4696,4700
<EOL>|4701,4702
linear|4702,4708
bibasilar|4709,4718
atelectasis|4719,4730
.|4730,4731
The|4733,4736
heart|4737,4742
is|4743,4745
top|4746,4749
normal|4750,4756
in|4757,4759
size|4760,4764
<EOL>|4765,4766
with|4766,4770
aortic|4771,4777
totuosity|4778,4787
.|4787,4788
<EOL>|4790,4791
<EOL>|4793,4794
IMPRESSION|4794,4804
:|4804,4805
Mild|4807,4811
pulmonary|4812,4821
edema|4822,4827
<EOL>|4829,4830
.|4830,4831
<EOL>|4831,4832
Urine|4832,4837
legionella|4838,4848
-|4848,4849
negative|4849,4857
<EOL>|4857,4858
.|4858,4859
<EOL>|4859,4860
Labs|4860,4864
on|4865,4867
Discharge|4868,4877
:|4877,4878
<EOL>|4878,4879
.|4879,4880
<EOL>|4880,4881
_|4881,4882
_|4882,4883
_|4883,4884
05|4885,4887
:|4887,4888
25AM|4888,4892
BLOOD|4893,4898
WBC|4899,4902
-|4902,4903
11|4903,4905
.|4905,4906
6|4906,4907
*|4907,4908
RBC|4909,4912
-|4912,4913
3|4913,4914
.|4914,4915
34|4915,4917
*|4917,4918
Hgb|4919,4922
-|4922,4923
9|4923,4924
.|4924,4925
3|4925,4926
*|4926,4927
Hct|4928,4931
-|4931,4932
28|4932,4934
.|4934,4935
5|4935,4936
*|4936,4937
<EOL>|4938,4939
MCV|4939,4942
-|4942,4943
86|4943,4945
MCH|4946,4949
-|4949,4950
27.9|4950,4954
MCHC|4955,4959
-|4959,4960
32.6|4960,4964
RDW|4965,4968
-|4968,4969
15|4969,4971
.|4971,4972
9|4972,4973
*|4973,4974
Plt|4975,4978
_|4979,4980
_|4980,4981
_|4981,4982
<EOL>|4982,4983
_|4983,4984
_|4984,4985
_|4985,4986
05|4987,4989
:|4989,4990
25AM|4990,4994
BLOOD|4995,5000
_|5001,5002
_|5002,5003
_|5003,5004
PTT|5005,5008
-|5008,5009
33.8|5009,5013
_|5014,5015
_|5015,5016
_|5016,5017
<EOL>|5017,5018
_|5018,5019
_|5019,5020
_|5020,5021
05|5022,5024
:|5024,5025
25AM|5025,5029
BLOOD|5030,5035
Glucose|5036,5043
-|5043,5044
106|5044,5047
*|5047,5048
UreaN|5049,5054
-|5054,5055
15|5055,5057
Creat|5058,5063
-|5063,5064
0.6|5064,5067
Na|5068,5070
-|5070,5071
134|5071,5074
<EOL>|5075,5076
K|5076,5077
-|5077,5078
3.8|5078,5081
Cl|5082,5084
-|5084,5085
96|5085,5087
HCO3|5088,5092
-|5092,5093
28|5093,5095
AnGap|5096,5101
-|5101,5102
14|5102,5104
<EOL>|5104,5105
_|5105,5106
_|5106,5107
_|5107,5108
06|5109,5111
:|5111,5112
15AM|5112,5116
BLOOD|5117,5122
ALT|5123,5126
-|5126,5127
68|5127,5129
*|5129,5130
AST|5131,5134
-|5134,5135
50|5135,5137
*|5137,5138
AlkPhos|5139,5146
-|5146,5147
66|5147,5149
TotBili|5150,5157
-|5157,5158
0.5|5158,5161
<EOL>|5161,5162
_|5162,5163
_|5163,5164
_|5164,5165
05|5166,5168
:|5168,5169
25AM|5169,5173
BLOOD|5174,5179
Calcium|5180,5187
-|5187,5188
8.7|5188,5191
Phos|5192,5196
-|5196,5197
2|5197,5198
.|5198,5199
4|5199,5200
*|5200,5201
Mg|5202,5204
-|5204,5205
1.8|5205,5208
<EOL>|5208,5209
_|5209,5210
_|5210,5211
_|5211,5212
10|5213,5215
:|5215,5216
47PM|5216,5220
URINE|5221,5226
Color|5227,5232
-|5232,5233
Yellow|5233,5239
Appear|5240,5246
-|5246,5247
Clear|5247,5252
Sp|5253,5255
_|5256,5257
_|5257,5258
_|5258,5259
<EOL>|5259,5260
_|5260,5261
_|5261,5262
_|5262,5263
10|5264,5266
:|5266,5267
47PM|5267,5271
URINE|5272,5277
Blood|5278,5283
-|5283,5284
NEG|5284,5287
Nitrite|5288,5295
-|5295,5296
NEG|5296,5299
Protein|5300,5307
-|5307,5308
NEG|5308,5311
<EOL>|5312,5313
Glucose|5313,5320
-|5320,5321
NEG|5321,5324
Ketone|5325,5331
-|5331,5332
NEG|5332,5335
Bilirub|5336,5343
-|5343,5344
NEG|5344,5347
Urobiln|5348,5355
-|5355,5356
NEG|5356,5359
pH|5360,5362
-|5362,5363
5.5|5363,5366
Leuks|5367,5372
-|5372,5373
TR|5373,5375
<EOL>|5375,5376
_|5376,5377
_|5377,5378
_|5378,5379
10|5380,5382
:|5382,5383
47PM|5383,5387
URINE|5388,5393
RBC|5394,5397
-|5397,5398
<|5398,5399
1|5399,5400
WBC|5401,5404
-|5404,5405
4|5405,5406
Bacteri|5407,5414
-|5414,5415
NONE|5415,5419
Yeast|5420,5425
-|5425,5426
NONE|5426,5430
<EOL>|5431,5432
Epi|5432,5435
-|5435,5436
_|5436,5437
_|5437,5438
_|5438,5439
with|5440,5444
diabetes|5445,5453
,|5453,5454
morbid|5455,5461
obesity|5462,5469
,|5469,5470
s|5471,5472
/|5472,5473
p|5473,5474
MI|5475,5477
,|5477,5478
HTN|5479,5482
who|5483,5486
presents|5487,5495
with|5496,5500
<EOL>|5501,5502
2|5502,5503
days|5504,5508
of|5509,5511
fevers|5512,5518
and|5519,5522
cough|5523,5528
productive|5529,5539
of|5540,5542
rust|5543,5547
colored|5548,5555
sputum|5556,5562
<EOL>|5563,5564
with|5564,5568
associated|5569,5579
SOB|5580,5583
.|5583,5584
<EOL>|5586,5587
.|5587,5588
<EOL>|5590,5591
#|5591,5592
Fevers|5593,5599
:|5599,5600
Likely|5601,5607
secondary|5608,5617
to|5618,5620
pneumonia|5621,5630
,|5630,5631
but|5632,5635
possibly|5636,5644
a|5645,5646
viral|5647,5652
<EOL>|5653,5654
illness|5654,5661
.|5661,5662
Most|5663,5667
likely|5668,5674
not|5675,5678
bacterial|5679,5688
process|5689,5696
but|5697,5700
no|5701,5703
leukocytosis|5704,5716
,|5716,5717
<EOL>|5718,5719
just|5719,5723
PMN|5724,5727
predominance|5728,5740
.|5740,5741
Urine|5742,5747
legionella|5748,5758
neg|5759,5762
.|5762,5763
CXR|5764,5767
underwhelming|5768,5781
<EOL>|5782,5783
for|5783,5786
pnuemonia|5787,5796
but|5797,5800
given|5801,5806
poor|5807,5811
PO|5812,5814
intake|5815,5821
and|5822,5825
overall|5826,5833
constellation|5834,5847
<EOL>|5848,5849
of|5849,5851
symptoms|5852,5860
without|5861,5868
other|5869,5874
localizing|5875,5885
source|5886,5892
and|5893,5896
neg|5897,5900
CT|5901,5903
,|5903,5904
so|5905,5907
<EOL>|5908,5909
patient|5909,5916
was|5917,5920
treated|5921,5928
presumptively|5929,5942
for|5943,5946
CAP|5947,5950
.|5950,5951
O2|5953,5955
sats|5956,5960
stable|5961,5967
on|5968,5970
<EOL>|5971,5972
room|5972,5976
air|5977,5980
during|5981,5987
the|5988,5991
day|5992,5995
,|5995,5996
but|5997,6000
at|6001,6003
night|6004,6009
de-satted|6010,6019
.|6019,6020
On|6022,6024
exam|6025,6029
,|6029,6030
lungs|6031,6036
<EOL>|6037,6038
with|6038,6042
improved|6043,6051
wheezing|6052,6060
since|6061,6066
yesterday|6067,6076
.|6076,6077
With|6078,6082
ambulation|6083,6093
,|6093,6094
O2|6095,6097
87|6098,6100
,|6100,6101
<EOL>|6102,6103
on|6103,6105
_|6106,6107
_|6107,6108
_|6108,6109
,|6109,6110
repeat|6111,6117
cxr|6118,6121
with|6122,6126
pulm|6127,6131
edema|6132,6137
likely|6138,6144
due|6145,6148
to|6149,6151
IV|6152,6154
fluid|6155,6160
bolus|6161,6166
<EOL>|6167,6168
day|6168,6171
prior|6172,6177
.|6177,6178
She|6179,6182
was|6183,6186
given|6187,6192
lasix|6193,6198
40mg|6199,6203
POx1|6204,6208
.|6208,6209
On|6211,6213
day|6214,6217
of|6218,6220
d|6221,6222
/|6222,6223
c|6223,6224
,|6224,6225
sats|6226,6230
<EOL>|6231,6232
mid|6232,6235
_|6236,6237
_|6237,6238
_|6238,6239
on|6240,6242
RA|6243,6245
,|6245,6246
down|6247,6251
to|6252,6254
88|6255,6257
%|6257,6258
with|6259,6263
prolonged|6264,6273
ambulation|6274,6284
.|6284,6285
Pt|6287,6289
not|6290,6293
<EOL>|6294,6295
subjectively|6295,6307
SOB|6308,6311
,|6311,6312
likely|6313,6319
this|6320,6324
is|6325,6327
baseline|6328,6336
given|6337,6342
pt|6343,6345
's|6345,6347
habitus|6348,6355
.|6355,6356
<EOL>|6358,6359
Treated|6359,6366
with|6367,6371
albuterol|6372,6381
nebs|6382,6386
and|6387,6390
Levofloxacin|6391,6403
750mg|6404,6409
PO|6410,6412
daily|6413,6418
.|6418,6419
On|6421,6423
<EOL>|6424,6425
d|6425,6426
/|6426,6427
c|6427,6428
,|6428,6429
will|6430,6434
complete|6435,6443
5|6444,6445
day|6446,6449
course|6450,6456
of|6457,6459
levofloxacin|6460,6472
.|6472,6473
<EOL>|6475,6476
.|6476,6477
<EOL>|6479,6480
#|6480,6481
Hypotnatremia|6482,6495
:|6495,6496
Na|6497,6499
134|6500,6503
on|6504,6506
am|6507,6509
of|6510,6512
discharge|6513,6522
,|6522,6523
improved|6524,6532
from|6533,6537
lowest|6538,6544
<EOL>|6545,6546
of|6546,6548
129|6549,6552
.|6553,6554
Based|6556,6561
on|6562,6564
urine|6565,6570
lytes|6571,6576
/|6576,6577
osm|6577,6580
and|6581,6584
serum|6585,6590
osm|6591,6594
,|6594,6595
most|6596,6600
likely|6601,6607
<EOL>|6608,6609
SIADH|6609,6614
secondary|6615,6624
to|6625,6627
pulmonary|6628,6637
process|6638,6645
.|6645,6646
<EOL>|6646,6647
.|6647,6648
<EOL>|6648,6649
#|6649,6650
Diabetes|6651,6659
:|6659,6660
Stable|6661,6667
.|6667,6668
Continued|6670,6679
home|6680,6684
Lantus|6685,6691
100U|6692,6696
qhs|6697,6700
and|6701,6704
ISS|6705,6708
.|6708,6709
<EOL>|6711,6712
Held|6712,6716
metformin|6717,6726
in|6727,6729
house|6730,6735
.|6735,6736
Was|6738,6741
on|6742,6744
diabetic|6745,6753
diet|6754,6758
.|6758,6759
<EOL>|6761,6762
.|6762,6763
<EOL>|6765,6766
#|6766,6767
HTN|6768,6771
:|6771,6772
Continued|6773,6782
home|6783,6787
lisinopril|6788,6798
,|6798,6799
metoprolol|6800,6810
.|6810,6811
Held|6813,6817
lasix|6818,6823
<EOL>|6824,6825
initially|6825,6834
in|6835,6837
setting|6838,6845
of|6846,6848
dehydration|6849,6860
initially|6861,6870
.|6870,6871
Re-started|6873,6883
on|6884,6886
<EOL>|6887,6888
d|6888,6889
/|6889,6890
c|6890,6891
.|6891,6892
<EOL>|6894,6895
.|6895,6896
<EOL>|6898,6899
#|6899,6900
CAD|6901,6904
:|6904,6905
No|6906,6908
CP|6909,6911
now|6912,6915
,|6915,6916
ECG|6917,6920
shows|6921,6926
<|6927,6928
1mm|6928,6931
STD|6932,6935
laterally|6936,6945
,|6945,6946
c|6947,6948
/|6948,6949
w|6949,6950
prior|6951,6956
.|6956,6957
<EOL>|6958,6959
Continued|6959,6968
home|6969,6973
asa|6974,6977
,|6977,6978
metoprolol|6979,6989
.|6989,6990
Heart|6991,6996
healthy|6997,7004
diet|7005,7009
.|7009,7010
<EOL>|7011,7012
.|7012,7013
<EOL>|7015,7016
#|7016,7017
HL|7018,7020
:|7020,7021
Stable|7022,7028
.|7028,7029
Continued|7031,7040
home|7041,7045
simvastatin|7046,7057
pending|7058,7065
med|7066,7069
rec|7070,7073
given|7074,7079
<EOL>|7080,7081
80mg|7081,7085
.|7085,7086
<EOL>|7088,7089
.|7089,7090
<EOL>|7092,7093
#|7093,7094
Anxiety|7095,7102
:|7102,7103
Stable|7104,7110
.|7110,7111
Continued|7113,7122
home|7123,7127
lorazepam|7128,7137
,|7137,7138
escitalopram|7139,7151
.|7151,7152
<EOL>|7154,7155
.|7155,7156
<EOL>|7158,7159
#|7159,7160
Anemia|7161,7167
:|7167,7168
Hct|7169,7172
now|7173,7176
at|7177,7179
baseline|7180,7188
35|7189,7191
.|7191,7192
<EOL>|7195,7196
.|7196,7197
<EOL>|7199,7200
#|7200,7201
GERD|7202,7206
:|7206,7207
Stable|7208,7214
.|7214,7215
Substituted|7217,7228
omeprazole|7229,7239
for|7240,7243
home|7244,7248
esomeprazole|7249,7261
.|7261,7262
<EOL>|7262,7263
.|7263,7264
<EOL>|7264,7265
#|7265,7266
incidental|7266,7276
radiographic|7277,7289
findings|7290,7298
-|7298,7299
pulmonary|7299,7308
nodule|7309,7315
.|7315,7316
Will|7317,7321
require|7322,7329
<EOL>|7330,7331
follow|7331,7337
up|7338,7340
.|7340,7341
<EOL>|7343,7344
.|7344,7345
<EOL>|7347,7348
TRANSITIONS|7348,7359
OF|7360,7362
CARE|7363,7367
:|7367,7368
<EOL>|7368,7369
-|7369,7370
will|7371,7375
complete|7376,7384
day|7385,7388
5|7389,7390
of|7391,7393
levofloxacin|7394,7406
course|7407,7413
on|7414,7416
_|7417,7418
_|7418,7419
_|7419,7420
<EOL>|7420,7421
-|7421,7422
will|7423,7427
have|7428,7432
labs|7433,7437
checked|7438,7445
(|7446,7447
particularly|7447,7459
Na|7460,7462
)|7462,7463
and|7464,7467
faxed|7468,7473
to|7474,7476
PCP|7477,7480
_|7481,7482
_|7482,7483
_|7483,7484
<EOL>|7485,7486
_|7486,7487
_|7487,7488
_|7488,7489
<EOL>|7489,7490
-|7490,7491
will|7492,7496
f|7497,7498
/|7498,7499
u|7499,7500
with|7501,7505
PCP|7506,7509
next|7510,7514
week|7515,7519
<EOL>|7519,7520
-|7520,7521
3mm|7522,7525
lung|7526,7530
nodule|7531,7537
seen|7538,7542
on|7543,7545
CXR|7546,7549
;|7549,7550
can|7551,7554
be|7555,7557
followed|7558,7566
as|7567,7569
outpt|7570,7575
<EOL>|7575,7576
-|7576,7577
CODE|7578,7582
:|7582,7583
Confirmed|7584,7593
full|7594,7598
<EOL>|7600,7601
-|7601,7602
CONTACT|7603,7610
:|7610,7611
Husband|7612,7619
_|7620,7621
_|7621,7622
_|7622,7623
_|7624,7625
_|7625,7626
_|7626,7627
<EOL>|7629,7630
<EOL>|7630,7631
<EOL>|7632,7633
_|7633,7634
_|7634,7635
_|7635,7636
on|7637,7639
Admission|7640,7649
:|7649,7650
<EOL>|7650,7651
Humalog|7651,7658
SSI|7659,7662
<EOL>|7664,7665
Lasix|7665,7670
40mg|7671,7675
daily|7676,7681
<EOL>|7683,7684
Dicyclomine|7684,7695
10mg|7696,7700
Q4|7701,7703
-|7703,7704
6H|7704,7706
:|7706,7707
PRN|7707,7710
<EOL>|7712,7713
Levothyroxine|7713,7726
25mcg|7727,7732
daily|7733,7738
<EOL>|7740,7741
Escitalopram|7741,7753
20mg|7754,7758
daily|7759,7764
<EOL>|7766,7767
Metoprolol|7767,7777
succinate|7778,7787
50mg|7788,7792
daily|7793,7798
<EOL>|7800,7801
Lantus|7801,7807
92|7808,7810
units|7811,7816
QHS|7817,7820
<EOL>|7822,7823
Vicodin|7823,7830
1|7831,7832
tab|7833,7836
Q4|7837,7839
-|7839,7840
6H|7840,7842
:|7842,7843
PRN|7843,7846
<EOL>|7848,7849
Lorazepam|7849,7858
2mg|7859,7862
QHS|7863,7866
:|7866,7867
PRN|7867,7870
<EOL>|7872,7873
Esomeprazole|7873,7885
40mg|7886,7890
BID|7891,7894
<EOL>|7896,7897
Lisinopril|7897,7907
20mg|7908,7912
daily|7913,7918
<EOL>|7920,7921
Simvastatin|7921,7932
80mg|7933,7937
QHS|7938,7941
<EOL>|7943,7944
Metformin|7944,7953
1000mg|7954,7960
BID|7961,7964
<EOL>|7966,7967
Ferrous|7967,7974
sulfate|7975,7982
325mg|7983,7988
TID|7989,7992
<EOL>|7994,7995
<EOL>|7995,7996
<EOL>|7997,7998
Discharge|7998,8007
Medications|8008,8019
:|8019,8020
<EOL>|8020,8021
1.|8021,8023
Escitalopram|8024,8036
Oxalate|8037,8044
20|8045,8047
mg|8048,8050
PO|8051,8053
DAILY|8054,8059
<EOL>|8060,8061
2.|8061,8063
Lisinopril|8064,8074
20|8075,8077
mg|8078,8080
PO|8081,8083
DAILY|8084,8089
<EOL>|8090,8091
hold|8091,8095
for|8096,8099
sbp|8100,8103
<|8103,8104
100|8104,8107
<EOL>|8108,8109
3.|8109,8111
esomeprazole|8112,8124
magnesium|8125,8134
*|8135,8136
NF|8136,8138
*|8138,8139
40|8140,8142
mg|8143,8145
Oral|8146,8150
BID|8151,8154
<EOL>|8155,8156
4.|8156,8158
Ferrous|8159,8166
Sulfate|8167,8174
325|8175,8178
mg|8179,8181
PO|8182,8184
TID|8185,8188
<EOL>|8189,8190
5.|8190,8192
DiCYCLOmine|8193,8204
10|8205,8207
mg|8208,8210
PO|8211,8213
QID|8214,8217
:|8217,8218
PRN|8218,8221
pain|8222,8226
<EOL>|8227,8228
6.|8228,8230
Levothyroxine|8231,8244
Sodium|8245,8251
25|8252,8254
mcg|8255,8258
PO|8259,8261
DAILY|8262,8267
<EOL>|8268,8269
7.|8269,8271
Metoprolol|8272,8282
Succinate|8283,8292
XL|8293,8295
50|8296,8298
mg|8299,8301
PO|8302,8304
DAILY|8305,8310
<EOL>|8311,8312
8.|8312,8314
Lorazepam|8315,8324
2|8325,8326
mg|8327,8329
PO|8330,8332
HS|8333,8335
:|8335,8336
PRN|8336,8339
insomnia|8340,8348
<EOL>|8349,8350
9.|8350,8352
Glargine|8353,8361
100|8362,8365
Units|8366,8371
Bedtime|8372,8379
<EOL>|8379,8380
Insulin|8380,8387
SC|8388,8390
Sliding|8391,8398
Scale|8399,8404
using|8405,8410
HUM|8411,8414
InsulinMax|8415,8425
Dose|8426,8430
Override|8431,8439
<EOL>|8440,8441
Reason|8441,8447
:|8447,8448
home|8449,8453
dosing|8454,8460
<EOL>|8460,8461
<EOL>|8461,8462
10.|8462,8465
Levofloxacin|8466,8478
750|8479,8482
mg|8483,8485
PO|8486,8488
DAILY|8489,8494
Start|8495,8500
:|8500,8501
In|8502,8504
am|8505,8507
<EOL>|8508,8509
last|8509,8513
day|8514,8517
is|8518,8520
_|8521,8522
_|8522,8523
_|8523,8524
<EOL>|8525,8526
RX|8526,8528
*|8529,8530
levofloxacin|8530,8542
750|8543,8546
mg|8547,8549
once|8550,8554
a|8555,8556
day|8557,8560
Disp|8561,8565
#|8566,8567
*|8567,8568
1|8568,8569
Tablet|8570,8576
Refills|8577,8584
:|8584,8585
*|8585,8586
0|8586,8587
<EOL>|8587,8588
11.|8588,8591
Hydrocodone|8592,8603
-|8603,8604
Acetaminophen|8604,8617
(|8618,8619
5mg|8619,8622
-|8622,8623
500mg|8623,8628
1|8629,8630
TAB|8631,8634
PO|8635,8637
Q6H|8638,8641
:|8641,8642
PRN|8642,8645
pain|8646,8650
<EOL>|8651,8652
hold|8652,8656
for|8657,8660
sedation|8661,8669
,|8669,8670
RR|8671,8673
<|8673,8674
10|8674,8676
<EOL>|8677,8678
12.|8678,8681
Simvastatin|8682,8693
80|8694,8696
mg|8697,8699
PO|8700,8702
DAILY|8703,8708
<EOL>|8709,8710
13.|8710,8713
MetFORMIN|8714,8723
(|8724,8725
Glucophage|8725,8735
)|8735,8736
1000|8737,8741
mg|8742,8744
PO|8745,8747
BID|8748,8751
<EOL>|8752,8753
14.|8753,8756
Furosemide|8757,8767
40|8768,8770
mg|8771,8773
PO|8774,8776
DAILY|8777,8782
<EOL>|8783,8784
15.|8784,8787
Outpatient|8788,8798
Lab|8799,8802
Work|8803,8807
<EOL>|8807,8808
Please|8808,8814
check|8815,8820
chem7|8821,8826
and|8827,8830
CBC|8831,8834
on|8835,8837
_|8838,8839
_|8839,8840
_|8840,8841
and|8842,8845
fax|8846,8849
results|8850,8857
to|8858,8860
:|8860,8861
<EOL>|8861,8862
Name|8862,8866
:|8866,8867
_|8868,8869
_|8869,8870
_|8870,8871
<EOL>|8872,8873
Fax|8873,8876
:|8876,8877
_|8878,8879
_|8879,8880
_|8880,8881
<EOL>|8882,8883
<EOL>|8883,8884
<EOL>|8885,8886
Discharge|8886,8895
Disposition|8896,8907
:|8907,8908
<EOL>|8908,8909
Home|8909,8913
<EOL>|8913,8914
<EOL>|8915,8916
Discharge|8916,8925
Diagnosis|8926,8935
:|8935,8936
<EOL>|8936,8937
Community|8937,8946
Acquired|8947,8955
Pneumonia|8956,8965
<EOL>|8965,8966
Diabetes|8966,8974
Mellitus|8975,8983
Type|8984,8988
2|8989,8990
<EOL>|8990,8991
<EOL>|8991,8992
<EOL>|8993,8994
Discharge|8994,9003
Condition|9004,9013
:|9013,9014
<EOL>|9014,9015
Mental|9015,9021
Status|9022,9028
:|9028,9029
Clear|9030,9035
and|9036,9039
coherent|9040,9048
.|9048,9049
<EOL>|9049,9050
Level|9050,9055
of|9056,9058
Consciousness|9059,9072
:|9072,9073
Alert|9074,9079
and|9080,9083
interactive|9084,9095
.|9095,9096
<EOL>|9096,9097
Activity|9097,9105
Status|9106,9112
:|9112,9113
Ambulatory|9114,9124
-|9125,9126
Independent|9127,9138
.|9138,9139
<EOL>|9139,9140
<EOL>|9140,9141
<EOL>|9142,9143
Discharge|9143,9152
Instructions|9153,9165
:|9165,9166
<EOL>|9166,9167
Dear|9167,9171
Ms.|9172,9175
_|9176,9177
_|9177,9178
_|9178,9179
,|9179,9180
<EOL>|9181,9182
<EOL>|9182,9183
You|9183,9186
were|9187,9191
admitted|9192,9200
to|9201,9203
the|9204,9207
hospital|9208,9216
for|9217,9220
a|9221,9222
pneumonia|9223,9232
.|9232,9233
You|9235,9238
were|9239,9243
<EOL>|9244,9245
started|9245,9252
on|9253,9255
antibiotics|9256,9267
which|9268,9273
you|9274,9277
will|9278,9282
need|9283,9287
to|9288,9290
continue|9291,9299
for|9300,9303
one|9304,9307
<EOL>|9308,9309
more|9309,9313
day|9314,9317
(|9318,9319
as|9319,9321
listed|9322,9328
below|9329,9334
)|9334,9335
.|9335,9336
You|9338,9341
were|9342,9346
also|9347,9351
a|9352,9353
little|9354,9360
bit|9361,9364
<EOL>|9365,9366
dehydrated|9366,9376
when|9377,9381
you|9382,9385
came|9386,9390
in|9391,9393
,|9393,9394
so|9395,9397
you|9398,9401
received|9402,9410
some|9411,9415
IV|9416,9418
fluids|9419,9425
to|9426,9428
<EOL>|9429,9430
help|9430,9434
hydrate|9435,9442
you|9443,9446
.|9446,9447
<EOL>|9448,9449
<EOL>|9449,9450
You|9450,9453
sodium|9454,9460
levels|9461,9467
in|9468,9470
your|9471,9475
blood|9476,9481
were|9482,9486
a|9487,9488
bit|9489,9492
low|9493,9496
.|9496,9497
This|9499,9503
was|9504,9507
most|9508,9512
<EOL>|9513,9514
likely|9514,9520
due|9521,9524
to|9525,9527
the|9528,9531
infection|9532,9541
in|9542,9544
your|9545,9549
lungs|9550,9555
.|9555,9556
As|9558,9560
we|9561,9563
treated|9564,9571
your|9572,9576
<EOL>|9577,9578
pneumonia|9578,9587
,|9587,9588
your|9589,9593
sodium|9594,9600
levels|9601,9607
improved|9608,9616
.|9616,9617
<EOL>|9617,9618
<EOL>|9618,9619
The|9619,9622
following|9623,9632
changes|9633,9640
were|9641,9645
made|9646,9650
to|9651,9653
your|9654,9658
medications|9659,9670
:|9670,9671
<EOL>|9672,9673
-|9673,9674
Please|9675,9681
START|9682,9687
levofloxacin|9688,9700
750mg|9701,9706
daily|9707,9712
for|9713,9716
1|9717,9718
more|9719,9723
day|9724,9727
<EOL>|9727,9728
<EOL>|9728,9729
If|9729,9731
you|9732,9735
begin|9736,9741
to|9742,9744
feel|9745,9749
more|9750,9754
short|9755,9760
of|9761,9763
breath|9764,9770
or|9771,9773
more|9774,9778
sick|9779,9783
,|9783,9784
please|9785,9791
<EOL>|9792,9793
do|9793,9795
n't|9795,9798
hesitate|9799,9807
to|9808,9810
call|9811,9815
your|9816,9820
primary|9821,9828
care|9829,9833
physician|9834,9843
.|9843,9844
<EOL>|9844,9845
<EOL>|9845,9846
Please|9846,9852
follow|9853,9859
up|9860,9862
with|9863,9867
your|9868,9872
primary|9873,9880
care|9881,9885
doctor|9886,9892
on|9893,9895
discharge|9896,9905
as|9906,9908
<EOL>|9909,9910
scheduled|9910,9919
below|9920,9925
.|9925,9926
<EOL>|9926,9927
<EOL>|9927,9928
Please|9928,9934
have|9935,9939
your|9940,9944
labs|9945,9949
checked|9950,9957
before|9958,9964
your|9965,9969
appointment|9970,9981
with|9982,9986
Dr|9987,9989
.|9989,9990
<EOL>|9991,9992
_|9992,9993
_|9993,9994
_|9994,9995
included|9996,10004
below|10005,10010
.|10010,10011
<EOL>|10011,10012
<EOL>|10012,10013
It|10013,10015
was|10016,10019
a|10020,10021
pleasure|10022,10030
taking|10031,10037
care|10038,10042
of|10043,10045
you|10046,10049
,|10049,10050
we|10051,10053
wish|10054,10058
you|10059,10062
all|10063,10066
the|10067,10070
best|10071,10075
!|10075,10076
<EOL>|10076,10077
<EOL>|10078,10079
Followup|10079,10087
Instructions|10088,10100
:|10100,10101
<EOL>|10101,10102
_|10102,10103
_|10103,10104
_|10104,10105
<EOL>|10105,10106

