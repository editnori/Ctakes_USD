 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Chief|276,281
Complaint|282,291
:|291,292
<EOL>|292,293
Shortness|293,302
of|303,305
Breath|306,312
<EOL>|312,313
<EOL>|313,314
<EOL>|315,316
Major|316,321
Surgical|322,330
or|331,333
Invasive|334,342
Procedure|343,352
:|352,353
<EOL>|353,354
N|354,355
/|355,356
A|356,357
<EOL>|357,358
<EOL>|358,359
<EOL>|360,361
History|361,368
of|369,371
Present|372,379
Illness|380,387
:|387,388
<EOL>|388,389
Ms.|389,392
_|393,394
_|394,395
_|395,396
is|397,399
a|400,401
_|402,403
_|403,404
_|404,405
female|406,412
with|413,417
history|418,425
of|426,428
<EOL>|429,430
COPD|430,434
on|435,437
home|438,442
O2|443,445
,|445,446
atrial|447,453
fibrillation|454,466
on|467,469
apixaban|470,478
,|478,479
hypertension|480,492
,|492,493
<EOL>|494,495
CAD|495,498
,|498,499
and|500,503
hyperlipidemia|504,518
who|519,522
presents|523,531
with|532,536
shortness|537,546
of|547,549
breath|550,556
,|556,557
<EOL>|558,559
cough|559,564
,|564,565
and|566,569
wheezing|570,578
for|579,582
one|583,586
day|587,590
.|590,591
<EOL>|591,592
<EOL>|592,593
The|593,596
patient|597,604
reports|605,612
shortness|613,622
of|623,625
breath|626,632
,|632,633
increased|634,643
cough|644,649
<EOL>|650,651
productive|651,661
of|662,664
_|665,666
_|666,667
_|667,668
red|669,672
-|672,673
flected|673,680
sputum|681,687
,|687,688
and|689,692
wheezing|693,701
since|702,707
<EOL>|708,709
yesterday|709,718
evening|719,726
.|726,727
She|729,732
has|733,736
been|737,741
using|742,747
albuterol|748,757
IH|758,760
more|761,765
<EOL>|766,767
frequently|767,777
(|778,779
_|779,780
_|780,781
_|781,782
)|782,783
with|784,788
ipratropium|789,800
nebs|801,805
every|806,811
4|812,813
hours|814,819
with|820,824
<EOL>|825,826
minimal|826,833
relief|834,840
.|840,841
She|842,845
had|846,849
to|850,852
increase|853,861
her|862,865
O2|866,868
flow|869,873
up|874,876
to|877,879
4L|880,882
without|883,890
<EOL>|891,892
significant|892,903
improvement|904,915
.|915,916
She|917,920
was|921,924
currently|925,934
taking|935,941
10mg|942,946
of|947,949
<EOL>|950,951
prednisone|951,961
.|961,962
She|963,966
has|967,970
also|971,975
been|976,980
taking|981,987
tiotropium|988,998
IH|999,1001
,|1001,1002
<EOL>|1003,1004
theophylline|1004,1016
,|1016,1017
advair|1018,1024
IH|1025,1027
at|1028,1030
home|1031,1035
as|1036,1038
prescribed|1039,1049
.|1049,1050
She|1051,1054
denies|1055,1061
sick|1062,1066
<EOL>|1067,1068
contacts|1068,1076
.|1076,1077
She|1078,1081
quit|1082,1086
smoking|1087,1094
approximately|1095,1108
1|1109,1110
month|1111,1116
ago|1117,1120
.|1120,1121
<EOL>|1121,1122
<EOL>|1122,1123
She|1123,1126
reports|1127,1134
an|1135,1137
episode|1138,1145
of|1146,1148
chest|1149,1154
pain|1155,1159
in|1160,1162
waiting|1163,1170
room|1171,1175
while|1176,1181
<EOL>|1182,1183
sitting|1183,1190
down|1191,1195
,|1195,1196
non-exertional|1197,1211
,|1211,1212
resolved|1213,1221
after|1222,1227
2|1228,1229
minutes|1230,1237
.|1237,1238
She|1239,1242
<EOL>|1243,1244
denies|1244,1250
fever|1251,1256
/|1256,1257
chills|1257,1263
,|1263,1264
abdominal|1265,1274
pain|1275,1279
,|1279,1280
nausea|1281,1287
/|1287,1288
vomiting|1288,1296
,|1296,1297
<EOL>|1298,1299
palpitations|1299,1311
,|1311,1312
and|1313,1316
diaphoresis|1317,1328
.|1328,1329
<EOL>|1331,1332
<EOL>|1332,1333
She|1333,1336
was|1337,1340
recently|1341,1349
admitted|1350,1358
from|1359,1363
_|1364,1365
_|1365,1366
_|1366,1367
to|1368,1370
_|1371,1372
_|1372,1373
_|1373,1374
for|1375,1378
dyspnea|1379,1386
that|1387,1391
<EOL>|1392,1393
was|1393,1396
thought|1397,1404
to|1405,1407
be|1408,1410
secondary|1411,1420
to|1421,1423
steroid|1424,1431
taper|1432,1437
for|1438,1441
recent|1442,1448
COPD|1449,1453
<EOL>|1454,1455
exacerbation|1455,1467
with|1468,1472
a|1473,1474
component|1475,1484
of|1485,1487
anxiety|1488,1495
(|1496,1497
not|1497,1500
an|1501,1503
acute|1504,1509
COPD|1510,1514
<EOL>|1515,1516
exacerbation|1516,1528
)|1528,1529
and|1530,1533
was|1534,1537
treated|1538,1545
with|1546,1550
steroids|1551,1559
and|1560,1563
duonebs|1564,1571
but|1572,1575
no|1576,1578
<EOL>|1579,1580
antibiotics|1580,1591
.|1591,1592
She|1593,1596
had|1597,1600
a|1601,1602
CT|1603,1605
that|1606,1610
showed|1611,1617
emphysema|1618,1627
but|1628,1631
no|1632,1634
evidence|1635,1643
<EOL>|1644,1645
of|1645,1647
infection|1648,1657
such|1658,1662
as|1663,1665
_|1666,1667
_|1667,1668
_|1668,1669
.|1669,1670
Pulmonary|1671,1680
was|1681,1684
consulted|1685,1694
and|1695,1698
<EOL>|1699,1700
recommended|1700,1711
increasing|1712,1722
her|1723,1726
Advair|1727,1733
dose|1734,1738
to|1739,1741
500|1742,1745
/|1745,1746
50|1746,1748
(|1749,1750
which|1750,1755
was|1756,1759
<EOL>|1760,1761
done|1761,1765
)|1765,1766
and|1767,1770
switching|1771,1780
from|1781,1785
theophylline|1786,1798
to|1799,1801
<EOL>|1802,1803
roflumilast|1803,1814
and|1815,1818
initiation|1819,1829
of|1830,1832
long|1833,1837
-|1837,1838
term|1838,1842
azithromycin|1843,1855
therapy|1856,1863
<EOL>|1864,1865
(|1865,1866
which|1866,1871
was|1872,1875
deferred|1876,1884
for|1885,1888
outpatient|1889,1899
follow|1900,1906
-|1906,1907
up|1907,1909
)|1909,1910
She|1911,1914
was|1915,1918
initiated|1919,1928
<EOL>|1929,1930
on|1930,1932
a|1933,1934
steroid|1935,1942
<EOL>|1943,1944
taper|1944,1949
on|1950,1952
_|1953,1954
_|1954,1955
_|1955,1956
of|1957,1959
prednisone|1960,1970
30|1971,1973
mg|1974,1976
for|1977,1980
3|1981,1982
days|1983,1987
,|1987,1988
then|1989,1993
20|1994,1996
mg|1997,1999
for|2000,2003
3|2004,2005
<EOL>|2006,2007
days|2007,2011
,|2011,2012
then|2013,2017
10|2018,2020
mg|2021,2023
until|2024,2029
outpatient|2030,2040
follow|2041,2047
-|2047,2048
up|2048,2050
.|2050,2051
<EOL>|2051,2052
<EOL>|2052,2053
In|2053,2055
the|2056,2059
ED|2060,2062
,|2062,2063
initial|2064,2071
vital|2072,2077
signs|2078,2083
were|2084,2088
:|2088,2089
97.6|2090,2094
67|2095,2097
132|2098,2101
/|2101,2102
82|2102,2104
22|2105,2107
97|2108,2110
%|2110,2111
4L|2112,2114
.|2114,2115
<EOL>|2116,2117
Exam|2117,2121
was|2122,2125
notable|2126,2133
for|2134,2137
limited|2138,2145
air|2146,2149
movement|2150,2158
with|2159,2163
wheezing|2164,2172
<EOL>|2173,2174
bilaterally|2174,2185
.|2185,2186
Labs|2187,2191
were|2192,2196
notable|2197,2204
for|2205,2208
WBC|2209,2212
7.1|2213,2216
,|2216,2217
H|2218,2219
/|2219,2220
H|2220,2221
12.8|2222,2226
/|2226,2227
41|2227,2229
.|2229,2230
1|2230,2231
,|2231,2232
Plt|2233,2236
<EOL>|2237,2238
233|2238,2241
,|2241,2242
Na|2243,2245
133|2246,2249
,|2249,2250
K|2251,2252
3.6|2253,2256
,|2256,2257
BUN|2258,2261
/|2261,2262
Cr|2262,2264
_|2265,2266
_|2266,2267
_|2267,2268
,|2268,2269
trop|2270,2274
<|2275,2276
0.01|2277,2281
,|2281,2282
BNP|2283,2286
181|2287,2290
,|2290,2291
lactate|2292,2299
<EOL>|2300,2301
1.5|2301,2304
,|2304,2305
VBG|2306,2309
7.43|2310,2314
/|2314,2315
_|2315,2316
_|2316,2317
_|2317,2318
.|2318,2319
Imaging|2320,2327
with|2328,2332
CXR|2333,2336
showed|2337,2343
mild|2344,2348
basilar|2349,2356
<EOL>|2357,2358
atelectasis|2358,2369
without|2370,2377
definite|2378,2386
focal|2387,2392
consolidation|2393,2406
.|2406,2407
The|2408,2411
patient|2412,2419
<EOL>|2420,2421
was|2421,2424
given|2425,2430
Duonebs|2431,2438
and|2439,2442
solumedrol|2443,2453
125mg|2454,2459
IV|2460,2462
.|2462,2463
Vitals|2464,2470
prior|2471,2476
to|2477,2479
<EOL>|2480,2481
transfer|2481,2489
were|2490,2494
:|2494,2495
<EOL>|2495,2496
<EOL>|2496,2497
Upon|2497,2501
arrival|2502,2509
to|2510,2512
the|2513,2516
floor|2517,2522
,|2522,2523
she|2524,2527
reports|2528,2535
her|2536,2539
breathing|2540,2549
is|2550,2552
<EOL>|2553,2554
improved|2554,2562
.|2562,2563
<EOL>|2563,2564
<EOL>|2564,2565
REVIEW|2565,2571
OF|2572,2574
SYSTEMS|2575,2582
:|2582,2583
Per|2584,2587
HPI|2588,2591
.|2591,2592
Denies|2593,2599
headache|2600,2608
,|2608,2609
visual|2610,2616
changes|2617,2624
,|2624,2625
<EOL>|2626,2627
pharyngitis|2627,2638
,|2638,2639
rhinorrhea|2640,2650
,|2650,2651
nasal|2652,2657
congestion|2658,2668
,|2668,2669
fevers|2670,2676
,|2676,2677
chills|2678,2684
,|2684,2685
<EOL>|2686,2687
sweats|2687,2693
,|2693,2694
weight|2695,2701
loss|2702,2706
,|2706,2707
abdominal|2708,2717
pain|2718,2722
,|2722,2723
nausea|2724,2730
,|2730,2731
vomiting|2732,2740
,|2740,2741
diarrhea|2742,2750
,|2750,2751
<EOL>|2752,2753
constipation|2753,2765
,|2765,2766
hematochezia|2767,2779
,|2779,2780
dysuria|2781,2788
,|2788,2789
rash|2790,2794
,|2794,2795
paresthesias|2796,2808
,|2808,2809
and|2810,2813
<EOL>|2814,2815
weakness|2815,2823
.|2823,2824
<EOL>|2824,2825
<EOL>|2826,2827
Past|2827,2831
Medical|2832,2839
History|2840,2847
:|2847,2848
<EOL>|2848,2849
-|2849,2850
COPD|2851,2855
/|2855,2856
Asthma|2856,2862
on|2863,2865
home|2866,2870
2L|2871,2873
O2|2874,2876
<EOL>|2876,2877
-|2877,2878
Atypical|2879,2887
Chest|2888,2893
Pain|2894,2898
<EOL>|2898,2899
-|2899,2900
Hypertension|2901,2913
<EOL>|2913,2914
-|2914,2915
Hyperlipidemia|2916,2930
<EOL>|2930,2931
-|2931,2932
Osteroarthritis|2933,2948
<EOL>|2948,2949
-|2949,2950
Atrial|2951,2957
Fibrillation|2958,2970
on|2971,2973
Apixaban|2974,2982
<EOL>|2982,2983
-|2983,2984
Anxiety|2985,2992
<EOL>|2992,2993
-|2993,2994
Cervical|2995,3003
Radiculitis|3004,3015
<EOL>|3015,3016
-|3016,3017
Cervical|3018,3026
Spondylosis|3027,3038
<EOL>|3038,3039
-|3039,3040
Coronary|3041,3049
Artery|3050,3056
Disease|3057,3064
<EOL>|3064,3065
-|3065,3066
Headache|3067,3075
<EOL>|3075,3076
-|3076,3077
Herpes|3078,3084
Zoster|3085,3091
<EOL>|3091,3092
-|3092,3093
GI|3094,3096
Bleeding|3097,3105
<EOL>|3105,3106
-|3106,3107
Peripheral|3108,3118
Vascular|3119,3127
Disease|3128,3135
s|3136,3137
/|3137,3138
p|3138,3139
bilateral|3140,3149
iliac|3150,3155
stents|3156,3162
<EOL>|3162,3163
-|3163,3164
s|3165,3166
/|3166,3167
p|3167,3168
hip|3169,3172
replacement|3173,3184
<EOL>|3184,3185
<EOL>|3186,3187
Social|3187,3193
History|3194,3201
:|3201,3202
<EOL>|3202,3203
_|3203,3204
_|3204,3205
_|3205,3206
<EOL>|3206,3207
Family|3207,3213
History|3214,3221
:|3221,3222
<EOL>|3222,3223
Mother|3223,3229
with|3230,3234
asthma|3235,3241
and|3242,3245
hypertension|3246,3258
.|3258,3259
Father|3260,3266
with|3267,3271
colon|3272,3277
cancer|3278,3284
.|3284,3285
<EOL>|3286,3287
Brother|3287,3294
with|3295,3299
leukemia|3300,3308
.|3308,3309
<EOL>|3309,3310
<EOL>|3310,3311
<EOL>|3312,3313
Physical|3313,3321
Exam|3322,3326
:|3326,3327
<EOL>|3327,3328
ADMISSION|3328,3337
PHYSICAL|3338,3346
EXAM|3347,3351
:|3351,3352
<EOL>|3352,3353
=|3353,3354
=|3354,3355
=|3355,3356
=|3356,3357
=|3357,3358
=|3358,3359
=|3359,3360
=|3360,3361
=|3361,3362
=|3362,3363
=|3363,3364
=|3364,3365
=|3365,3366
=|3366,3367
=|3367,3368
=|3368,3369
=|3369,3370
=|3370,3371
=|3371,3372
=|3372,3373
=|3373,3374
=|3374,3375
=|3375,3376
=|3376,3377
=|3377,3378
=|3378,3379
<EOL>|3379,3380
VITALS|3380,3386
:|3386,3387
Temp|3388,3392
97.3|3393,3397
,|3397,3398
HR|3399,3401
76|3402,3404
,|3404,3405
O2|3406,3408
sat|3409,3412
160|3413,3416
/|3416,3417
80|3417,3419
,|3419,3420
RR|3421,3423
20|3424,3426
,|3426,3427
O2|3428,3430
sat|3431,3434
94|3435,3437
%|3437,3438
4L|3439,3441
<EOL>|3441,3442
GENERAL|3442,3449
:|3449,3450
AOx3|3451,3455
,|3455,3456
speaking|3457,3465
in|3466,3468
full|3469,3473
sentences|3474,3483
,|3483,3484
NAD|3485,3488
,|3488,3489
resting|3490,3497
in|3498,3500
bed|3501,3504
<EOL>|3505,3506
comfortably|3506,3517
.|3517,3518
<EOL>|3518,3519
HEENT|3519,3524
:|3524,3525
NCAT|3526,3530
.|3530,3531
PERRL|3532,3537
.|3537,3538
EOMI|3539,3543
.|3543,3544
Sclera|3545,3551
anicteric|3552,3561
and|3562,3565
not|3566,3569
injected|3570,3578
.|3578,3579
<EOL>|3580,3581
MMM|3581,3584
.|3584,3585
Oropharynx|3586,3596
is|3597,3599
clear|3600,3605
.|3605,3606
<EOL>|3606,3607
NECK|3607,3611
:|3611,3612
Supple|3613,3619
.|3619,3620
No|3621,3623
LAD|3624,3627
.|3627,3628
JVP|3629,3632
not|3633,3636
appreciated|3637,3648
at|3649,3651
45|3652,3654
degrees|3655,3662
.|3662,3663
<EOL>|3663,3664
CARDIAC|3664,3671
:|3671,3672
Irregularly|3673,3684
irregular|3685,3694
,|3694,3695
normal|3696,3702
rate|3703,3707
.|3707,3708
_|3709,3710
_|3710,3711
_|3711,3712
systolic|3713,3721
murmur|3722,3728
<EOL>|3729,3730
<EOL>|3730,3731
at|3731,3733
the|3734,3737
RUSB|3738,3742
.|3742,3743
No|3744,3746
rubs|3747,3751
or|3752,3754
gallops|3755,3762
.|3762,3763
<EOL>|3763,3764
LUNGS|3764,3769
:|3769,3770
Expiratory|3771,3781
wheezes|3782,3789
throughout|3790,3800
with|3801,3805
poor|3806,3810
air|3811,3814
movement|3815,3823
.|3823,3824
<EOL>|3824,3825
ABDOMEN|3825,3832
:|3832,3833
+|3834,3835
BS|3835,3837
,|3837,3838
soft|3839,3843
,|3843,3844
nontender|3845,3854
,|3854,3855
and|3856,3859
nondistended|3860,3872
.|3872,3873
<EOL>|3873,3874
EXTREMITIES|3874,3885
:|3885,3886
Warm|3887,3891
and|3892,3895
well|3896,3900
-|3900,3901
perfused|3901,3909
.|3909,3910
No|3911,3913
edema|3914,3919
.|3919,3920
2|3921,3922
+|3922,3923
DP|3924,3926
pulses|3927,3933
<EOL>|3934,3935
bilaterally|3935,3946
.|3946,3947
<EOL>|3948,3949
NEUROLOGIC|3949,3959
:|3959,3960
A|3961,3962
&|3962,3963
Ox3|3963,3966
,|3966,3967
CNII|3968,3972
-|3972,3973
XII|3973,3976
intact|3977,3983
,|3983,3984
strength|3985,3993
and|3994,3997
sensation|3998,4007
<EOL>|4008,4009
grossly|4009,4016
intact|4017,4023
bilaterally|4024,4035
.|4035,4036
<EOL>|4036,4037
<EOL>|4037,4038
DISCHARGE|4038,4047
PHYSICAL|4048,4056
EXAM|4057,4061
:|4061,4062
<EOL>|4062,4063
=|4063,4064
=|4064,4065
=|4065,4066
=|4066,4067
=|4067,4068
=|4068,4069
=|4069,4070
=|4070,4071
=|4071,4072
=|4072,4073
=|4073,4074
=|4074,4075
=|4075,4076
=|4076,4077
=|4077,4078
=|4078,4079
=|4079,4080
=|4080,4081
=|4081,4082
=|4082,4083
=|4083,4084
=|4084,4085
=|4085,4086
=|4086,4087
=|4087,4088
=|4088,4089
=|4089,4090
<EOL>|4090,4091
VITALS|4091,4097
:|4097,4098
Tm|4099,4101
99.1|4102,4106
,|4106,4107
146|4108,4111
/|4111,4112
69|4112,4114
(|4115,4116
143|4116,4119
-|4119,4120
159|4120,4123
/|4123,4124
69|4124,4126
-|4126,4127
77|4127,4129
)|4129,4130
,|4130,4131
94|4132,4134
,|4134,4135
22|4136,4138
,|4138,4139
94|4140,4142
-|4142,4143
95|4143,4145
%|4145,4146
%|4146,4147
2L|4148,4150
<EOL>|4150,4151
GENERAL|4151,4158
:|4158,4159
speaking|4160,4168
in|4169,4171
full|4172,4176
sentences|4177,4186
,|4186,4187
NAD|4188,4191
,|4191,4192
resting|4193,4200
in|4201,4203
bed|4204,4207
<EOL>|4208,4209
comfortably|4209,4220
.|4220,4221
<EOL>|4221,4222
CARDIAC|4222,4229
:|4229,4230
rrr|4231,4234
,|4234,4235
normal|4236,4242
rate|4243,4247
.|4247,4248
_|4249,4250
_|4250,4251
_|4251,4252
systolic|4253,4261
murmur|4262,4268
at|4269,4271
the|4272,4275
RUSB|4276,4280
<EOL>|4280,4281
LUNGS|4281,4286
:|4286,4287
+|4288,4289
mild|4289,4293
wheezes|4294,4301
throughout|4302,4312
<EOL>|4312,4313
ABDOMEN|4313,4320
:|4320,4321
+|4322,4323
BS|4323,4325
,|4325,4326
soft|4327,4331
,|4331,4332
nontender|4333,4342
,|4342,4343
and|4344,4347
nondistended|4348,4360
.|4360,4361
<EOL>|4361,4362
EXTREMITIES|4362,4373
:|4373,4374
Warm|4375,4379
and|4380,4383
well|4384,4388
-|4388,4389
perfused|4389,4397
.|4397,4398
1|4399,4400
+|4400,4401
b|4402,4403
/|4403,4404
l|4404,4405
_|4406,4407
_|4407,4408
_|4408,4409
edema|4410,4415
.|4415,4416
<EOL>|4417,4418
NEUROLOGIC|4418,4428
:|4428,4429
grossly|4430,4437
nonfocal|4438,4446
,|4446,4447
aaox3|4448,4453
<EOL>|4453,4454
<EOL>|4455,4456
Pertinent|4456,4465
Results|4466,4473
:|4473,4474
<EOL>|4474,4475
ADMISSION|4475,4484
LABS|4485,4489
:|4489,4490
<EOL>|4491,4492
=|4492,4493
=|4493,4494
=|4494,4495
=|4495,4496
=|4496,4497
=|4497,4498
=|4498,4499
=|4499,4500
=|4500,4501
=|4501,4502
=|4502,4503
=|4503,4504
=|4504,4505
=|4505,4506
=|4506,4507
=|4507,4508
=|4508,4509
=|4509,4510
=|4510,4511
=|4511,4512
=|4512,4513
=|4513,4514
=|4514,4515
=|4515,4516
=|4516,4517
<EOL>|4517,4518
_|4518,4519
_|4519,4520
_|4520,4521
05|4522,4524
:|4524,4525
54PM|4525,4529
BLOOD|4530,4535
WBC|4536,4539
-|4539,4540
7.1|4540,4543
RBC|4544,4547
-|4547,4548
4|4548,4549
.|4549,4550
74|4550,4552
Hgb|4553,4556
-|4556,4557
12.8|4557,4561
Hct|4562,4565
-|4565,4566
41.1|4566,4570
MCV|4571,4574
-|4574,4575
87|4575,4577
<EOL>|4578,4579
MCH|4579,4582
-|4582,4583
27.0|4583,4587
MCHC|4588,4592
-|4592,4593
31|4593,4595
.|4595,4596
1|4596,4597
*|4597,4598
RDW|4599,4602
-|4602,4603
22|4603,4605
.|4605,4606
6|4606,4607
*|4607,4608
RDWSD|4609,4614
-|4614,4615
69|4615,4617
.|4617,4618
0|4618,4619
*|4619,4620
Plt|4621,4624
_|4625,4626
_|4626,4627
_|4627,4628
<EOL>|4628,4629
_|4629,4630
_|4630,4631
_|4631,4632
05|4633,4635
:|4635,4636
54PM|4636,4640
BLOOD|4641,4646
Neuts|4647,4652
-|4652,4653
81|4653,4655
.|4655,4656
8|4656,4657
*|4657,4658
Lymphs|4659,4665
-|4665,4666
9|4666,4667
.|4667,4668
6|4668,4669
*|4669,4670
Monos|4671,4676
-|4676,4677
7.6|4677,4680
<EOL>|4681,4682
Eos|4682,4685
-|4685,4686
0|4686,4687
.|4687,4688
3|4688,4689
*|4689,4690
Baso|4691,4695
-|4695,4696
0.1|4696,4699
Im|4700,4702
_|4703,4704
_|4704,4705
_|4705,4706
AbsNeut|4707,4714
-|4714,4715
5|4715,4716
.|4716,4717
82|4717,4719
AbsLymp|4720,4727
-|4727,4728
0|4728,4729
.|4729,4730
68|4730,4732
*|4732,4733
<EOL>|4734,4735
AbsMono|4735,4742
-|4742,4743
0|4743,4744
.|4744,4745
54|4745,4747
AbsEos|4748,4754
-|4754,4755
0|4755,4756
.|4756,4757
02|4757,4759
*|4759,4760
AbsBaso|4761,4768
-|4768,4769
0.01|4769,4773
<EOL>|4773,4774
_|4774,4775
_|4775,4776
_|4776,4777
06|4778,4780
:|4780,4781
35AM|4781,4785
BLOOD|4786,4791
Calcium|4792,4799
-|4799,4800
9.9|4800,4803
Phos|4804,4808
-|4808,4809
4.1|4809,4812
Mg|4813,4815
-|4815,4816
2.0|4816,4819
<EOL>|4819,4820
_|4820,4821
_|4821,4822
_|4822,4823
05|4824,4826
:|4826,4827
54PM|4827,4831
BLOOD|4832,4837
_|4838,4839
_|4839,4840
_|4840,4841
pO2|4842,4845
-|4845,4846
52|4846,4848
*|4848,4849
pCO2|4850,4854
-|4854,4855
49|4855,4857
*|4857,4858
pH|4859,4861
-|4861,4862
7.43|4862,4866
<EOL>|4867,4868
calTCO2|4868,4875
-|4875,4876
34|4876,4878
*|4878,4879
Base|4880,4884
XS|4885,4887
-|4887,4888
6|4888,4889
<EOL>|4889,4890
_|4890,4891
_|4891,4892
_|4892,4893
05|4894,4896
:|4896,4897
54PM|4897,4901
BLOOD|4902,4907
Lactate|4908,4915
-|4915,4916
1.5|4916,4919
<EOL>|4919,4920
_|4920,4921
_|4921,4922
_|4922,4923
05|4924,4926
:|4926,4927
54PM|4927,4931
BLOOD|4932,4937
proBNP|4938,4944
-|4944,4945
181|4945,4948
<EOL>|4948,4949
_|4949,4950
_|4950,4951
_|4951,4952
05|4953,4955
:|4955,4956
54PM|4956,4960
BLOOD|4961,4966
cTropnT|4967,4974
-|4974,4975
<|4975,4976
0|4976,4977
.|4977,4978
01|4978,4980
<EOL>|4980,4981
<EOL>|4981,4982
STUDIES|4982,4989
:|4989,4990
<EOL>|4991,4992
=|4992,4993
=|4993,4994
=|4994,4995
=|4995,4996
=|4996,4997
=|4997,4998
=|4998,4999
=|4999,5000
=|5000,5001
=|5001,5002
=|5002,5003
=|5003,5004
=|5004,5005
=|5005,5006
=|5006,5007
=|5007,5008
=|5008,5009
=|5009,5010
=|5010,5011
=|5011,5012
=|5012,5013
=|5013,5014
=|5014,5015
=|5015,5016
=|5016,5017
<EOL>|5017,5018
+|5018,5019
CXR|5020,5023
(|5024,5025
_|5025,5026
_|5026,5027
_|5027,5028
)|5028,5029
:|5029,5030
Mild|5031,5035
basilar|5036,5043
atelectasis|5044,5055
without|5056,5063
definite|5064,5072
focal|5073,5078
<EOL>|5079,5080
consolidation|5080,5093
.|5093,5094
<EOL>|5094,5095
+|5095,5096
EKG|5097,5100
:|5100,5101
Sinus|5102,5107
rhythm|5108,5114
at|5115,5117
69|5118,5120
,|5120,5121
left|5122,5126
bundle|5127,5133
branch|5134,5140
block|5141,5146
,|5146,5147
no|5148,5150
acute|5151,5156
ST|5157,5159
<EOL>|5160,5161
or|5161,5163
T|5164,5165
wave|5166,5170
changes|5171,5178
.|5178,5179
<EOL>|5179,5180
<EOL>|5180,5181
DISCHARGE|5181,5190
LABS|5191,5195
:|5195,5196
<EOL>|5197,5198
=|5198,5199
=|5199,5200
=|5200,5201
=|5201,5202
=|5202,5203
=|5203,5204
=|5204,5205
=|5205,5206
=|5206,5207
=|5207,5208
=|5208,5209
=|5209,5210
=|5210,5211
=|5211,5212
=|5212,5213
=|5213,5214
=|5214,5215
=|5215,5216
=|5216,5217
=|5217,5218
=|5218,5219
=|5219,5220
=|5220,5221
=|5221,5222
=|5222,5223
<EOL>|5223,5224
_|5224,5225
_|5225,5226
_|5226,5227
06|5228,5230
:|5230,5231
38AM|5231,5235
BLOOD|5236,5241
WBC|5242,5245
-|5245,5246
14|5246,5248
.|5248,5249
4|5249,5250
*|5250,5251
#|5251,5252
RBC|5253,5256
-|5256,5257
4|5257,5258
.|5258,5259
34|5259,5261
Hgb|5262,5265
-|5265,5266
11.8|5266,5270
Hct|5271,5274
-|5274,5275
37.6|5275,5279
<EOL>|5280,5281
MCV|5281,5284
-|5284,5285
87|5285,5287
MCH|5288,5291
-|5291,5292
27.2|5292,5296
MCHC|5297,5301
-|5301,5302
31|5302,5304
.|5304,5305
4|5305,5306
*|5306,5307
RDW|5308,5311
-|5311,5312
22|5312,5314
.|5314,5315
5|5315,5316
*|5316,5317
RDWSD|5318,5323
-|5323,5324
69|5324,5326
.|5326,5327
4|5327,5328
*|5328,5329
Plt|5330,5333
_|5334,5335
_|5335,5336
_|5336,5337
<EOL>|5337,5338
_|5338,5339
_|5339,5340
_|5340,5341
06|5342,5344
:|5344,5345
38AM|5345,5349
BLOOD|5350,5355
Glucose|5356,5363
-|5363,5364
113|5364,5367
*|5367,5368
UreaN|5369,5374
-|5374,5375
18|5375,5377
Creat|5378,5383
-|5383,5384
0.8|5384,5387
Na|5388,5390
-|5390,5391
137|5391,5394
<EOL>|5395,5396
K|5396,5397
-|5397,5398
3.1|5398,5401
(|5401,5402
repleted|5402,5410
)|5410,5411
*|5411,5412
Cl|5413,5415
-|5415,5416
94|5416,5418
*|5418,5419
HCO3|5420,5424
-|5424,5425
31|5425,5427
AnGap|5428,5433
-|5433,5434
15|5434,5436
<EOL>|5436,5437
<EOL>|5437,5438
<EOL>|5439,5440
Brief|5440,5445
Hospital|5446,5454
Course|5455,5461
:|5461,5462
<EOL>|5462,5463
Ms.|5463,5466
_|5467,5468
_|5468,5469
_|5469,5470
is|5471,5473
a|5474,5475
_|5476,5477
_|5477,5478
_|5478,5479
female|5480,5486
with|5487,5491
history|5492,5499
of|5500,5502
<EOL>|5503,5504
COPD|5504,5508
on|5509,5511
home|5512,5516
O2|5517,5519
,|5519,5520
atrial|5521,5527
fibrillation|5528,5540
on|5541,5543
apixaban|5544,5552
,|5552,5553
hypertension|5554,5566
,|5566,5567
<EOL>|5568,5569
CAD|5569,5572
,|5572,5573
and|5574,5577
hyperlipidemia|5578,5592
who|5593,5596
presents|5597,5605
with|5606,5610
shortness|5611,5620
of|5621,5623
breath|5624,5630
,|5630,5631
<EOL>|5632,5633
cough|5633,5638
,|5638,5639
and|5640,5643
wheezing|5644,5652
for|5653,5656
one|5657,5660
day|5661,5664
.|5664,5665
Pt|5666,5668
recently|5669,5677
DC|5678,5680
'd|5680,5682
from|5683,5687
hospital|5688,5696
<EOL>|5697,5698
for|5698,5701
dyspnea|5702,5709
,|5709,5710
treated|5711,5718
only|5719,5723
w|5724,5725
/|5725,5726
nebs|5726,5730
and|5731,5734
steroids|5735,5743
as|5744,5746
not|5747,5750
thought|5751,5758
_|5759,5760
_|5760,5761
_|5761,5762
<EOL>|5763,5764
true|5764,5768
COPD|5769,5773
exacerbation|5774,5786
,|5786,5787
c|5788,5789
/|5789,5790
f|5790,5791
anxiety|5792,5799
component|5800,5809
.|5809,5810
Pt|5811,5813
re-admitted|5814,5825
<EOL>|5826,5827
w|5827,5828
/|5828,5829
similar|5829,5836
Sx|5837,5839
,|5839,5840
thought|5841,5848
_|5849,5850
_|5850,5851
_|5851,5852
COPD|5853,5857
exacerbation|5858,5870
,|5870,5871
received|5872,5880
nebs|5881,5885
,|5885,5886
<EOL>|5887,5888
steroids|5888,5896
,|5896,5897
azithromycin|5898,5910
.|5910,5911
Pt|5912,5914
's|5914,5916
wheezing|5917,5925
,|5925,5926
cough|5927,5932
,|5932,5933
SOB|5934,5937
improved|5938,5946
<EOL>|5947,5948
shortly|5948,5955
after|5956,5961
admission|5962,5971
,|5971,5972
O2|5973,5975
titrated|5976,5984
down|5985,5989
&|5990,5991
satting|5992,5999
well|6000,6004
on|6005,6007
2L|6008,6010
<EOL>|6011,6012
in|6012,6014
mid-90s|6015,6022
which|6023,6028
is|6029,6031
baseline|6032,6040
.|6040,6041
Evaluated|6042,6051
by|6052,6054
_|6055,6056
_|6056,6057
_|6057,6058
,|6058,6059
recommended|6060,6071
DC|6072,6074
to|6075,6077
<EOL>|6078,6079
pulmonary|6079,6088
rehab|6089,6094
,|6094,6095
pt|6096,6098
was|6099,6102
agreeable|6103,6112
.|6112,6113
<EOL>|6114,6115
<EOL>|6115,6116
ACTIVE|6116,6122
ISSUES|6123,6129
<EOL>|6129,6130
=|6130,6131
=|6131,6132
=|6132,6133
=|6133,6134
=|6134,6135
=|6135,6136
=|6136,6137
=|6137,6138
=|6138,6139
=|6139,6140
=|6140,6141
=|6141,6142
=|6142,6143
=|6143,6144
=|6144,6145
=|6145,6146
=|6146,6147
<EOL>|6147,6148
#|6148,6149
Shortness|6150,6159
of|6160,6162
Breath|6163,6169
:|6169,6170
Patient|6171,6178
with|6179,6183
history|6184,6191
of|6192,6194
COPD|6195,6199
and|6200,6203
recent|6204,6210
<EOL>|6211,6212
admission|6212,6221
for|6222,6225
dyspnea|6226,6233
in|6234,6236
the|6237,6240
setting|6241,6248
of|6249,6251
steroid|6252,6259
taper|6260,6265
.|6265,6266
Her|6267,6270
<EOL>|6271,6272
symptoms|6272,6280
on|6281,6283
presentation|6284,6296
were|6297,6301
consistent|6302,6312
with|6313,6317
severe|6318,6324
COPD|6325,6329
given|6330,6335
<EOL>|6336,6337
diffuse|6337,6344
wheezing|6345,6353
and|6354,6357
poor|6358,6362
air|6363,6366
movement|6367,6375
.|6375,6376
She|6377,6380
likely|6381,6387
had|6388,6391
an|6392,6394
<EOL>|6395,6396
exacerbation|6396,6408
in|6409,6411
the|6412,6415
setting|6416,6423
of|6424,6426
a|6427,6428
decrease|6429,6437
in|6438,6440
her|6441,6444
steroids|6445,6453
.|6453,6454
There|6455,6460
<EOL>|6461,6462
may|6462,6465
also|6466,6470
be|6471,6473
a|6474,6475
component|6476,6485
of|6486,6488
anxiety|6489,6496
.|6496,6497
She|6498,6501
underwent|6502,6511
CT|6512,6514
last|6515,6519
<EOL>|6520,6521
admission|6521,6530
that|6531,6535
was|6536,6539
negative|6540,6548
for|6549,6552
infections|6553,6563
such|6564,6568
as|6569,6571
_|6572,6573
_|6573,6574
_|6574,6575
.|6575,6576
She|6577,6580
was|6581,6584
<EOL>|6585,6586
continued|6586,6595
on|6596,6598
home|6599,6603
spiriva|6604,6611
,|6611,6612
theophylline|6613,6625
,|6625,6626
advair|6627,6633
.|6633,6634
She|6635,6638
was|6639,6642
started|6643,6650
<EOL>|6651,6652
on|6652,6654
standing|6655,6663
duonebs|6664,6671
q6h|6672,6675
and|6676,6679
albuterol|6680,6689
q2h|6690,6693
prn|6694,6697
and|6698,6701
prednisone|6702,6712
was|6713,6716
<EOL>|6717,6718
started|6718,6725
at|6726,6728
40mg|6729,6733
daily|6734,6739
with|6740,6744
slow|6745,6749
taper|6750,6755
.|6755,6756
She|6757,6760
was|6761,6764
also|6765,6769
given|6770,6775
<EOL>|6776,6777
azithromycin|6777,6789
to|6790,6792
complete|6793,6801
5|6802,6803
day|6804,6807
course|6808,6814
.|6814,6815
She|6816,6819
had|6820,6823
improvement|6824,6835
in|6836,6838
<EOL>|6839,6840
her|6840,6843
wheezing|6844,6852
and|6853,6856
returned|6857,6865
to|6866,6868
baseline|6869,6877
O2|6878,6880
requirement|6881,6892
after|6893,6898
48|6899,6901
<EOL>|6902,6903
hours|6903,6908
.|6908,6909
She|6910,6913
was|6914,6917
seen|6918,6922
by|6923,6925
_|6926,6927
_|6927,6928
_|6928,6929
who|6930,6933
felt|6934,6938
that|6939,6943
she|6944,6947
would|6948,6953
benefit|6954,6961
from|6962,6966
<EOL>|6967,6968
discharge|6968,6977
to|6978,6980
inpatient|6981,6990
pulmonary|6991,7000
rehabilitation|7001,7015
program|7016,7023
.|7023,7024
On|7025,7027
DC|7028,7030
<EOL>|7031,7032
to|7032,7034
_|7035,7036
_|7036,7037
_|7037,7038
rehab|7039,7044
,|7044,7045
recommended|7046,7057
continued|7058,7067
Prendisone|7068,7078
40mg|7079,7083
<EOL>|7084,7085
daily|7085,7090
for|7091,7094
1x|7095,7097
week|7098,7102
with|7103,7107
slow|7108,7112
taper|7113,7118
by|7119,7121
5mg|7122,7125
every|7126,7131
5|7132,7133
days|7134,7138
.|7138,7139
_|7140,7141
_|7141,7142
_|7142,7143
also|7144,7148
<EOL>|7149,7150
consider|7150,7158
starting|7159,7167
bactrim|7168,7175
ppx|7176,7179
with|7180,7184
extended|7185,7193
duration|7194,7202
of|7203,7205
steroids|7206,7214
<EOL>|7215,7216
if|7216,7218
unable|7219,7225
to|7226,7228
wean|7229,7233
less|7234,7238
than|7239,7243
20mg|7244,7248
qd|7249,7251
.|7251,7252
Will|7253,7257
also|7258,7262
f|7263,7264
/|7264,7265
u|7265,7266
as|7267,7269
outpatient|7270,7280
<EOL>|7281,7282
with|7282,7286
pulm|7287,7291
.|7291,7292
<EOL>|7292,7293
<EOL>|7293,7294
CHRONIC|7294,7301
ISSUES|7302,7308
:|7308,7309
<EOL>|7310,7311
=|7311,7312
=|7312,7313
=|7313,7314
=|7314,7315
=|7315,7316
=|7316,7317
=|7317,7318
=|7318,7319
=|7319,7320
=|7320,7321
=|7321,7322
=|7322,7323
=|7323,7324
=|7324,7325
=|7325,7326
=|7326,7327
=|7327,7328
=|7328,7329
<EOL>|7329,7330
#|7330,7331
Anxiety|7332,7339
/|7339,7340
Insomnia|7340,7348
:|7348,7349
Continued|7350,7359
home|7360,7364
lorazepam|7365,7374
.|7374,7375
Consider|7376,7384
starting|7385,7393
<EOL>|7394,7395
SRRI|7395,7399
as|7400,7402
an|7403,7405
outpatient|7406,7416
.|7416,7417
<EOL>|7418,7419
#|7419,7420
Atrial|7421,7427
Fibrillation|7428,7440
:|7440,7441
Continued|7442,7451
dilt|7452,7456
for|7457,7460
rate|7461,7465
control|7466,7473
and|7474,7477
<EOL>|7478,7479
apixaban|7479,7487
for|7488,7491
anticoagulation|7492,7507
.|7507,7508
<EOL>|7508,7509
#|7509,7510
Hypertension|7511,7523
:|7523,7524
Continued|7525,7534
home|7535,7539
imdur|7540,7545
,|7545,7546
hydrochlorothiazide|7547,7566
,|7566,7567
and|7568,7571
<EOL>|7572,7573
diltiazem|7573,7582
.|7582,7583
<EOL>|7583,7584
#|7584,7585
CAD|7586,7589
:|7589,7590
Cardiac|7591,7598
catheterization|7599,7614
in|7615,7617
_|7618,7619
_|7619,7620
_|7620,7621
without|7622,7629
evidence|7630,7638
of|7639,7641
<EOL>|7642,7643
significant|7643,7654
stenosis|7655,7663
of|7664,7666
coronaries|7667,7677
.|7677,7678
ECHO|7679,7683
on|7684,7686
_|7687,7688
_|7688,7689
_|7689,7690
with|7691,7695
EF|7696,7698
>|7699,7700
<EOL>|7701,7702
55|7702,7704
%|7704,7705
and|7706,7709
no|7710,7712
regional|7713,7721
or|7722,7724
global|7725,7731
wall|7732,7736
motion|7737,7743
abnormalities|7744,7757
.|7757,7758
<EOL>|7759,7760
Continued|7760,7769
home|7770,7774
aspirin|7775,7782
and|7783,7786
atorvastatin|7787,7799
.|7799,7800
<EOL>|7800,7801
#|7801,7802
Anemia|7803,7809
:|7809,7810
Continued|7811,7820
home|7821,7825
iron|7826,7830
supplements|7831,7842
.|7842,7843
<EOL>|7843,7844
<EOL>|7844,7845
TRANSITIONAL|7845,7857
ISSUES|7858,7864
:|7864,7865
<EOL>|7865,7866
=|7866,7867
=|7867,7868
=|7868,7869
=|7869,7870
=|7870,7871
=|7871,7872
=|7872,7873
=|7873,7874
=|7874,7875
=|7875,7876
=|7876,7877
=|7877,7878
=|7878,7879
=|7879,7880
=|7880,7881
=|7881,7882
=|7882,7883
=|7883,7884
=|7884,7885
=|7885,7886
=|7886,7887
=|7887,7888
=|7888,7889
=|7889,7890
=|7890,7891
=|7891,7892
<EOL>|7892,7893
[|7893,7894
]|7894,7895
For|7896,7899
pt|7900,7902
's|7902,7904
continued|7905,7914
COPD|7915,7919
exacerbations|7920,7933
,|7933,7934
recommend|7935,7944
finishing|7945,7954
5d|7955,7957
<EOL>|7958,7959
course|7959,7965
of|7966,7968
Azithromycin|7969,7981
,|7981,7982
250mg|7983,7988
qd|7989,7991
until|7992,7997
_|7998,7999
_|7999,8000
_|8000,8001
<EOL>|8001,8002
[|8002,8003
]|8003,8004
Recommend|8005,8014
extended|8015,8023
prednisone|8024,8034
taper|8035,8040
for|8041,8044
pt|8045,8047
,|8047,8048
5d|8049,8051
40mg|8052,8056
<EOL>|8057,8058
Prednisone|8058,8068
(|8069,8070
to|8070,8072
finish|8073,8079
_|8080,8081
_|8081,8082
_|8082,8083
followed|8084,8092
by|8093,8095
10mg|8096,8100
taper|8101,8106
every|8107,8112
5|8113,8114
days|8115,8119
<EOL>|8120,8121
(|8121,8122
35mg|8122,8126
from|8127,8131
_|8132,8133
_|8133,8134
_|8134,8135
,|8135,8136
30mg|8137,8141
_|8142,8143
_|8143,8144
_|8144,8145
,|8145,8146
etc|8147,8150
...|8150,8153
)|8153,8154
.|8154,8155
<EOL>|8156,8157
[|8157,8158
]|8158,8159
Would|8160,8165
consider|8166,8174
PCP|8175,8178
prophylaxis|8179,8190
with|8191,8195
_|8196,8197
_|8197,8198
_|8198,8199
if|8200,8202
unable|8203,8209
to|8210,8212
wean|8213,8217
<EOL>|8218,8219
prednisone|8219,8229
to|8230,8232
less|8233,8237
than|8238,8242
20mg|8243,8247
daily|8248,8253
.|8253,8254
<EOL>|8255,8256
[|8256,8257
]|8257,8258
Pt|8259,8261
's|8261,8263
SOB|8264,8267
may|8268,8271
have|8272,8276
an|8277,8279
anxiety|8280,8287
component|8288,8297
,|8297,8298
may|8299,8302
benefit|8303,8310
from|8311,8315
<EOL>|8316,8317
starting|8317,8325
SSRI|8326,8330
in|8331,8333
addition|8334,8342
to|8343,8345
home|8346,8350
benzos|8351,8357
already|8358,8365
prescribed|8366,8376
<EOL>|8376,8377
<EOL>|8377,8378
#|8378,8379
CONTACT|8380,8387
:|8387,8388
Full|8389,8393
Code|8394,8398
<EOL>|8398,8399
#|8399,8400
CODE|8401,8405
STATUS|8406,8412
:|8412,8413
_|8414,8415
_|8415,8416
_|8416,8417
(|8418,8419
husband|8419,8426
/|8426,8427
HCP|8427,8430
)|8430,8431
_|8432,8433
_|8433,8434
_|8434,8435
<EOL>|8435,8436
<EOL>|8437,8438
_|8438,8439
_|8439,8440
_|8440,8441
on|8442,8444
Admission|8445,8454
:|8454,8455
<EOL>|8455,8456
The|8456,8459
Preadmission|8460,8472
Medication|8473,8483
list|8484,8488
is|8489,8491
accurate|8492,8500
and|8501,8504
complete|8505,8513
.|8513,8514
<EOL>|8514,8515
1.|8515,8517
Acetaminophen|8518,8531
325|8532,8535
mg|8536,8538
PO|8539,8541
Q4H|8542,8545
:|8545,8546
PRN|8546,8549
Pain|8550,8554
<EOL>|8555,8556
2.|8556,8558
Apixaban|8559,8567
5|8568,8569
mg|8570,8572
PO|8573,8575
BID|8576,8579
<EOL>|8580,8581
3.|8581,8583
Aspirin|8584,8591
81|8592,8594
mg|8595,8597
PO|8598,8600
DAILY|8601,8606
<EOL>|8607,8608
4.|8608,8610
Atorvastatin|8611,8623
10|8624,8626
mg|8627,8629
PO|8630,8632
QPM|8633,8636
<EOL>|8637,8638
5.|8638,8640
Diltiazem|8641,8650
Extended|8651,8659
-|8659,8660
Release|8660,8667
240|8668,8671
mg|8672,8674
PO|8675,8677
BID|8678,8681
<EOL>|8682,8683
6.|8683,8685
Docusate|8686,8694
Sodium|8695,8701
100|8702,8705
mg|8706,8708
PO|8709,8711
BID|8712,8715
<EOL>|8716,8717
7.|8717,8719
Dorzolamide|8720,8731
2|8732,8733
%|8733,8734
Ophth|8735,8740
.|8740,8741
Soln.|8742,8747
1|8748,8749
DROP|8750,8754
BOTH|8755,8759
EYES|8760,8764
BID|8765,8768
<EOL>|8769,8770
8.|8770,8772
Ferrous|8773,8780
Sulfate|8781,8788
325|8789,8792
mg|8793,8795
PO|8796,8798
DAILY|8799,8804
<EOL>|8805,8806
9.|8806,8808
Fluticasone|8809,8820
Propionate|8821,8831
NASAL|8832,8837
2|8838,8839
SPRY|8840,8844
NU|8845,8847
DAILY|8848,8853
:|8853,8854
PRN|8854,8857
allergies|8858,8867
<EOL>|8868,8869
10.|8869,8872
Hydrochlorothiazide|8873,8892
50|8893,8895
mg|8896,8898
PO|8899,8901
DAILY|8902,8907
<EOL>|8908,8909
11.|8909,8912
Isosorbide|8913,8923
Mononitrate|8924,8935
(|8936,8937
Extended|8937,8945
Release|8946,8953
)|8953,8954
240|8955,8958
mg|8959,8961
PO|8962,8964
DAILY|8965,8970
<EOL>|8971,8972
12.|8972,8975
Latanoprost|8976,8987
0.005|8988,8993
%|8993,8994
Ophth|8995,9000
.|9000,9001
Soln.|9002,9007
1|9008,9009
DROP|9010,9014
BOTH|9015,9019
EYES|9020,9024
QHS|9025,9028
<EOL>|9029,9030
13.|9030,9033
Multivitamins|9034,9047
1|9048,9049
TAB|9050,9053
PO|9054,9056
DAILY|9057,9062
<EOL>|9063,9064
14.|9064,9067
PredniSONE|9068,9078
10|9079,9081
mg|9082,9084
PO|9085,9087
DAILY|9088,9093
<EOL>|9094,9095
15.|9095,9098
Ranitidine|9099,9109
300|9110,9113
mg|9114,9116
PO|9117,9119
DAILY|9120,9125
<EOL>|9126,9127
16|9127,9129
.|9129,9130
Theophylline|9131,9143
SR|9144,9146
300|9147,9150
mg|9151,9153
PO|9154,9156
BID|9157,9160
<EOL>|9161,9162
17.|9162,9165
Tiotropium|9166,9176
Bromide|9177,9184
1|9185,9186
CAP|9187,9190
IH|9191,9193
DAILY|9194,9199
<EOL>|9200,9201
18.|9201,9204
Ipratropium|9205,9216
Bromide|9217,9224
Neb|9225,9228
1|9229,9230
NEB|9231,9234
IH|9235,9237
Q6H|9238,9241
:|9241,9242
PRN|9242,9245
Wheezing|9246,9254
<EOL>|9255,9256
19.|9256,9259
cod|9260,9263
liver|9264,9269
oil|9270,9273
1|9274,9275
capsule|9276,9283
oral|9285,9289
BID|9290,9293
<EOL>|9294,9295
20|9295,9297
.|9297,9298
Calcitrate|9299,9309
-|9309,9310
Vitamin|9310,9317
D|9318,9319
(|9320,9321
calcium|9321,9328
citrate|9329,9336
-|9336,9337
vitamin|9337,9344
D3|9345,9347
)|9347,9348
315|9349,9352
mg|9353,9355
-|9356,9357
<EOL>|9358,9359
200|9359,9362
units|9363,9368
oral|9370,9374
DAILY|9375,9380
<EOL>|9381,9382
21.|9382,9385
albuterol|9386,9395
sulfate|9396,9403
90|9404,9406
mcg|9407,9410
/|9410,9411
actuation|9411,9420
inhalation|9421,9431
Q4H|9432,9435
<EOL>|9436,9437
22.|9437,9440
Fluticasone|9441,9452
-|9452,9453
Salmeterol|9453,9463
Diskus|9464,9470
(|9471,9472
500|9472,9475
/|9475,9476
50|9476,9478
)|9478,9479
1|9481,9482
INH|9483,9486
IH|9487,9489
BID|9490,9493
<EOL>|9494,9495
23|9495,9497
.|9497,9498
Lorazepam|9499,9508
0.5|9509,9512
mg|9513,9515
PO|9516,9518
Q8H|9519,9522
:|9522,9523
PRN|9523,9526
Anxiety|9527,9534
<EOL>|9535,9536
24|9536,9538
.|9538,9539
Guaifenesin|9540,9551
_|9552,9553
_|9553,9554
_|9554,9555
mL|9556,9558
PO|9559,9561
Q4H|9562,9565
:|9565,9566
PRN|9566,9569
cough|9570,9575
<EOL>|9576,9577
<EOL>|9577,9578
<EOL>|9579,9580
Discharge|9580,9589
Medications|9590,9601
:|9601,9602
<EOL>|9602,9603
1.|9603,9605
Acetaminophen|9606,9619
325|9620,9623
mg|9624,9626
PO|9627,9629
Q4H|9630,9633
:|9633,9634
PRN|9634,9637
Pain|9638,9642
<EOL>|9643,9644
2.|9644,9646
albuterol|9647,9656
sulfate|9657,9664
90|9665,9667
mcg|9668,9671
/|9671,9672
actuation|9672,9681
inhalation|9682,9692
Q4H|9693,9696
<EOL>|9697,9698
3.|9698,9700
Apixaban|9701,9709
5|9710,9711
mg|9712,9714
PO|9715,9717
BID|9718,9721
<EOL>|9722,9723
4.|9723,9725
Aspirin|9726,9733
81|9734,9736
mg|9737,9739
PO|9740,9742
DAILY|9743,9748
<EOL>|9749,9750
5.|9750,9752
Atorvastatin|9753,9765
10|9766,9768
mg|9769,9771
PO|9772,9774
QPM|9775,9778
<EOL>|9779,9780
6.|9780,9782
Diltiazem|9783,9792
Extended|9793,9801
-|9801,9802
Release|9802,9809
240|9810,9813
mg|9814,9816
PO|9817,9819
BID|9820,9823
<EOL>|9824,9825
7.|9825,9827
Docusate|9828,9836
Sodium|9837,9843
100|9844,9847
mg|9848,9850
PO|9851,9853
BID|9854,9857
<EOL>|9858,9859
8.|9859,9861
Dorzolamide|9862,9873
2|9874,9875
%|9875,9876
Ophth|9877,9882
.|9882,9883
Soln.|9884,9889
1|9890,9891
DROP|9892,9896
BOTH|9897,9901
EYES|9902,9906
BID|9907,9910
<EOL>|9911,9912
9.|9912,9914
Ferrous|9915,9922
Sulfate|9923,9930
325|9931,9934
mg|9935,9937
PO|9938,9940
DAILY|9941,9946
<EOL>|9947,9948
10.|9948,9951
Fluticasone|9952,9963
Propionate|9964,9974
NASAL|9975,9980
2|9981,9982
SPRY|9983,9987
NU|9988,9990
DAILY|9991,9996
:|9996,9997
PRN|9997,10000
allergies|10001,10010
<EOL>|10011,10012
11|10012,10014
.|10014,10015
Fluticasone|10016,10027
-|10027,10028
Salmeterol|10028,10038
Diskus|10039,10045
(|10046,10047
500|10047,10050
/|10050,10051
50|10051,10053
)|10053,10054
1|10056,10057
INH|10058,10061
IH|10062,10064
BID|10065,10068
<EOL>|10069,10070
12.|10070,10073
Guaifenesin|10074,10085
_|10086,10087
_|10087,10088
_|10088,10089
mL|10090,10092
PO|10093,10095
Q4H|10096,10099
:|10099,10100
PRN|10100,10103
cough|10104,10109
<EOL>|10110,10111
13.|10111,10114
Hydrochlorothiazide|10115,10134
50|10135,10137
mg|10138,10140
PO|10141,10143
DAILY|10144,10149
<EOL>|10150,10151
14.|10151,10154
Isosorbide|10155,10165
Mononitrate|10166,10177
(|10178,10179
Extended|10179,10187
Release|10188,10195
)|10195,10196
240|10197,10200
mg|10201,10203
PO|10204,10206
DAILY|10207,10212
<EOL>|10213,10214
15.|10214,10217
Latanoprost|10218,10229
0.005|10230,10235
%|10235,10236
Ophth|10237,10242
.|10242,10243
Soln.|10244,10249
1|10250,10251
DROP|10252,10256
BOTH|10257,10261
EYES|10262,10266
QHS|10267,10270
<EOL>|10271,10272
16|10272,10274
.|10274,10275
Lorazepam|10276,10285
0.5|10286,10289
mg|10290,10292
PO|10293,10295
Q8H|10296,10299
:|10299,10300
PRN|10300,10303
Anxiety|10304,10311
<EOL>|10312,10313
17.|10313,10316
Multivitamins|10317,10330
1|10331,10332
TAB|10333,10336
PO|10337,10339
DAILY|10340,10345
<EOL>|10346,10347
18.|10347,10350
Ranitidine|10351,10361
300|10362,10365
mg|10366,10368
PO|10369,10371
DAILY|10372,10377
<EOL>|10378,10379
19|10379,10381
.|10381,10382
Theophylline|10383,10395
SR|10396,10398
300|10399,10402
mg|10403,10405
PO|10406,10408
BID|10409,10412
<EOL>|10413,10414
20|10414,10416
.|10416,10417
Tiotropium|10418,10428
Bromide|10429,10436
1|10437,10438
CAP|10439,10442
IH|10443,10445
DAILY|10446,10451
<EOL>|10452,10453
21|10453,10455
.|10455,10456
Calcitrate|10457,10467
-|10467,10468
Vitamin|10468,10475
D|10476,10477
(|10478,10479
calcium|10479,10486
citrate|10487,10494
-|10494,10495
vitamin|10495,10502
D3|10503,10505
)|10505,10506
315|10507,10510
mg|10511,10513
-|10514,10515
<EOL>|10516,10517
200|10517,10520
units|10521,10526
oral|10528,10532
DAILY|10533,10538
<EOL>|10539,10540
22.|10540,10543
cod|10544,10547
liver|10548,10553
oil|10554,10557
1|10558,10559
capsule|10560,10567
oral|10569,10573
BID|10574,10577
<EOL>|10578,10579
23|10579,10581
.|10581,10582
Ipratropium|10583,10594
Bromide|10595,10602
Neb|10603,10606
1|10607,10608
NEB|10609,10612
IH|10613,10615
Q6H|10616,10619
:|10619,10620
PRN|10620,10623
Wheezing|10624,10632
<EOL>|10633,10634
24|10634,10636
.|10636,10637
Nicotine|10638,10646
Patch|10647,10652
7|10653,10654
mg|10655,10657
TD|10658,10660
DAILY|10661,10666
<EOL>|10667,10668
25|10668,10670
.|10670,10671
Azithromycin|10672,10684
250|10685,10688
mg|10689,10691
PO|10692,10694
Q24H|10695,10699
Duration|10700,10708
:|10708,10709
4|10710,10711
Doses|10712,10717
<EOL>|10718,10719
please|10719,10725
take|10726,10730
until|10731,10736
_|10737,10738
_|10738,10739
_|10739,10740
.|10740,10741
PredniSONE|10742,10752
40|10753,10755
mg|10756,10758
PO|10759,10761
DAILY|10762,10767
Duration|10768,10776
:|10776,10777
5|10778,10779
Days|10780,10784
<EOL>|10785,10786
40mg|10786,10790
until|10791,10796
_|10797,10798
_|10798,10799
_|10799,10800
<EOL>|10801,10802
Tapered|10802,10809
dose|10810,10814
-|10815,10816
DOWN|10817,10821
<EOL>|10822,10823
<EOL>|10823,10824
<EOL>|10825,10826
Discharge|10826,10835
Disposition|10836,10847
:|10847,10848
<EOL>|10848,10849
Extended|10849,10857
Care|10858,10862
<EOL>|10862,10863
<EOL>|10864,10865
Facility|10865,10873
:|10873,10874
<EOL>|10874,10875
_|10875,10876
_|10876,10877
_|10877,10878
<EOL>|10878,10879
<EOL>|10880,10881
_|10881,10882
_|10882,10883
_|10883,10884
Diagnosis|10885,10894
:|10894,10895
<EOL>|10895,10896
PRIMARY|10896,10903
:|10903,10904
<EOL>|10904,10905
COPD|10905,10909
Exacerbation|10910,10922
<EOL>|10922,10923
<EOL>|10923,10924
SECONDARY|10924,10933
:|10933,10934
<EOL>|10934,10935
Afib|10935,10939
<EOL>|10939,10940
Anxiety|10940,10947
<EOL>|10947,10948
HTN|10948,10951
<EOL>|10951,10952
CAD|10952,10955
<EOL>|10955,10956
<EOL>|10956,10957
<EOL>|10958,10959
Discharge|10959,10968
Condition|10969,10978
:|10978,10979
<EOL>|10979,10980
Mental|10980,10986
Status|10987,10993
:|10993,10994
Clear|10995,11000
and|11001,11004
coherent|11005,11013
.|11013,11014
<EOL>|11014,11015
Level|11015,11020
of|11021,11023
Consciousness|11024,11037
:|11037,11038
Alert|11039,11044
and|11045,11048
interactive|11049,11060
.|11060,11061
<EOL>|11061,11062
Activity|11062,11070
Status|11071,11077
:|11077,11078
Ambulatory|11079,11089
-|11090,11091
requires|11092,11100
assistance|11101,11111
or|11112,11114
aid|11115,11118
(|11119,11120
walker|11120,11126
<EOL>|11127,11128
or|11128,11130
cane|11131,11135
)|11135,11136
.|11136,11137
<EOL>|11137,11138
<EOL>|11138,11139
<EOL>|11140,11141
Discharge|11141,11150
Instructions|11151,11163
:|11163,11164
<EOL>|11164,11165
Dear|11165,11169
Ms.|11170,11173
_|11174,11175
_|11175,11176
_|11176,11177
,|11177,11178
<EOL>|11178,11179
<EOL>|11179,11180
You|11180,11183
were|11184,11188
admitted|11189,11197
to|11198,11200
_|11201,11202
_|11202,11203
_|11203,11204
after|11205,11210
you|11211,11214
developed|11215,11224
<EOL>|11225,11226
shortness|11226,11235
of|11236,11238
breath|11239,11245
and|11246,11249
wheezing|11250,11258
at|11259,11261
home|11262,11266
shortly|11267,11274
after|11275,11280
your|11281,11285
last|11286,11290
<EOL>|11291,11292
discharge|11292,11301
.|11301,11302
You|11303,11306
were|11307,11311
treated|11312,11319
for|11320,11323
a|11324,11325
COPD|11326,11330
exacerbation|11331,11343
and|11344,11347
your|11348,11352
<EOL>|11353,11354
breathing|11354,11363
quickly|11364,11371
got|11372,11375
better|11376,11382
.|11382,11383
Our|11384,11387
physical|11388,11396
therapists|11397,11407
evaluated|11408,11417
<EOL>|11418,11419
you|11419,11422
and|11423,11426
recommended|11427,11438
that|11439,11443
you|11444,11447
have|11448,11452
a|11453,11454
short|11455,11460
stay|11461,11465
at|11466,11468
Pulmonary|11469,11478
<EOL>|11479,11480
_|11480,11481
_|11481,11482
_|11482,11483
before|11484,11490
going|11491,11496
home|11497,11501
to|11502,11504
improve|11505,11512
your|11513,11517
breathing|11518,11527
.|11527,11528
<EOL>|11529,11530
<EOL>|11530,11531
We|11531,11533
wish|11534,11538
you|11539,11542
all|11543,11546
the|11547,11550
best|11551,11555
at|11556,11558
rehab|11559,11564
and|11565,11568
send|11569,11573
our|11574,11577
condolences|11578,11589
to|11590,11592
<EOL>|11593,11594
your|11594,11598
family|11599,11605
on|11606,11608
your|11609,11613
recent|11614,11620
loss|11621,11625
.|11625,11626
<EOL>|11626,11627
<EOL>|11627,11628
It|11628,11630
was|11631,11634
truly|11635,11640
a|11641,11642
pleasure|11643,11651
taking|11652,11658
care|11659,11663
of|11664,11666
you|11667,11670
.|11670,11671
<EOL>|11671,11672
<EOL>|11672,11673
Your|11673,11677
_|11678,11679
_|11679,11680
_|11680,11681
Team|11682,11686
<EOL>|11686,11687
<EOL>|11688,11689
Followup|11689,11697
Instructions|11698,11710
:|11710,11711
<EOL>|11711,11712
_|11712,11713
_|11713,11714
_|11714,11715
<EOL>|11715,11716

