CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Hallucinations, Visual|Finding|false|false||Visual hallucinationsnull|Visual|Finding|false|false||Visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Disease|Disorder|false|false||diseasenull|Dyslipidemias|Disorder|false|false||dyslipidemianull|Medical History|Finding|false|false|C0033572;C4266527|history ofnull|History of present illness (finding)|Finding|false|false|C0033572;C4266527|history
null|History of previous events|Finding|false|false|C0033572;C4266527|history
null|Historical aspects qualifier|Finding|false|false|C0033572;C4266527|history
null|Medical History|Finding|false|false|C0033572;C4266527|history
null|Concept History|Finding|false|false|C0033572;C4266527|historynull|History|Subject|false|false||historynull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0262926;C0376358;C0600139;C0006826;C0262926;C1705255;C0019665;C0262512;C2004062;C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0262926;C0376358;C0600139;C0006826;C0262926;C1705255;C0019665;C0262512;C2004062;C0496923;C0154088;C0033575;C0154009|prostatenull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Prostatectomy|Procedure|false|false||prostatectomynull|Neurologists|Subject|false|false||neurologistnull|Gait|Finding|false|false||gaitnull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Chart evaluation by healthcare professional|Procedure|false|false||chart reviewnull|Charts (publication)|Finding|false|false||chartnull|chart [medical device]|Device|false|false||chartnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Neurologists|Subject|false|false||neurologistnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Gait|Finding|false|false||gaitnull|Frozen behavior|Finding|false|false||freezingnull|Freezing|Phenomenon|false|false||freezingnull|Gait|Finding|false|false||gaitnull|Frozen behavior|Finding|false|false||freezingnull|Freezing|Phenomenon|false|false||freezingnull|Mirapex|Drug|false|false||mirapex
null|Mirapex|Drug|false|false||mirapexnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Neurologists|Subject|false|false||neurologistnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Mirapex|Drug|false|false||Mirapex
null|Mirapex|Drug|false|false||Mirapexnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Daughter|Subject|false|false||daughternull|Progressive|Finding|false|false||progressivenull|Gait|Finding|false|false||gaitnull|Stiffness|Finding|false|false||stiffnessnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Difficult (qualifier value)|Finding|false|false||difficulty withnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Bathroom|Device|false|false||bathroom
null|Toilet Facilities|Device|false|false||bathroomnull|Episode of|Time|false|false||episodesnull|Incontinence|Disorder|false|false||incontinencenull|Reassuring (procedure)|Procedure|false|false||reassuringnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Presentation|Finding|false|false||presentationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Experience (Practice)|Finding|false|false||experience
null|Experience|Finding|false|false||experiencenull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Cross syndrome|Disorder|false|false||crossnull|Traverse|Finding|false|false||crossnull|AMACR wt Allele|Finding|false|false||race
null|AMACR gene|Finding|false|false||racenull|Rapid Amplification of cDNA Ends|Procedure|false|false||racenull|null|Attribute|false|false||racenull|Race (classification)|Subject|false|false||race
null|Race|Subject|false|false||racenull|History of fall|Finding|false|false||a fallnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|wife|Subject|false|false||wifenull|Unable|Finding|false|false|C3714591|unablenull|Floor (anatomic)|Anatomy|false|false|C1299582|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076|head
null|Head|Anatomy|false|false|C0876917;C0362076|headnull|Head Device|Device|false|false||headnull|Strikes, Employee|Event|true|false||strikenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|wife|Subject|false|false||wifenull|Gait|Finding|false|false||gaitnull|Hour|Time|false|false||hoursnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Unable|Finding|false|false||unablenull|Ambulate|Finding|false|false||ambulatenull|Own|Finding|false|false||ownnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Daughter|Subject|false|false||daughternull|Neurologists|Subject|false|false||neurologistnull|Presentation|Finding|false|false||presentationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|HGS protein, human|Drug|false|false||HRs
null|HGS protein, human|Drug|false|false||HRsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||HRsnull|HARS1 wt Allele|Finding|false|false||HRs
null|HARS1 gene|Finding|false|false||HRs
null|HGS wt Allele|Finding|false|false||HRs
null|HGS gene|Finding|false|false||HRs
null|ATN1 wt Allele|Finding|false|false||HRs
null|SRSF5 gene|Finding|false|false||HRsnull|Hour|Time|false|false||HRsnull|Saturation of Peripheral Oxygen|Attribute|false|false||SpO2null|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Cogwheel Rigidity|Finding|false|false||cogwheelingnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|All extremities|Anatomy|false|false|C0392756;C0808080|extremities
null|Limb structure|Anatomy|false|false|C0392756;C0808080|extremitiesnull|Reduced|Finding|false|false|C0278454;C0015385|decreasenull|Decrease|LabModifier|false|false||decreasenull|Strength (attribute)|Finding|false|false|C0278454;C0015385|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Laboratory test finding|Lab|false|false||Labsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|TOX protein, human|Drug|false|false||tox
null|TOX protein, human|Drug|false|false||toxnull|TOX gene|Finding|false|false||toxnull|Toxicity aspects|Modifier|false|false||toxnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|null|Modifier|false|false||unremarkablenull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C0009555|CBCnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0741025|Chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|Chestnull|Diagnostic radiologic examination|Procedure|false|false||Xraynull|Roentgen Rays|Phenomenon|false|false||Xraynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Process Pharmacologic Substance|Drug|false|false|C1184743|processnull|Process (qualifier value)|Finding|false|false|C1184743|processnull|bony process|Anatomy|false|false|C1538070;C1413792;C4521054;C1951340;C1522240|processnull|Process|Phenomenon|false|false|C1184743|processnull|CTH protein, human|Drug|false|false||CTH
null|CTH protein, human|Drug|false|false||CTHnull|CTH gene|Finding|false|false|C1184743|CTH
null|VSIG2 gene|Finding|false|false|C1184743|CTHnull|Reassuring (procedure)|Procedure|false|false||reassuringnull|Neurology speciality|Title|false|false||neurologynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Patient's home|Device|false|false||patient's homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Metabolic Process, Cellular|Finding|false|false||metabolic
null|Metabolic|Finding|false|false||metabolicnull|Multisection metabolic|Procedure|false|false||metabolicnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|pramipexole|Drug|false|false||pramipexole
null|pramipexole|Drug|false|false||pramipexolenull|pravastatin|Drug|false|false||pravastatin
null|pravastatin|Drug|false|false||pravastatinnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feeling comfortable|Finding|false|false||comfortablenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Published Interview|Finding|false|false||interviewnull|Interview|Event|false|false||interviewnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|SURE Test|Finding|true|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Party|Finding|false|false||partynull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Cross syndrome|Disorder|false|false||crossnull|Traverse|Finding|false|false||crossnull|AMACR wt Allele|Finding|false|false||race
null|AMACR gene|Finding|false|false||racenull|Rapid Amplification of cDNA Ends|Procedure|false|false||racenull|null|Attribute|false|false||racenull|Race (classification)|Subject|false|false||race
null|Race|Subject|false|false||racenull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|History of fall|Finding|false|false||a fallnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|year|Time|false|false||yearsnull|Fever|Finding|false|false||feversnull|Chills|Finding|false|false||chillsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C1549543;C0030193;C0008031;C0741025;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C1549543;C0030193;C0008031;C0741025;C2926613|chestnull|Abdominal Pain|Finding|false|false|C0000726|pain, abdominalnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Dysuria|Finding|false|false||dysurianull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Disease|Disorder|false|false||diseasenull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C1551342;C0497327;C0011265|Body
null|Human body structure|Anatomy|false|false|C1551342;C0497327;C0011265|Body
null|Body structure|Anatomy|false|false|C1551342;C0497327;C0011265|Body
null|Adult human body|Anatomy|false|false|C1551342;C0497327;C0011265|Body
null|Whole body|Anatomy|false|false|C1551342;C0497327;C0011265|Bodynull|Human body|Subject|false|false||Bodynull|Presenile dementia|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Dementia
null|Dementia|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Dementianull|Dyslipidemias|Disorder|false|false||dyslipidemianull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0376358;C0600139;C0496923;C0154088;C0033575;C0154009;C0006826|prostate
null|Prostate|Anatomy|false|false|C0376358;C0600139;C0496923;C0154088;C0033575;C0154009;C0006826|prostatenull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Prostatectomy|Procedure|false|false||prostatectomynull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Senility|Finding|false|false||old agenull|Old age|Time|false|false||old agenull|Old|Time|false|false||oldnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0006826;C0496923;C0154088;C0033575;C0154009;C0376358;C0600139|prostate
null|Prostate|Anatomy|false|false|C0006826;C0496923;C0154088;C0033575;C0154009;C0376358;C0600139|prostatenull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Sister - courtesy title|Finding|false|false||sister
null|Relationship - Sister|Finding|false|false||sisternull|Sister|Subject|false|false||sisternull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Younger sister|Subject|false|false||younger sisternull|Sister - courtesy title|Finding|false|false||sister
null|Relationship - Sister|Finding|false|false||sisternull|Sister|Subject|false|false||sisternull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Brother - courtesy title|Finding|false|false||brother
null|Relationship - Brother|Finding|false|false||brothernull|Brothers|Subject|false|false||brothernull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Daughter|Subject|false|false||daughtersnull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Neurologic (qualifier value)|Modifier|false|false||neurologicnull|Illness (finding)|Finding|false|false||illnessnull|Presenile dementia|Disorder|false|false||dementia
null|Dementia|Disorder|false|false||dementianull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Mental disorders|Disorder|false|false||mental disordersnull|Psyche structure|Finding|false|false||mentalnull|Disease|Disorder|false|false||disordersnull|Learning|Finding|false|false||learningnull|Knowledge acquisition|Procedure|false|false||learningnull|Disability|Finding|false|false||disabilitynull|null|Attribute|false|false||disabilitynull|Attention deficit hyperactivity disorder|Disorder|false|false||ADHDnull|Family Medical History|Finding|true|false||family history ofnull|Family Medical History|Finding|true|false||family historynull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|true|true||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Referral type - Psychiatric|Finding|true|true||psychiatric
null|Psychiatric|Finding|true|true||psychiatricnull|Psychiatric service|Procedure|true|true||psychiatricnull|Psychiatry Specialty|Title|false|false||psychiatricnull|Problems - What subject filter|Finding|false|false||problemsnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|ATP5F1A gene|Finding|false|false||OMRnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|patient appears in no acute distress (physical finding)|Finding|false|false||In no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C1828121;C0021485;C1533685;C2228481;C0036412;C0205180|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Injection|Drug|true|false||injectionnull|Injection Route of Administration|Finding|true|false|C0036410|injectionnull|Injection of therapeutic agent|Procedure|true|false|C0036410|injection
null|Injection procedure|Procedure|true|false|C0036410|injectionnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Cervical lymphadenopathy|Disorder|true|false|C0027530|cervical lymphadenopathynull|Swollen lymph nodes in the neck|Finding|true|false|C0027530|cervical lymphadenopathynull|Neck|Anatomy|false|false|C4551446;C0497156;C0235592;C4282165|cervicalnull|Cervical|Modifier|false|false||cervicalnull|Lymphadenopathy|Disorder|true|false|C0027530|lymphadenopathynull|Swollen Lymph Node|Finding|true|false|C0027530|lymphadenopathynull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Regular|Modifier|false|false||Regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Heart murmur|Finding|false|false||murmursnull|Pericardial friction rub|Finding|false|false||rubsnull|Lung|Anatomy|false|false||LUNGSnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Increased work of breathing|Finding|true|false||increased work of breathingnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|false|false||increasednull|Work of Breathing|Finding|true|false||work of breathingnull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Renal angle tenderness|Finding|true|false||CVA tendernessnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0153662;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|ABDOMENnull|Intestines|Anatomy|false|false||bowelsnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Palpation|Procedure|false|false||palpationnull|Four quadrants|Modifier|false|false||four quadrantsnull|Organomegaly|Finding|true|false||organomegalynull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|null|Drug|false|false||Pulsesnull|Physiologic pulse|Finding|false|false||Pulsesnull|Pulse taking|Procedure|false|false||Pulsesnull|Radial|Finding|false|false||Radial
null|Circumpennate|Finding|false|false||Radialnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|refill|Finding|false|false||refillnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Neurologic (qualifier value)|Modifier|false|false||NEUROLOGICnull|CNDP2 gene|Finding|false|false||CN2null|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Muscle Hypertonia|Finding|false|false||Increased tonenull|Lewis Blood-Group System|Finding|false|false|C0227192|LEsnull|Inferior esophageal sphincter structure|Anatomy|false|false|C0023595|LEsnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|Last|Modifier|false|false||lastnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|patient appears in no acute distress (physical finding)|Finding|false|false||In no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Very|Modifier|false|false||verynull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Regular|Modifier|false|false||Regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Heart murmur|Finding|false|false||murmursnull|Pericardial friction rub|Finding|false|false||rubsnull|Lung|Anatomy|false|false||LUNGSnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Increased work of breathing|Finding|true|false||increased work of breathingnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|false|false||increasednull|Work of Breathing|Finding|true|false||work of breathingnull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Intestines|Anatomy|false|false||bowelsnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Palpation|Procedure|false|false||palpationnull|Four quadrants|Modifier|false|false||four quadrantsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|null|Drug|false|false||Pulsesnull|Physiologic pulse|Finding|false|false||Pulsesnull|Pulse taking|Procedure|false|false||Pulsesnull|Radial|Finding|false|false||Radial
null|Circumpennate|Finding|false|false||Radialnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Neurologic (qualifier value)|Modifier|false|false||NEUROLOGICnull|CNDP2 gene|Finding|false|false||CN2null|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Muscle Hypertonia|Finding|false|false||Increased tonenull|Lewis Blood-Group System|Finding|false|false|C0227192|LEsnull|Inferior esophageal sphincter structure|Anatomy|false|false|C0023595|LEsnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1266129;C1370889;C2257651;C1415274;C1140170;C4553172;C0004002;C0242192;C1121182;C4522245;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|AB(S) hearing assessment list|Device|false|false||Abnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||Ethanol
null|CNS depressants ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanolnull|Toxic effect of ethyl alcohol|Disorder|false|false||Ethanolnull|Ethanol measurement|Procedure|false|false||Ethanolnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Imaging problem|Finding|false|false|C0018670;C0152336|Imagingnull|Diagnostic Imaging|Procedure|false|false|C0018670;C0152336|Imaging
null|Imaging Techniques|Procedure|false|false|C0018670;C0152336|Imagingnull|Imaging Technology|Title|false|false||Imagingnull|CAT scan of head|Procedure|false|false|C0018670;C0152336|CT HEADnull|null|Attribute|false|false|C0018670;C0152336|CT HEADnull|Problems with head|Disorder|false|false|C0018670;C0152336|HEADnull|Procedure on head|Procedure|false|false|C0018670;C0152336|HEADnull|Structure of head of caudate nucleus|Anatomy|false|false|C0740845;C0881943;C0202691;C0079595;C0011923;C0362076;C0876917|HEAD
null|Head|Anatomy|false|false|C0740845;C0881943;C0202691;C0079595;C0011923;C0362076;C0876917|HEADnull|Head Device|Device|false|false||HEADnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Infarction|Finding|true|false||infarctionnull|Hemorrhage|Finding|true|false||hemorrhagenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Mass of body structure|Finding|true|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false||mass
null|null|Finding|true|false||mass
null|FBN1 wt Allele|Finding|true|false||mass
null|FBN1 gene|Finding|true|false||mass
null|Mass of body region|Finding|true|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Heart Ventricle|Anatomy|false|false||ventriclesnull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Fracture|Disorder|true|false||fracturenull|Part|Modifier|false|false||portionnull|Nasal sinus|Anatomy|false|false|C2228461;C1550016;C0016169;C0496788;C0271428;C0851354;C1510420;C0011334;C1546608;C1550629;C1552826|paranasal sinusesnull|pathologic fistula|Disorder|false|false|C0030471;C4071871;C0030471;C0013455|sinusesnull|Head>Sinuses|Anatomy|false|false|C0851354;C0016169;C0496788;C0271428;C1552826;C2228461;C1510420;C0011334;C1550016;C1546608;C1550629|sinuses
null|Nasal sinus|Anatomy|false|false|C0851354;C0016169;C0496788;C0271428;C1552826;C2228461;C1510420;C0011334;C1550016;C1546608;C1550629|sinusesnull|Malignant neoplasm of middle ear|Disorder|false|false|C4071871;C0030471;C0030471;C0333343;C0013455;C0013443;C0521421|middle ear
null|Disorder of middle ear|Disorder|false|false|C4071871;C0030471;C0030471;C0333343;C0013455;C0013443;C0521421|middle earnull|examination of middle ear|Procedure|false|false|C0030471;C0333343;C0013443;C0521421;C0013455;C4071871;C0030471|middle earnull|middle ear|Anatomy|false|false|C1550016;C0851354;C0016169;C2228461;C1552826;C0496788;C0271428;C1510420;C0011334|middle earnull|Table Cell Vertical Align - middle|Finding|false|false|C0013455;C4071871;C0030471;C0030471|middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Ear and labyrinth disorders|Disorder|false|false|C4071871;C0030471;C0013455;C0013443;C0521421;C0030471;C0333343|earnull|SpecimenType - Ear|Finding|false|false|C0333343;C0013443;C0521421;C0030471;C4071871;C0030471|ear
null|null|Finding|false|false|C0333343;C0013443;C0521421;C0030471;C4071871;C0030471|earnull|Ear structure|Anatomy|false|false|C2228461;C0851354;C1546608;C1550629;C0496788;C0271428|ear
null|null|Anatomy|false|false|C2228461;C0851354;C1546608;C1550629;C0496788;C0271428|earnull|Dental caries|Disorder|false|false|C0030471;C0333343;C4071871;C0030471;C0013455|cavities
null|Cavitation|Disorder|false|false|C0030471;C0333343;C4071871;C0030471;C0013455|cavitiesnull|Body cavities|Anatomy|false|false|C1550016;C1546608;C1550629;C2228461;C0496788;C0271428;C1510420;C0011334;C0851354|cavitiesnull|Remote control command - Clear|Finding|false|false|C0333343;C0030471;C0013455;C4071871;C0030471|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Part|Modifier|false|false||portionnull|Ocular orbit|Anatomy|false|false||orbitsnull|null|Modifier|false|false||unremarkablenull|Bilateral|Modifier|false|false||bilateralnull|Lens Diseases|Disorder|false|false|C0023317|lensnull|examination of lens|Procedure|false|false|C0023317|lensnull|Lens, Crystalline|Anatomy|false|false|C0035139;C2239142;C0023308|lensnull|Lens Device|Device|false|false||lensnull|Lens <eudicots>|Entity|false|false||lens
null|Lens <bivalves>|Entity|false|false||lensnull|Surgical Replantation|Procedure|false|false|C0023317|replacementsnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false|C0524466|intracranialnull|Intracranial|Anatomy|false|false|C0000768;C1522213|intracranialnull|Congenital Abnormality|Disorder|true|false|C0524466|abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Hydrocephalus|Disorder|true|false||hydrocephalusnull|Imaging problem|Finding|false|false|C1527391;C0817096|Imagingnull|Diagnostic Imaging|Procedure|false|false|C1527391;C0817096|Imaging
null|Imaging Techniques|Procedure|false|false|C1527391;C0817096|Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Chest problem|Finding|false|false|C1527391;C0817096|CHESTnull|Chest|Anatomy|false|false|C0740845;C0079595;C0011923;C0741025|CHEST
null|Anterior thoracic region|Anatomy|false|false|C0740845;C0079595;C0011923;C0741025|CHESTnull|LAT protein, human|Drug|false|false||LAT
null|L-Type Amino Acid Transporter|Drug|false|false||LAT
null|L-Type Amino Acid Transporter|Drug|false|false||LAT
null|ORC3 protein, human|Drug|false|false||LAT
null|ORC3 protein, human|Drug|false|false||LAT
null|LAT protein, human|Drug|false|false||LATnull|LAT gene|Finding|false|false||LAT
null|ORC3 wt Allele|Finding|false|false||LAT
null|ORC3 gene|Finding|false|false||LAT
null|SPNS1 gene|Finding|false|false||LATnull|Latin Language|Entity|false|false||LATnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Atelectasis|Finding|false|false||atelectasisnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C0740941;C0024115|lungnull|Base|Drug|false|false||basesnull|Base - unit of product usage|LabModifier|false|false||basesnull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|true|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Glycation End Products, Advanced|Drug|false|false||Age
null|Glycation End Products, Advanced|Drug|false|false||Agenull|null|Attribute|false|false||Agenull|Age|Subject|false|false||Agenull|Indeterminate|Modifier|false|false||indeterminatenull|Moderate to severe|Modifier|false|false||moderate to severenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Deformity|Disorder|false|false||deformity
null|Congenital Abnormality|Disorder|false|false||deformitynull|null|Finding|false|false||deformitynull|IPSS-R Risk Category Low|Finding|false|false|C0223084;C0817096;C1305451;C0223199|low
null|IPSS Risk Category Low|Finding|false|false|C0223084;C0817096;C1305451;C0223199|low
null|low confidentiality|Finding|false|false|C0223084;C0817096;C1305451;C0223199|lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|null|Anatomy|false|false|C5779551;C5203106;C4522223;C1550472;C1551342|thoracic vertebral body
null|Structure of body of thoracic vertebra|Anatomy|false|false|C5779551;C5203106;C4522223;C1550472;C1551342|thoracic vertebral bodynull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false|C1305451;C0223199;C0223084;C0817096|thoracicnull|Chest|Anatomy|false|false|C5203106;C4522223;C1550472;C1551342;C5779551|thoracicnull|Body of vertebra|Anatomy|false|false|C5203106;C4522223;C1550472;C1551342;C5779551|vertebral bodynull|Bone structure of spine|Anatomy|false|false|C1551342|vertebralnull|Document Body|Finding|false|false|C0223084;C0817096;C0549207;C1305451;C0223199;C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C1551342|body
null|Human body structure|Anatomy|false|false|C1551342|body
null|Body structure|Anatomy|false|false|C1551342|body
null|Adult human body|Anatomy|false|false|C1551342|body
null|Whole body|Anatomy|false|false|C1551342|bodynull|Human body|Subject|false|false||bodynull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Disease|Disorder|false|false||diseasenull|Dyslipidemias|Disorder|false|false||dyslipidemianull|Medical History|Finding|false|false|C0033572;C4266527|history ofnull|History of present illness (finding)|Finding|false|false|C0033572;C4266527|history
null|History of previous events|Finding|false|false|C0033572;C4266527|history
null|Historical aspects qualifier|Finding|false|false|C0033572;C4266527|history
null|Medical History|Finding|false|false|C0033572;C4266527|history
null|Concept History|Finding|false|false|C0033572;C4266527|historynull|History|Subject|false|false||historynull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0262926;C0006826;C0262926;C1705255;C0019665;C0262512;C2004062;C0376358;C0600139;C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0262926;C0006826;C0262926;C1705255;C0019665;C0262512;C2004062;C0376358;C0600139;C0496923;C0154088;C0033575;C0154009|prostatenull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Prostatectomy|Procedure|false|false||prostatectomynull|Neurologists|Subject|false|false||neurologistnull|Gait|Finding|false|false||gaitnull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|nervous system disorder|Disorder|false|false||neurologic disordernull|Neurologic (qualifier value)|Modifier|false|false||neurologicnull|Disease|Disorder|false|false||disordernull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Disease|Disorder|false|false||diseasenull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C0497327;C0011265;C1551342|Body
null|Human body structure|Anatomy|false|false|C0497327;C0011265;C1551342|Body
null|Body structure|Anatomy|false|false|C0497327;C0011265;C1551342|Body
null|Adult human body|Anatomy|false|false|C0497327;C0011265;C1551342|Body
null|Whole body|Anatomy|false|false|C0497327;C0011265;C1551342|Bodynull|Human body|Subject|false|false||Bodynull|Presenile dementia|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Dementia
null|Dementia|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|Dementianull|Hallucinations, Visual|Finding|false|false||Visual Hallucinationsnull|Visual|Finding|false|false||Visualnull|Hallucinations|Disorder|false|false||Hallucinationsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Acute-on-chronic|Time|false|false||acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|false|false||disease progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Mirapex|Drug|false|false||mirapex
null|Mirapex|Drug|false|false||mirapexnull|rasagiline|Drug|false|false||rasagiline
null|rasagiline|Drug|false|false||rasagilinenull|rivastigmine|Drug|false|false||rivastigmine
null|rivastigmine|Drug|false|false||rivastigminenull|Neurology speciality|Title|false|false||Neurologynull|Seroquel|Drug|false|false||Seroquel
null|Seroquel|Drug|false|false||Seroquelnull|Hallucinations|Disorder|false|false||hallucinationsnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Rehabilitation therapy|Procedure|false|false||rehabnull|Recommendation|Finding|false|false||recommendationnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Discharge to home|Procedure|false|false||discharge to homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Goals of Care|Procedure|false|false||goals of carenull|What subject filter - Goals|Finding|false|false||goals
null|objective (goal)|Finding|false|false||goals
null|treatment goals|Finding|false|false||goalsnull|null|Attribute|false|false||goalsnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Hallucinations, Visual|Finding|false|false||visual hallucinationnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Seroquel|Drug|false|false||Seroquel
null|Seroquel|Drug|false|false||Seroquelnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|rasagiline|Drug|false|false||Rasagiline
null|rasagiline|Drug|false|false||Rasagilinenull|Daily|Time|false|false||DAILYnull|pramipexole|Drug|false|false||Pramipexole
null|pramipexole|Drug|false|false||Pramipexolenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|rivastigmine|Drug|false|false||rivastigmine
null|rivastigmine|Drug|false|false||rivastigminenull|Transdermal Route of Administration|Finding|false|false||transdermal
null|transdermal|Finding|false|false||transdermal
null|Transdermal (intended site)|Finding|false|false||transdermalnull|Daily|Time|false|false||DAILYnull|pravastatin|Drug|false|false||Pravastatin
null|pravastatin|Drug|false|false||Pravastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalaminnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|unknown vaccine or immune globulin|Drug|false|false||Unknown
null|Unknown - Vaccines administered|Drug|false|false||Unknown
null|Unknown - Vaccines administered|Drug|false|false||Unknown
null|unknown vaccine or immune globulin|Drug|false|false||Unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||Unknown
null|Unknown - Special Program Code|Finding|false|false||Unknown
null|Unknown - Production Class Code|Finding|false|false||Unknown
null|Unknown - Patient Outcome|Finding|false|false||Unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||Unknown
null|Unknown - Escort Required|Finding|false|false||Unknown
null|Unknown - Transport Arranged|Finding|false|false||Unknown
null|Unknown - Living Arrangement|Finding|false|false||Unknown
null|Unknown - Employment Status|Finding|false|false||Unknown
null|Unknown - Relationship|Finding|false|false||Unknown
null|Unknown - publishing section|Finding|false|false||Unknown
null|Unknown Publicity Code|Finding|false|false||Unknown
null|Unknown - Event reason|Finding|false|false||Unknown
null|Unknown - Religion|Finding|false|false||Unknown
null|Unknown - Organ Donor Code|Finding|false|false||Unknown
null|unknown - NullFlavor|Finding|false|false||Unknown
null|Unknown - Notify Clergy Code|Finding|false|false||Unknown
null|Unknown - Administrative Gender|Finding|false|false||Unknown
null|Unknown - Patient Condition Code|Finding|false|false||Unknown
null|Unknown - Living Will Code|Finding|false|false||Unknown
null|Marital Status - Unknown|Finding|false|false||Unknown
null|Unknown - mode of arrival code|Finding|false|false||Unknown
null|Unknown - Patient Class|Finding|false|false||Unknown
null|Unknown - Event Expected|Finding|false|false||Unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||Unknown
null|Unknown - Immunization Registry Status|Finding|false|false||Unknown
null|Unknown - Container status|Finding|false|false||Unknown
null|Unknown - CWE statuses|Finding|false|false||Unknown
null|Unknown - Job Status|Finding|false|false||Unknown
null|Unknown - Precaution Code|Finding|false|false||Unknown
null|Unknown - Contact Role|Finding|false|false||Unknown
null|Unknown - Living Dependency|Finding|false|false||Unknownnull|Ethnic group unknown|Subject|false|false||Unknownnull|Unknown - Allergy Severity|Modifier|false|false||Unknown
null|Unknown - HL7 update mode|Modifier|false|false||Unknown
null|Unknown|Modifier|false|false||Unknownnull|Daily|Time|false|false||DAILYnull|loratadine|Drug|false|false||Loratadine
null|loratadine|Drug|false|false||Loratadinenull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|quetiapine fumarate|Drug|false|false||QUEtiapine Fumarate
null|quetiapine fumarate|Drug|false|false||QUEtiapine Fumaratenull|quetiapine|Drug|false|false||QUEtiapine
null|quetiapine|Drug|false|false||QUEtiapinenull|fumarate|Drug|false|false||Fumarate
null|fumarate|Drug|false|false||Fumaratenull|Once a day, at bedtime|Time|false|false||QHSnull|quetiapine|Drug|false|false||quetiapine
null|quetiapine|Drug|false|false||quetiapinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Night time|Time|false|false||AT NIGHTnull|Night time|Time|false|false||NIGHTnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|loratadine|Drug|false|false||Loratadine
null|loratadine|Drug|false|false||Loratadinenull|Daily|Time|false|false||DAILYnull|pramipexole|Drug|false|false||Pramipexole
null|pramipexole|Drug|false|false||Pramipexolenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|pravastatin|Drug|false|false||Pravastatin
null|pravastatin|Drug|false|false||Pravastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|rasagiline|Drug|false|false||Rasagiline
null|rasagiline|Drug|false|false||Rasagilinenull|Daily|Time|false|false||DAILYnull|rivastigmine|Drug|false|false||rivastigmine
null|rivastigmine|Drug|false|false||rivastigminenull|Transdermal Route of Administration|Finding|false|false||transdermal
null|transdermal|Finding|false|false||transdermal
null|Transdermal (intended site)|Finding|false|false||transdermalnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Confusion|Disorder|false|false||Confusednull|Precaution Code - Confused|Finding|false|false||Confused
null|Clouded consciousness|Finding|false|false||Confusednull|Sometimes|Time|false|false||sometimesnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Role Privilege|Finding|false|false||privilege
null|User Privilege|Finding|false|false||privilege
null|Privilege|Finding|false|false||privilegenull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Encounter Referral Source - emergency room|Finding|false|false||emergency roomnull|Accident and Emergency department|Device|false|false||emergency roomnull|Accident and Emergency department|Entity|false|false||emergency roomnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Neurologists|Subject|false|false||neurologistnull|Hallucinations, Visual|Finding|false|false||visual hallucinationsnull|Visual|Finding|false|false||visualnull|Hallucinations|Disorder|false|false||hallucinationsnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Continuous|Finding|false|false||Continuenull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Appointments|Event|false|false||appointmentsnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions