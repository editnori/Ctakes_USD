 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Nonexertional|293,306
Chest|307,312
pain|313,317
<EOL>|317,318
<EOL>|319,320
Major|320,325
Surgical|326,334
or|335,337
Invasive|338,346
Procedure|347,356
:|356,357
<EOL>|357,358
none|358,362
<EOL>|362,363
<EOL>|363,364
<EOL>|365,366
This|394,398
is|399,401
a|402,403
_|404,405
_|405,406
_|406,407
year|408,412
old|413,416
female|417,423
with|424,428
PMHx|429,433
CAD|434,437
,|437,438
PVD|439,442
and|443,446
COPD|447,451
<EOL>|452,453
presenting|453,463
with|464,468
chest|469,474
pain|475,479
.|479,480
She|481,484
reports|485,492
that|493,497
she|498,501
woke|502,506
up|507,509
at|510,512
3|513,514
am|515,517
<EOL>|518,519
with|519,523
substernal|524,534
pressure|535,543
like|544,548
pain|549,553
which|554,559
was|560,563
associated|564,574
with|575,579
<EOL>|580,581
shortness|581,590
of|591,593
breath|594,600
.|600,601
She|602,605
rated|606,611
the|612,615
pain|616,620
a|621,622
_|623,624
_|624,625
_|625,626
and|627,630
reports|631,638
that|639,643
<EOL>|644,645
it|645,647
lasted|648,654
for|655,658
about|659,664
5|665,666
minutes|667,674
and|675,678
resolved|679,687
spontaneously|688,701
.|701,702
She|703,706
<EOL>|707,708
had|708,711
several|712,719
more|720,724
episodes|725,733
of|734,736
the|737,740
same|741,745
pain|746,750
lasting|751,758
about|759,764
5|765,766
<EOL>|767,768
minutes|768,775
at|776,778
a|779,780
time|781,785
throughout|786,796
the|797,800
morning|801,808
but|809,812
which|813,818
were|819,823
much|824,828
<EOL>|829,830
less|830,834
severe|835,841
.|841,842
She|843,846
has|847,850
n't|850,853
had|854,857
an|858,860
episode|861,868
of|869,871
pain|872,876
since|877,882
1|883,884
pm|885,887
.|887,888
She|889,892
<EOL>|893,894
denies|894,900
palpitations|901,913
,|913,914
lightheadedness|915,930
,|930,931
dizziness|932,941
,|941,942
nausea|943,949
,|949,950
<EOL>|951,952
vomiting|952,960
,|960,961
diaphoresis|962,973
.|973,974
<EOL>|976,977
In|977,979
the|980,983
ED|984,986
,|986,987
initial|988,995
vitals|996,1002
were|1003,1007
:|1007,1008
98.0|1009,1013
50|1014,1016
156|1017,1020
/|1020,1021
73|1021,1023
20|1024,1026
99|1027,1029
%|1029,1030
<EOL>|1032,1033
-|1033,1034
Labs|1035,1039
were|1040,1044
significant|1045,1056
for|1057,1060
:|1060,1061
<EOL>|1063,1064
-|1064,1065
Na|1066,1068
137|1069,1072
K|1073,1074
3.0|1075,1078
Cl|1079,1081
94|1082,1084
CO2|1085,1088
32|1089,1091
BUN|1092,1095
16|1096,1098
Cr|1099,1101
0.8|1102,1105
<EOL>|1107,1108
-|1108,1109
Ca|1110,1112
:|1112,1113
10.6|1114,1118
Mg|1119,1121
:|1121,1122
1.9|1123,1126
P|1127,1128
:|1128,1129
2.9|1130,1133
<EOL>|1135,1136
-|1136,1137
WBC|1138,1141
5.9|1142,1145
Hgb|1146,1149
13.6|1150,1154
Hct|1155,1158
41.1|1159,1163
Plt|1164,1167
238|1168,1171
<EOL>|1173,1174
-|1174,1175
_|1176,1177
_|1177,1178
_|1178,1179
:|1179,1180
10.7|1181,1185
PTT|1186,1189
:|1189,1190
28.7|1191,1195
INR|1196,1199
:|1199,1200
1.0|1201,1204
<EOL>|1206,1207
-|1207,1208
Lactate|1209,1216
:|1216,1217
2.0|1217,1220
<EOL>|1222,1223
-|1223,1224
Trop|1225,1229
-|1229,1230
T|1230,1231
:|1231,1232
<|1233,1234
0.01|1234,1238
<EOL>|1240,1241
-|1241,1242
Imaging|1243,1250
revealed|1251,1259
:|1259,1260
<EOL>|1262,1263
-|1263,1264
CXR|1265,1268
:|1268,1269
No|1270,1272
acute|1273,1278
cardiopulmonary|1279,1294
process|1295,1302
<EOL>|1304,1305
-|1305,1306
The|1307,1310
patient|1311,1318
was|1319,1322
given|1323,1328
:|1328,1329
PO|1330,1332
Aspirin|1333,1340
243|1341,1344
,|1344,1345
IH|1346,1348
Albuterol|1349,1358
0.083|1359,1364
%|1364,1365
<EOL>|1366,1367
Neb|1367,1370
,|1370,1371
IH|1372,1374
Ipratropium|1375,1386
Bromide|1387,1394
Neb|1395,1398
,|1398,1399
PO|1400,1402
Potassium|1403,1412
Chloride|1413,1421
40|1422,1424
mEq|1425,1428
,|1428,1429
<EOL>|1430,1431
40|1431,1433
mEq|1434,1437
Potassium|1438,1447
Chloride|1448,1456
/|1457,1458
1000|1459,1463
mL|1464,1466
NS|1467,1469
<EOL>|1471,1472
-|1472,1473
Vitals|1474,1480
prior|1481,1486
to|1487,1489
transfer|1490,1498
were|1499,1503
:|1503,1504
98.1|1505,1509
84|1510,1512
163|1513,1516
/|1516,1517
118|1517,1520
17|1521,1523
100|1524,1527
%|1527,1528
RA|1529,1531
<EOL>|1533,1534
Upon|1534,1538
arrival|1539,1546
to|1547,1549
the|1550,1553
floor|1554,1559
,|1559,1560
patient|1561,1568
denies|1569,1575
chest|1576,1581
pain|1582,1586
,|1586,1587
shortness|1588,1597
<EOL>|1598,1599
of|1599,1601
breath|1602,1608
,|1608,1609
palpitations|1610,1622
,|1622,1623
lightheadedness|1624,1639
,|1639,1640
dizziness|1641,1650
.|1650,1651
<EOL>|1653,1654
REVIEW|1654,1660
OF|1661,1663
SYSTEMS|1664,1671
:|1671,1672
<EOL>|1674,1675
(|1675,1676
+|1676,1677
)|1677,1678
Per|1679,1682
HPI|1683,1686
<EOL>|1688,1689
<EOL>|1689,1690
<EOL>|1691,1692
ASTHMA|1714,1720
/|1720,1721
COPD|1721,1725
/|1725,1726
Tobacco|1726,1733
use|1734,1737
,|1737,1738
Peripheral|1739,1749
Arterial|1750,1758
disease|1759,1766
s|1767,1768
/|1768,1769
p|1769,1770
recent|1771,1777
<EOL>|1778,1779
common|1779,1785
iliac|1786,1791
stenting|1792,1800
,|1800,1801
ATRIAL|1802,1808
TACHYCARDIA|1809,1820
,|1820,1821
ATYPICAL|1822,1830
CHEST|1831,1836
PAIN|1837,1841
,|1841,1842
<EOL>|1843,1844
CERVICAL|1844,1852
RADICULITIS|1853,1864
,|1864,1865
CERVICAL|1866,1874
SPONDYLOSIS|1875,1886
,|1886,1887
CORONARY|1888,1896
ARTERY|1897,1903
<EOL>|1904,1905
DISEASE|1905,1912
<EOL>|1914,1915
HEADACHE|1915,1923
,|1923,1924
HIP|1925,1928
REPLACEMENT|1929,1940
,|1940,1941
HYPERLIPIDEMIA|1942,1956
,|1956,1957
HYPERTENSION|1958,1970
,|1970,1971
<EOL>|1972,1973
OSTEOARTHRITIS|1973,1987
,|1987,1988
HERPES|1989,1995
ZOSTER|1996,2002
,|2002,2003
TOBACCO|2004,2011
ABUSE|2012,2017
,|2017,2018
ATRIAL|2019,2025
<EOL>|2026,2027
FIBRILLATION|2027,2039
<EOL>|2041,2042
ANXIETY|2042,2049
,|2049,2050
GASTROINTESTINAL|2050,2066
BLEEDING|2067,2075
,|2075,2076
OSTEOARTHRITIS|2077,2091
,|2091,2092
<EOL>|2093,2094
ATHEROSCLEROTIC|2094,2109
CARDIOVASCULAR|2110,2124
DISEASE|2125,2132
,|2132,2133
PERIPHERAL|2134,2144
VASCULAR|2145,2153
<EOL>|2154,2155
DISEASE|2155,2162
,|2162,2163
CATARACT|2164,2172
SURGERY|2173,2180
_|2181,2182
_|2182,2183
_|2183,2184
<EOL>|2186,2187
Surgery|2187,2194
:|2194,2195
<EOL>|2197,2198
BILATERAL|2198,2207
COMMON|2208,2214
ILIAC|2215,2220
ARTERY|2221,2227
STENTING|2228,2236
_|2237,2238
_|2238,2239
_|2239,2240
<EOL>|2242,2243
BUNIONECTOMY|2243,2255
<EOL>|2257,2258
HIP|2258,2261
REPLACEMENT|2262,2273
<EOL>|2275,2276
PRIOR|2276,2281
CESAREAN|2282,2290
SECTION|2291,2298
<EOL>|2300,2301
GANGLION|2301,2309
CYST|2310,2314
<EOL>|2314,2315
<EOL>|2316,2317
:|2331,2332
<EOL>|2332,2333
_|2333,2334
_|2334,2335
_|2335,2336
<EOL>|2336,2337
:|2351,2352
<EOL>|2352,2353
Mother|2353,2359
:|2359,2360
_|2361,2362
_|2362,2363
_|2363,2364
,|2364,2365
HTN|2366,2369
<EOL>|2371,2372
Father|2372,2378
:|2378,2379
_|2380,2381
_|2381,2382
_|2382,2383
CA|2384,2386
<EOL>|2388,2389
Brother|2389,2396
:|2396,2397
CA|2398,2400
?|2400,2401
<EOL>|2403,2404
Brother|2404,2411
:|2411,2412
_|2413,2414
_|2414,2415
_|2415,2416
<EOL>|2417,2418
<EOL>|2419,2420
Physical|2420,2428
_|2429,2430
_|2430,2431
_|2431,2432
:|2432,2433
<EOL>|2433,2434
Admission|2434,2443
PE|2444,2446
:|2446,2447
<EOL>|2447,2448
Vitals|2448,2454
:|2454,2455
98.4|2456,2460
159|2461,2464
/|2464,2465
66|2465,2467
91|2468,2470
16|2471,2473
93|2474,2476
%|2476,2477
RA|2478,2480
Wt|2483,2485
:|2485,2486
66.2|2487,2491
<EOL>|2491,2492
General|2492,2499
:|2499,2500
Alert|2501,2506
,|2506,2507
oriented|2508,2516
,|2516,2517
no|2518,2520
acute|2521,2526
distress|2527,2535
<EOL>|2537,2538
HEENT|2538,2543
:|2543,2544
Sclera|2545,2551
anicteric|2552,2561
,|2561,2562
MMM|2563,2566
,|2566,2567
oropharynx|2568,2578
clear|2579,2584
,|2584,2585
EOMI|2586,2590
,|2590,2591
PERRL|2592,2597
<EOL>|2599,2600
Neck|2600,2604
:|2604,2605
Supple|2606,2612
,|2612,2613
JVP|2614,2617
not|2618,2621
elevated|2622,2630
,|2630,2631
no|2632,2634
LAD|2635,2638
<EOL>|2640,2641
CV|2641,2643
:|2643,2644
Regular|2645,2652
rate|2653,2657
and|2658,2661
rhythm|2662,2668
,|2668,2669
normal|2670,2676
S1|2677,2679
+|2680,2681
S2|2682,2684
,|2684,2685
_|2686,2687
_|2687,2688
_|2688,2689
systolic|2690,2698
murmur|2699,2705
<EOL>|2706,2707
heard|2707,2712
best|2713,2717
at|2718,2720
RUSB|2721,2725
,|2725,2726
no|2727,2729
rubs|2730,2734
or|2735,2737
gallops|2738,2745
<EOL>|2747,2748
Lungs|2748,2753
:|2753,2754
inspiratory|2755,2766
and|2767,2770
expiratory|2771,2781
wheezes|2782,2789
,|2789,2790
no|2791,2793
rales|2794,2799
or|2800,2802
rhonchi|2803,2810
<EOL>|2812,2813
Abdomen|2813,2820
:|2820,2821
Soft|2822,2826
,|2826,2827
non-tender|2828,2838
,|2838,2839
non-distended|2840,2853
,|2853,2854
bowel|2855,2860
sounds|2861,2867
present|2868,2875
,|2875,2876
<EOL>|2877,2878
no|2878,2880
organomegaly|2881,2893
,|2893,2894
no|2895,2897
rebound|2898,2905
or|2906,2908
guarding|2909,2917
<EOL>|2919,2920
GU|2920,2922
:|2922,2923
No|2924,2926
foley|2927,2932
<EOL>|2934,2935
Ext|2935,2938
:|2938,2939
Warm|2940,2944
,|2944,2945
well|2946,2950
perfused|2951,2959
,|2959,2960
2|2961,2962
+|2962,2963
pulses|2964,2970
,|2970,2971
no|2972,2974
clubbing|2975,2983
,|2983,2984
cyanosis|2985,2993
or|2994,2996
<EOL>|2997,2998
edema|2998,3003
<EOL>|3003,3004
<EOL>|3004,3005
Discharge|3005,3014
PE|3015,3017
:|3017,3018
<EOL>|3018,3019
Vitals|3019,3025
:|3025,3026
98.5|3027,3031
_|3032,3033
_|3033,3034
_|3034,3035
20|3036,3038
_|3039,3040
_|3040,3041
_|3041,3042
98|3043,3045
%|3045,3046
RA|3046,3048
<EOL>|3049,3050
Weight|3050,3056
:|3056,3057
64.5|3058,3062
<EOL>|3062,3063
Weight|3063,3069
on|3070,3072
admission|3073,3082
:|3082,3083
66.2|3084,3088
<EOL>|3088,3089
General|3089,3096
:|3096,3097
NAD|3098,3101
<EOL>|3102,3103
HEENT|3103,3108
:|3108,3109
Sclera|3110,3116
anicteric|3117,3126
<EOL>|3127,3128
Neck|3128,3132
:|3132,3133
JVP|3134,3137
not|3138,3141
elevated|3142,3150
<EOL>|3152,3153
CV|3153,3155
:|3155,3156
Regular|3157,3164
rhythm|3165,3171
with|3172,3176
frequent|3177,3185
skipped|3186,3193
beats|3194,3199
,|3199,3200
normal|3201,3207
S1|3208,3210
+|3211,3212
S2|3213,3215
,|3215,3216
<EOL>|3217,3218
_|3218,3219
_|3219,3220
_|3220,3221
systolic|3222,3230
murmur|3231,3237
heard|3238,3243
best|3244,3248
at|3249,3251
RUSB|3252,3256
,|3256,3257
no|3258,3260
rubs|3261,3265
or|3266,3268
gallops|3269,3276
<EOL>|3278,3279
Lungs|3279,3284
:|3284,3285
mild|3286,3290
expiratory|3291,3301
wheezes|3302,3309
,|3309,3310
diffuse|3311,3318
mild|3319,3323
rhonchi|3324,3331
<EOL>|3332,3333
(|3333,3334
pre-nebulizer|3334,3347
)|3347,3348
<EOL>|3349,3350
Abdomen|3350,3357
:|3357,3358
Soft|3359,3363
,|3363,3364
non-tender|3365,3375
,|3375,3376
non-distended|3377,3390
,|3390,3391
bowel|3392,3397
sounds|3398,3404
present|3405,3412
,|3412,3413
<EOL>|3414,3415
no|3415,3417
organomegaly|3418,3430
,|3430,3431
no|3432,3434
rebound|3435,3442
or|3443,3445
guarding|3446,3454
<EOL>|3457,3458
Ext|3458,3461
:|3461,3462
Warm|3463,3467
,|3467,3468
well|3469,3473
perfused|3474,3482
,|3482,3483
no|3484,3486
edema|3487,3492
<EOL>|3493,3494
<EOL>|3494,3495
<EOL>|3496,3497
Pertinent|3497,3506
Results|3507,3514
:|3514,3515
<EOL>|3515,3516
Admission|3516,3525
Labs|3526,3530
:|3530,3531
<EOL>|3532,3533
<EOL>|3533,3534
_|3534,3535
_|3535,3536
_|3536,3537
07|3538,3540
:|3540,3541
49PM|3541,3545
_|3548,3549
_|3549,3550
_|3550,3551
PTT|3552,3555
-|3555,3556
28.7|3556,3560
_|3561,3562
_|3562,3563
_|3563,3564
<EOL>|3564,3565
_|3565,3566
_|3566,3567
_|3567,3568
07|3569,3571
:|3571,3572
05PM|3572,3576
LACTATE|3579,3586
-|3586,3587
2.0|3587,3590
<EOL>|3590,3591
_|3591,3592
_|3592,3593
_|3593,3594
05|3595,3597
:|3597,3598
58PM|3598,3602
GLUCOSE|3605,3612
-|3612,3613
103|3613,3616
*|3616,3617
UREA|3618,3622
N|3623,3624
-|3624,3625
16|3625,3627
CREAT|3628,3633
-|3633,3634
0.8|3634,3637
SODIUM|3638,3644
-|3644,3645
137|3645,3648
<EOL>|3649,3650
POTASSIUM|3650,3659
-|3659,3660
3|3660,3661
.|3661,3662
0|3662,3663
*|3663,3664
CHLORIDE|3665,3673
-|3673,3674
94|3674,3676
*|3676,3677
TOTAL|3678,3683
CO2|3684,3687
-|3687,3688
32|3688,3690
ANION|3691,3696
GAP|3697,3700
-|3700,3701
14|3701,3703
<EOL>|3703,3704
_|3704,3705
_|3705,3706
_|3706,3707
05|3708,3710
:|3710,3711
58PM|3711,3715
estGFR|3718,3724
-|3724,3725
Using|3725,3730
this|3731,3735
<EOL>|3735,3736
_|3736,3737
_|3737,3738
_|3738,3739
05|3740,3742
:|3742,3743
58PM|3743,3747
cTropnT|3750,3757
-|3757,3758
<|3758,3759
0|3759,3760
.|3760,3761
01|3761,3763
<EOL>|3763,3764
_|3764,3765
_|3765,3766
_|3766,3767
05|3768,3770
:|3770,3771
58PM|3771,3775
CALCIUM|3778,3785
-|3785,3786
10|3786,3788
.|3788,3789
6|3789,3790
*|3790,3791
PHOSPHATE|3792,3801
-|3801,3802
2.9|3802,3805
MAGNESIUM|3806,3815
-|3815,3816
1.9|3816,3819
<EOL>|3819,3820
_|3820,3821
_|3821,3822
_|3822,3823
05|3824,3826
:|3826,3827
58PM|3827,3831
WBC|3834,3837
-|3837,3838
5.9|3838,3841
RBC|3842,3845
-|3845,3846
4|3846,3847
.|3847,3848
62|3848,3850
HGB|3851,3854
-|3854,3855
13.6|3855,3859
HCT|3860,3863
-|3863,3864
41.1|3864,3868
MCV|3869,3872
-|3872,3873
89|3873,3875
<EOL>|3876,3877
MCH|3877,3880
-|3880,3881
29.4|3881,3885
MCHC|3886,3890
-|3890,3891
33.1|3891,3895
RDW|3896,3899
-|3899,3900
14.7|3900,3904
RDWSD|3905,3910
-|3910,3911
47|3911,3913
.|3913,3914
1|3914,3915
*|3915,3916
<EOL>|3916,3917
_|3917,3918
_|3918,3919
_|3919,3920
05|3921,3923
:|3923,3924
58PM|3924,3928
NEUTS|3931,3936
-|3936,3937
57.8|3937,3941
_|3942,3943
_|3943,3944
_|3944,3945
MONOS|3946,3951
-|3951,3952
9.3|3952,3955
EOS|3956,3959
-|3959,3960
0|3960,3961
.|3961,3962
3|3962,3963
*|3963,3964
<EOL>|3965,3966
BASOS|3966,3971
-|3971,3972
0.2|3972,3975
IM|3976,3978
_|3979,3980
_|3980,3981
_|3981,3982
AbsNeut|3983,3990
-|3990,3991
3|3991,3992
.|3992,3993
41|3993,3995
AbsLymp|3996,4003
-|4003,4004
1|4004,4005
.|4005,4006
88|4006,4008
AbsMono|4009,4016
-|4016,4017
0|4017,4018
.|4018,4019
55|4019,4021
<EOL>|4022,4023
AbsEos|4023,4029
-|4029,4030
0|4030,4031
.|4031,4032
02|4032,4034
*|4034,4035
AbsBaso|4036,4043
-|4043,4044
0.01|4044,4048
<EOL>|4048,4049
_|4049,4050
_|4050,4051
_|4051,4052
05|4053,4055
:|4055,4056
58PM|4056,4060
PLT|4063,4066
COUNT|4067,4072
-|4072,4073
238|4073,4076
<EOL>|4076,4077
<EOL>|4077,4078
Discharge|4078,4087
Labs|4088,4092
:|4092,4093
<EOL>|4093,4094
<EOL>|4094,4095
_|4095,4096
_|4096,4097
_|4097,4098
06|4099,4101
:|4101,4102
20AM|4102,4106
BLOOD|4107,4112
WBC|4113,4116
-|4116,4117
6.1|4117,4120
RBC|4121,4124
-|4124,4125
4|4125,4126
.|4126,4127
60|4127,4129
Hgb|4130,4133
-|4133,4134
13.4|4134,4138
Hct|4139,4142
-|4142,4143
41.2|4143,4147
MCV|4148,4151
-|4151,4152
90|4152,4154
<EOL>|4155,4156
MCH|4156,4159
-|4159,4160
29.1|4160,4164
MCHC|4165,4169
-|4169,4170
32.5|4170,4174
RDW|4175,4178
-|4178,4179
14.9|4179,4183
RDWSD|4184,4189
-|4189,4190
47|4190,4192
.|4192,4193
8|4193,4194
*|4194,4195
Plt|4196,4199
_|4200,4201
_|4201,4202
_|4202,4203
<EOL>|4203,4204
_|4204,4205
_|4205,4206
_|4206,4207
06|4208,4210
:|4210,4211
20AM|4211,4215
BLOOD|4216,4221
Plt|4222,4225
_|4226,4227
_|4227,4228
_|4228,4229
<EOL>|4229,4230
_|4230,4231
_|4231,4232
_|4232,4233
06|4234,4236
:|4236,4237
20AM|4237,4241
BLOOD|4242,4247
Glucose|4248,4255
-|4255,4256
97|4256,4258
UreaN|4259,4264
-|4264,4265
17|4265,4267
Creat|4268,4273
-|4273,4274
1.0|4274,4277
Na|4278,4280
-|4280,4281
134|4281,4284
<EOL>|4285,4286
K|4286,4287
-|4287,4288
4.2|4288,4291
Cl|4292,4294
-|4294,4295
96|4295,4297
HCO3|4298,4302
-|4302,4303
24|4303,4305
AnGap|4306,4311
-|4311,4312
18|4312,4314
<EOL>|4314,4315
_|4315,4316
_|4316,4317
_|4317,4318
06|4319,4321
:|4321,4322
25AM|4322,4326
BLOOD|4327,4332
ALT|4333,4336
-|4336,4337
19|4337,4339
AST|4340,4343
-|4343,4344
22|4344,4346
LD|4347,4349
(|4349,4350
LDH|4350,4353
)|4353,4354
-|4354,4355
260|4355,4358
*|4358,4359
AlkPhos|4360,4367
-|4367,4368
81|4368,4370
<EOL>|4371,4372
TotBili|4372,4379
-|4379,4380
0.4|4380,4383
<EOL>|4383,4384
_|4384,4385
_|4385,4386
_|4386,4387
06|4388,4390
:|4390,4391
20AM|4391,4395
BLOOD|4396,4401
Calcium|4402,4409
-|4409,4410
9.7|4410,4413
Phos|4414,4418
-|4418,4419
3.7|4419,4422
Mg|4423,4425
-|4425,4426
1.9|4426,4429
<EOL>|4429,4430
<EOL>|4430,4431
Studies|4431,4438
:|4438,4439
<EOL>|4439,4440
1.|4440,4442
CXR|4443,4446
_|4447,4448
_|4448,4449
_|4449,4450
:|4450,4451
No|4452,4454
acute|4455,4460
cardiopulmonary|4461,4476
process|4477,4484
<EOL>|4486,4487
2.|4487,4489
_|4490,4491
_|4491,4492
_|4492,4493
:|4493,4494
Exercise|4495,4503
stress|4504,4510
test|4511,4515
<EOL>|4517,4518
INTERPRETATION|4518,4532
:|4532,4533
This|4534,4538
_|4539,4540
_|4540,4541
_|4541,4542
year|4543,4547
old|4548,4551
woman|4552,4557
with|4558,4562
a|4563,4564
history|4565,4572
of|4573,4575
PAD|4576,4579
and|4580,4583
<EOL>|4584,4585
<EOL>|4586,4587
LBBB|4587,4591
was|4592,4595
referred|4596,4604
to|4605,4607
the|4608,4611
lab|4612,4615
from|4616,4620
the|4621,4624
ER|4625,4627
following|4628,4637
negative|4638,4646
<EOL>|4647,4648
serial|4648,4654
<EOL>|4656,4657
cardiac|4657,4664
markers|4665,4672
for|4673,4676
evaluation|4677,4687
of|4688,4690
chest|4691,4696
discomfort|4697,4707
.|4707,4708
The|4709,4712
patient|4713,4720
<EOL>|4721,4722
was|4722,4725
<EOL>|4727,4728
referred|4728,4736
for|4737,4740
a|4741,4742
dipyridamole|4743,4755
stress|4756,4762
test|4763,4767
but|4768,4771
due|4772,4775
to|4776,4778
her|4779,4782
<EOL>|4783,4784
theophylline|4784,4796
<EOL>|4798,4799
therapy|4799,4806
we|4807,4809
were|4810,4814
not|4815,4818
able|4819,4823
to|4824,4826
proceed|4827,4834
.|4834,4835
Due|4836,4839
to|4840,4842
her|4843,4846
frequent|4847,4855
atrial|4856,4862
<EOL>|4863,4864
ectopy|4864,4870
we|4871,4873
chose|4874,4879
not|4880,4883
to|4884,4886
give|4887,4891
her|4892,4895
dobutamine|4896,4906
but|4907,4910
had|4911,4914
her|4915,4918
walk|4919,4923
on|4924,4926
<EOL>|4927,4928
the|4928,4931
treadmill|4932,4941
instead|4942,4949
.|4949,4950
She|4951,4954
exercised|4955,4964
for|4965,4968
3|4969,4970
minutes|4971,4978
of|4979,4981
a|4982,4983
modified|4984,4992
<EOL>|4993,4994
_|4994,4995
_|4995,4996
_|4996,4997
protocol|4998,5006
and|5007,5010
stopped|5011,5018
due|5019,5022
to|5023,5025
leg|5026,5029
claudication|5030,5042
.|5042,5043
The|5044,5047
<EOL>|5048,5049
estimated|5049,5058
peak|5059,5063
MET|5064,5067
capacity|5068,5076
was|5077,5080
2.5|5081,5084
which|5085,5090
represents|5091,5101
a|5102,5103
poor|5104,5108
<EOL>|5109,5110
functional|5110,5120
capacity|5121,5129
for|5130,5133
her|5134,5137
age|5138,5141
.|5141,5142
No|5143,5145
arm|5146,5149
,|5149,5150
neck|5151,5155
,|5155,5156
back|5157,5161
or|5162,5164
chest|5165,5170
<EOL>|5171,5172
discomfort|5172,5182
was|5183,5186
reported|5187,5195
by|5196,5198
the|5199,5202
patient|5203,5210
throughout|5211,5221
the|5222,5225
study|5226,5231
.|5231,5232
The|5233,5236
<EOL>|5237,5238
ST|5238,5240
segments|5241,5249
are|5250,5253
uninterpretable|5254,5269
for|5270,5273
ischemia|5274,5282
in|5283,5285
the|5286,5289
setting|5290,5297
of|5298,5300
<EOL>|5301,5302
the|5302,5305
baseline|5306,5314
LBBB|5315,5319
.|5319,5320
The|5321,5324
rhythm|5325,5331
was|5332,5335
sinus|5336,5341
with|5342,5346
frequent|5347,5355
isolated|5356,5364
<EOL>|5365,5366
apbs|5366,5370
,|5370,5371
occasional|5372,5382
atrial|5383,5389
couplets|5390,5398
and|5399,5402
a|5403,5404
6|5405,5406
beat|5407,5411
run|5412,5415
of|5416,5418
PSVT|5419,5423
.|5423,5424
Rare|5425,5429
<EOL>|5430,5431
isolated|5431,5439
vpbs|5440,5444
were|5445,5449
also|5450,5454
noted|5455,5460
.|5460,5461
Resting|5462,5469
mild|5470,5474
systolic|5475,5483
<EOL>|5484,5485
hypertension|5485,5497
with|5498,5502
a|5503,5504
pprorpriate|5505,5516
increase|5517,5525
in|5526,5528
BP|5529,5531
with|5532,5536
exercise|5537,5545
and|5546,5549
<EOL>|5550,5551
recovery|5551,5559
.|5559,5560
<EOL>|5562,5563
IMPRESSION|5563,5573
:|5573,5574
No|5575,5577
anginal|5578,5585
type|5586,5590
symptoms|5591,5599
or|5600,5602
interpretable|5603,5616
ST|5617,5619
<EOL>|5620,5621
segments|5621,5629
at|5630,5632
a|5633,5634
high|5635,5639
cardiac|5640,5647
demand|5648,5654
and|5655,5658
poor|5659,5663
functional|5664,5674
capacity|5675,5683
.|5683,5684
<EOL>|5685,5686
Nuclear|5686,5693
report|5694,5700
sent|5701,5705
separately|5706,5716
.|5716,5717
<EOL>|5719,5720
3.|5720,5722
_|5723,5724
_|5724,5725
_|5725,5726
CATH|5727,5731
:|5731,5732
<EOL>|5734,5735
LMCA|5735,5739
:|5739,5740
short|5741,5746
,|5746,5747
no|5748,5750
CAD|5751,5754
.|5754,5755
LAD|5756,5759
:|5759,5760
mild|5761,5765
<EOL>|5767,5768
focal|5768,5773
origin|5774,5780
disease|5781,5788
(|5789,5790
20|5790,5792
%|5792,5793
)|5793,5794
and|5795,5798
mild|5799,5803
proximal|5804,5812
disease|5813,5820
(|5821,5822
30|5822,5824
%|5824,5825
)|5825,5826
.|5826,5827
LCX|5828,5831
:|5831,5832
<EOL>|5833,5834
<EOL>|5835,5836
minimal|5836,5843
luminal|5844,5851
irregularities|5852,5866
.|5866,5867
RCA|5868,5871
:|5871,5872
30|5873,5875
%|5875,5876
.|5876,5877
<EOL>|5879,5880
4.|5880,5882
ECG|5883,5886
_|5887,5888
_|5888,5889
_|5889,5890
:|5890,5891
sinus|5892,5897
rhythm|5898,5904
with|5905,5909
multiple|5910,5918
PACs|5919,5923
,|5923,5924
left|5925,5929
axis|5930,5934
<EOL>|5935,5936
deviation|5936,5945
,|5945,5946
old|5947,5950
LBBB|5951,5955
<EOL>|5956,5957
5.|5957,5959
ECG|5960,5963
_|5964,5965
_|5965,5966
_|5966,5967
:|5967,5968
Likely|5969,5975
atrial|5976,5982
tachycardia|5983,5994
.|5994,5995
Left|5996,6000
bundle|6001,6007
-|6007,6008
branch|6008,6014
<EOL>|6015,6016
block|6016,6021
.|6021,6022
Compared|6023,6031
to|6032,6034
the|6035,6038
previous|6039,6047
tracing|6048,6055
atrial|6056,6062
tachycardia|6063,6074
has|6075,6078
<EOL>|6079,6080
replaced|6080,6088
sinus|6089,6094
rhythm|6095,6101
with|6102,6106
premature|6107,6116
atrial|6117,6123
contractions|6124,6136
.|6136,6137
Left|6138,6142
<EOL>|6143,6144
bundle|6144,6150
-|6150,6151
branch|6151,6157
block|6158,6163
was|6164,6167
previously|6168,6178
noted|6179,6184
.|6184,6185
<EOL>|6186,6187
6.|6187,6189
ECHO|6190,6194
_|6195,6196
_|6196,6197
_|6197,6198
:|6198,6199
Conclusions|6200,6211
<EOL>|6213,6214
The|6214,6217
left|6218,6222
atrium|6223,6229
is|6230,6232
normal|6233,6239
in|6240,6242
size|6243,6247
.|6247,6248
No|6249,6251
atrial|6252,6258
septal|6259,6265
defect|6266,6272
is|6273,6275
<EOL>|6276,6277
seen|6277,6281
by|6282,6284
2D|6285,6287
or|6288,6290
color|6291,6296
Doppler|6297,6304
.|6304,6305
The|6306,6309
estimated|6310,6319
right|6320,6325
atrial|6326,6332
pressure|6333,6341
<EOL>|6342,6343
is|6343,6345
_|6346,6347
_|6347,6348
_|6348,6349
mmHg|6350,6354
.|6354,6355
Left|6356,6360
ventricular|6361,6372
wall|6373,6377
thickness|6378,6387
,|6387,6388
cavity|6389,6395
size|6396,6400
and|6401,6404
<EOL>|6405,6406
regional|6406,6414
/|6414,6415
global|6415,6421
systolic|6422,6430
function|6431,6439
are|6440,6443
normal|6444,6450
(|6451,6452
LVEF|6452,6456
>|6457,6458
55|6458,6460
%|6460,6461
)|6461,6462
.|6462,6463
There|6464,6469
<EOL>|6470,6471
is|6471,6473
considerable|6474,6486
beat|6487,6491
-|6491,6492
to|6492,6494
-|6494,6495
beat|6495,6499
variability|6500,6511
of|6512,6514
the|6515,6518
left|6519,6523
ventricular|6524,6535
<EOL>|6536,6537
ejection|6537,6545
fraction|6546,6554
due|6555,6558
to|6559,6561
an|6562,6564
irregular|6565,6574
rhythm|6575,6581
/|6581,6582
premature|6582,6591
beats|6592,6597
.|6597,6598
<EOL>|6599,6600
Tissue|6600,6606
Doppler|6607,6614
imaging|6615,6622
suggests|6623,6631
a|6632,6633
normal|6634,6640
left|6641,6645
ventricular|6646,6657
<EOL>|6658,6659
filling|6659,6666
pressure|6667,6675
(|6676,6677
PCWP|6677,6681
<|6681,6682
12mmHg|6682,6688
)|6688,6689
.|6689,6690
Right|6691,6696
ventricular|6697,6708
chamber|6709,6716
size|6717,6721
<EOL>|6722,6723
and|6723,6726
free|6727,6731
wall|6732,6736
motion|6737,6743
are|6744,6747
normal|6748,6754
.|6754,6755
The|6756,6759
aortic|6760,6766
valve|6767,6772
leaflets|6773,6781
are|6782,6785
<EOL>|6786,6787
mildly|6787,6793
thickened|6794,6803
(|6804,6805
?|6805,6806
#|6806,6807
)|6807,6808
.|6808,6809
There|6810,6815
is|6816,6818
no|6819,6821
aortic|6822,6828
valve|6829,6834
stenosis|6835,6843
.|6843,6844
No|6845,6847
<EOL>|6848,6849
aortic|6849,6855
regurgitation|6856,6869
is|6870,6872
seen|6873,6877
.|6877,6878
The|6879,6882
mitral|6883,6889
valve|6890,6895
leaflets|6896,6904
are|6905,6908
<EOL>|6909,6910
mildly|6910,6916
thickened|6917,6926
.|6926,6927
There|6928,6933
is|6934,6936
no|6937,6939
mitral|6940,6946
valve|6947,6952
prolapse|6953,6961
.|6961,6962
Physiologic|6963,6974
<EOL>|6975,6976
mitral|6976,6982
regurgitation|6983,6996
is|6997,6999
seen|7000,7004
(|7005,7006
within|7006,7012
normal|7013,7019
limits|7020,7026
)|7026,7027
.|7027,7028
The|7029,7032
left|7033,7037
<EOL>|7038,7039
ventricular|7039,7050
inflow|7051,7057
pattern|7058,7065
suggests|7066,7074
impaired|7075,7083
relaxation|7084,7094
.|7094,7095
The|7096,7099
<EOL>|7100,7101
estimated|7101,7110
pulmonary|7111,7120
artery|7121,7127
systolic|7128,7136
pressure|7137,7145
is|7146,7148
normal|7149,7155
.|7155,7156
There|7157,7162
is|7163,7165
<EOL>|7166,7167
no|7167,7169
pericardial|7170,7181
effusion|7182,7190
.|7190,7191
<EOL>|7192,7193
Compared|7193,7201
with|7202,7206
the|7207,7210
prior|7211,7216
study|7217,7222
(|7223,7224
images|7224,7230
reviewed|7231,7239
)|7239,7240
of|7241,7243
_|7244,7245
_|7245,7246
_|7246,7247
,|7247,7248
<EOL>|7249,7250
frequent|7250,7258
atrial|7259,7265
ectopy|7266,7272
is|7273,7275
seen|7276,7280
;|7280,7281
biventricular|7282,7295
function|7296,7304
appears|7305,7312
<EOL>|7313,7314
similar|7314,7321
.|7321,7322
<EOL>|7325,7326
<EOL>|7326,7327
Micro|7327,7332
:|7332,7333
_|7334,7335
_|7335,7336
_|7336,7337
:|7337,7338
Bcx|7339,7342
pending|7343,7350
<EOL>|7350,7351
<EOL>|7352,7353
<EOL>|7375,7376
=|7398,7399
=|7399,7400
=|7400,7401
=|7401,7402
=|7402,7403
=|7403,7404
=|7404,7405
=|7405,7406
=|7406,7407
=|7407,7408
=|7408,7409
=|7409,7410
=|7410,7411
=|7411,7412
=|7412,7413
=|7413,7414
=|7414,7415
=|7415,7416
=|7416,7417
=|7417,7418
=|7418,7419
=|7419,7420
=|7420,7421
=|7421,7422
=|7422,7423
=|7423,7424
=|7424,7425
=|7425,7426
=|7426,7427
=|7427,7428
=|7428,7429
=|7429,7430
=|7430,7431
=|7431,7432
=|7432,7433
=|7433,7434
=|7434,7435
=|7435,7436
=|7436,7437
=|7437,7438
=|7438,7439
=|7439,7440
=|7440,7441
=|7441,7442
=|7442,7443
=|7443,7444
=|7444,7445
=|7445,7446
=|7446,7447
=|7447,7448
=|7448,7449
=|7449,7450
=|7450,7451
=|7451,7452
=|7452,7453
=|7453,7454
=|7454,7455
=|7455,7456
=|7456,7457
<EOL>|7457,7458
_|7458,7459
_|7459,7460
_|7460,7461
PMH|7462,7465
of|7466,7468
CAD|7469,7472
,|7472,7473
PVD|7474,7477
,|7477,7478
and|7479,7482
COPD|7483,7487
presenting|7488,7498
with|7499,7503
recurrent|7504,7513
<EOL>|7514,7515
non-exertional|7515,7529
substernal|7530,7540
chest|7541,7546
pain|7547,7551
.|7551,7552
The|7553,7556
patient|7557,7564
has|7565,7568
a|7569,7570
history|7571,7578
<EOL>|7579,7580
of|7580,7582
mild|7583,7587
CAD|7588,7591
but|7592,7595
labs|7596,7600
were|7601,7605
significant|7606,7617
for|7618,7621
negative|7622,7630
troponins|7631,7640
and|7641,7644
<EOL>|7645,7646
EKG|7646,7649
was|7650,7653
without|7654,7661
ischemic|7662,7670
changes|7671,7678
.|7678,7679
During|7680,7686
her|7687,7690
admission|7691,7700
,|7700,7701
she|7702,7705
also|7706,7710
<EOL>|7711,7712
developed|7712,7721
multiple|7722,7730
episodes|7731,7739
of|7740,7742
atrial|7743,7749
tachycardia|7750,7761
(|7762,7763
AFib|7763,7767
vs|7768,7770
.|7770,7771
<EOL>|7772,7773
Aflutter|7773,7781
)|7781,7782
and|7783,7786
was|7787,7790
started|7791,7798
on|7799,7801
Amiodarone|7802,7812
for|7813,7816
rate|7817,7821
/|7821,7822
rhythm|7822,7828
control|7829,7836
<EOL>|7837,7838
and|7838,7841
Rivaroxaban|7842,7853
for|7854,7857
anticoagulation|7858,7873
,|7873,7874
and|7875,7878
kept|7879,7883
on|7884,7886
home|7887,7891
dose|7892,7896
of|7897,7899
<EOL>|7900,7901
Diltiazem|7901,7910
also|7911,7915
for|7916,7919
rate|7920,7924
control|7925,7932
.|7932,7933
She|7934,7937
did|7938,7941
not|7942,7945
have|7946,7950
any|7951,7954
episodes|7955,7963
<EOL>|7964,7965
of|7965,7967
chest|7968,7973
pain|7974,7978
during|7979,7985
hospitalization|7986,8001
,|8001,8002
so|8003,8005
was|8006,8009
discharged|8010,8020
once|8021,8025
<EOL>|8026,8027
atrial|8027,8033
fibrillation|8034,8046
/|8046,8047
flutter|8047,8054
was|8055,8058
controlled|8059,8069
.|8069,8070
She|8071,8074
will|8075,8079
need|8080,8084
to|8085,8087
<EOL>|8088,8089
follow|8089,8095
up|8096,8098
with|8099,8103
her|8104,8107
primary|8108,8115
care|8116,8120
doctor|8121,8127
regarding|8128,8137
vague|8138,8143
chest|8144,8149
<EOL>|8150,8151
pain|8151,8155
which|8156,8161
led|8162,8165
to|8166,8168
admission|8169,8178
.|8178,8179
<EOL>|8179,8180
<EOL>|8180,8181
Acute|8181,8186
Issues|8187,8193
:|8193,8194
<EOL>|8194,8195
=|8195,8196
=|8196,8197
=|8197,8198
=|8198,8199
=|8199,8200
=|8200,8201
=|8201,8202
=|8202,8203
=|8203,8204
=|8204,8205
=|8205,8206
=|8206,8207
=|8207,8208
=|8208,8209
=|8209,8210
=|8210,8211
=|8211,8212
=|8212,8213
=|8213,8214
=|8214,8215
=|8215,8216
=|8216,8217
=|8217,8218
=|8218,8219
=|8219,8220
=|8220,8221
=|8221,8222
=|8222,8223
=|8223,8224
=|8224,8225
=|8225,8226
=|8226,8227
=|8227,8228
=|8228,8229
=|8229,8230
=|8230,8231
=|8231,8232
=|8232,8233
=|8233,8234
=|8234,8235
=|8235,8236
=|8236,8237
=|8237,8238
=|8238,8239
=|8239,8240
=|8240,8241
=|8241,8242
=|8242,8243
=|8243,8244
=|8244,8245
=|8245,8246
=|8246,8247
=|8247,8248
=|8248,8249
=|8249,8250
=|8250,8251
<EOL>|8251,8252
#|8252,8253
Atrial|8253,8259
Tachycardia|8260,8271
:|8271,8272
During|8273,8279
admission|8280,8289
pt|8290,8292
had|8293,8296
runs|8297,8301
of|8302,8304
wide|8305,8309
<EOL>|8310,8311
complex|8311,8318
tachyarrythmia|8319,8333
,|8333,8334
thought|8335,8342
likely|8343,8349
supraventricular|8350,8366
in|8367,8369
<EOL>|8370,8371
origin|8371,8377
:|8377,8378
rapid|8379,8384
Atrial|8385,8391
Fibrillation|8392,8404
/|8404,8405
Flutter|8406,8413
vs|8414,8416
.|8416,8417
atrial|8418,8424
<EOL>|8425,8426
tachycardia|8426,8437
,|8437,8438
with|8439,8443
abberancy|8444,8453
(|8454,8455
complexes|8455,8464
with|8465,8469
similar|8470,8477
morphology|8478,8488
<EOL>|8489,8490
to|8490,8492
native|8493,8499
LBBB|8500,8504
)|8504,8505
.|8505,8506
She|8507,8510
was|8511,8514
treated|8515,8522
with|8523,8527
Diltiazem|8528,8537
and|8538,8541
Amiodarone|8542,8552
<EOL>|8553,8554
and|8554,8557
had|8558,8561
fewer|8562,8567
episodes|8568,8576
of|8577,8579
tachycardia|8580,8591
.|8591,8592
EP|8593,8595
team|8596,8600
evaluated|8601,8610
patient|8611,8618
<EOL>|8619,8620
and|8620,8623
recommended|8624,8635
anticoagulation|8636,8651
and|8652,8655
outpatient|8656,8666
follow|8667,8673
up|8674,8676
to|8677,8679
<EOL>|8680,8681
consider|8681,8689
EP|8690,8692
study|8693,8698
and|8699,8702
possible|8703,8711
ablation|8712,8720
of|8721,8723
Atrial|8724,8730
Flutter|8731,8738
.|8738,8739
<EOL>|8740,8741
Patient|8741,8748
was|8749,8752
discharged|8753,8763
with|8764,8768
_|8769,8770
_|8770,8771
_|8771,8772
of|8773,8775
Hearts|8776,8782
monitor|8783,8790
,|8790,8791
Amiodarone|8792,8802
<EOL>|8803,8804
200mg|8804,8809
twice|8810,8815
daily|8816,8821
x|8822,8823
1|8824,8825
week|8826,8830
followed|8831,8839
by|8840,8842
200|8843,8846
mg|8847,8849
daily|8850,8855
thereafter|8856,8866
.|8866,8867
<EOL>|8868,8869
Diltiazem|8869,8878
continued|8879,8888
at|8889,8891
home|8892,8896
dose|8897,8901
.|8901,8902
Rivaroxaban|8903,8914
added|8915,8920
for|8921,8924
<EOL>|8925,8926
anticoagulation|8926,8941
.|8941,8942
As|8943,8945
per|8946,8949
outpatient|8950,8960
cardiologist|8961,8973
(|8974,8975
Dr|8975,8977
.|8977,8978
_|8979,8980
_|8980,8981
_|8981,8982
,|8982,8983
<EOL>|8984,8985
plavix|8985,8991
was|8992,8995
discontinued|8996,9008
in|9009,9011
light|9012,9017
of|9018,9020
addition|9021,9029
of|9030,9032
Rivaroxaban|9033,9044
and|9045,9048
<EOL>|9049,9050
interest|9050,9058
in|9059,9061
avoiding|9062,9070
triple|9071,9077
therapy|9078,9085
in|9086,9088
this|9089,9093
patient|9094,9101
.|9101,9102
Pt|9103,9105
was|9106,9109
<EOL>|9110,9111
given|9111,9116
follow|9117,9123
up|9124,9126
appointments|9127,9139
with|9140,9144
Drs.|9145,9149
_|9150,9151
_|9151,9152
_|9152,9153
.|9153,9154
She|9155,9158
was|9159,9162
<EOL>|9163,9164
scheduled|9164,9173
to|9174,9176
see|9177,9180
Dr.|9181,9184
_|9185,9186
_|9186,9187
_|9187,9188
EP|9189,9191
evaluation|9192,9202
in|9203,9205
2|9206,9207
months|9208,9214
.|9214,9215
<EOL>|9215,9216
<EOL>|9216,9217
#|9217,9218
Chest|9218,9223
pain|9224,9228
:|9228,9229
Pt|9230,9232
presented|9233,9242
with|9243,9247
substernal|9248,9258
chest|9259,9264
pain|9265,9269
that|9270,9274
<EOL>|9275,9276
occurred|9276,9284
at|9285,9287
rest|9288,9292
and|9293,9296
was|9297,9300
ruled|9301,9306
out|9307,9310
for|9311,9314
MI|9315,9317
with|9318,9322
no|9323,9325
troponin|9326,9334
<EOL>|9335,9336
elevation|9336,9345
or|9346,9348
significant|9349,9360
new|9361,9364
ECG|9365,9368
changes|9369,9376
.|9376,9377
Likely|9378,9384
her|9385,9388
chest|9389,9394
pain|9395,9399
<EOL>|9400,9401
was|9401,9404
related|9405,9412
to|9413,9415
periods|9416,9423
of|9424,9426
tachycardia|9427,9438
,|9438,9439
although|9440,9448
while|9449,9454
in|9455,9457
the|9458,9461
<EOL>|9462,9463
hospital|9463,9471
the|9472,9475
runs|9476,9480
of|9481,9483
atrial|9484,9490
tachycardia|9491,9502
did|9503,9506
not|9507,9510
reproduce|9511,9520
chest|9521,9526
<EOL>|9527,9528
pain|9528,9532
.|9532,9533
She|9534,9537
did|9538,9541
not|9542,9545
have|9546,9550
any|9551,9554
episodes|9555,9563
of|9564,9566
chest|9567,9572
pain|9573,9577
during|9578,9584
<EOL>|9585,9586
hospitalization|9586,9601
,|9601,9602
so|9603,9605
was|9606,9609
discharged|9610,9620
once|9621,9625
atrial|9626,9632
<EOL>|9633,9634
fibrillation|9634,9646
/|9646,9647
flutter|9647,9654
was|9655,9658
controlled|9659,9669
.|9669,9670
She|9671,9674
will|9675,9679
need|9680,9684
to|9685,9687
follow|9688,9694
up|9695,9697
<EOL>|9698,9699
with|9699,9703
her|9704,9707
primary|9708,9715
care|9716,9720
doctor|9721,9727
regarding|9728,9737
vague|9738,9743
chest|9744,9749
pain|9750,9754
which|9755,9760
<EOL>|9761,9762
led|9762,9765
to|9766,9768
admission|9769,9778
.|9778,9779
<EOL>|9779,9780
<EOL>|9780,9781
#|9781,9782
Dry|9782,9785
eyes|9786,9790
:|9790,9791
pt|9792,9794
had|9795,9798
erythema|9799,9807
and|9808,9811
pain|9812,9816
of|9817,9819
R|9820,9821
eye|9822,9825
,|9825,9826
found|9827,9832
to|9833,9835
have|9836,9840
dry|9841,9844
<EOL>|9845,9846
eyes|9846,9850
per|9851,9854
optholmology|9855,9867
.|9867,9868
Sent|9869,9873
out|9874,9877
with|9878,9882
Artificial|9883,9893
tears|9894,9899
and|9900,9903
<EOL>|9904,9905
erythromycin|9905,9917
eye|9918,9921
drops|9922,9927
.|9927,9928
Patient|9929,9936
had|9937,9940
follow|9941,9947
up|9948,9950
appointment|9951,9962
<EOL>|9963,9964
already|9964,9971
scheduled|9972,9981
with|9982,9986
optholmology|9987,9999
and|10000,10003
was|10004,10007
instructed|10008,10018
to|10019,10021
attend|10022,10028
<EOL>|10029,10030
appointment|10030,10041
.|10041,10042
<EOL>|10042,10043
<EOL>|10043,10044
Chronic|10044,10051
Issues|10052,10058
:|10058,10059
<EOL>|10059,10060
=|10060,10061
=|10061,10062
=|10062,10063
=|10063,10064
=|10064,10065
=|10065,10066
=|10066,10067
=|10067,10068
=|10068,10069
=|10069,10070
=|10070,10071
=|10071,10072
=|10072,10073
=|10073,10074
=|10074,10075
=|10075,10076
=|10076,10077
=|10077,10078
=|10078,10079
=|10079,10080
=|10080,10081
=|10081,10082
=|10082,10083
=|10083,10084
=|10084,10085
=|10085,10086
=|10086,10087
=|10087,10088
=|10088,10089
=|10089,10090
=|10090,10091
=|10091,10092
=|10092,10093
=|10093,10094
=|10094,10095
=|10095,10096
=|10096,10097
=|10097,10098
=|10098,10099
=|10099,10100
=|10100,10101
=|10101,10102
=|10102,10103
=|10103,10104
=|10104,10105
=|10105,10106
=|10106,10107
=|10107,10108
=|10108,10109
=|10109,10110
=|10110,10111
=|10111,10112
=|10112,10113
=|10113,10114
=|10114,10115
=|10115,10116
=|10116,10117
=|10117,10118
=|10118,10119
=|10119,10120
=|10120,10121
<EOL>|10121,10122
#|10122,10123
COPD|10124,10128
Pt|10130,10132
appeared|10133,10141
to|10142,10144
be|10145,10147
at|10148,10150
baseline|10151,10159
respiratory|10160,10171
status|10172,10178
.|10178,10179
She|10180,10183
<EOL>|10184,10185
was|10185,10188
sent|10189,10193
home|10194,10198
with|10199,10203
her|10204,10207
home|10208,10212
albuterol|10213,10222
neb|10223,10226
,|10226,10227
albuterol|10228,10237
inhaler|10238,10245
,|10245,10246
<EOL>|10247,10248
Fluticasone|10248,10259
nasal|10260,10265
spray|10266,10271
,|10271,10272
fluticasone|10273,10284
-|10284,10285
salmeterol|10285,10295
diskus|10296,10302
,|10302,10303
<EOL>|10304,10305
tiotropium|10305,10315
bromide|10316,10323
nebs|10324,10328
,|10328,10329
and|10330,10333
theophylline|10334,10346
<EOL>|10346,10347
<EOL>|10347,10348
#|10348,10349
PAD|10350,10353
:|10353,10354
<EOL>|10355,10356
As|10356,10358
above|10359,10364
,|10364,10365
we|10366,10368
stopped|10369,10376
Clopidogrel|10377,10388
as|10389,10391
patient|10392,10399
is|10400,10402
now|10403,10406
on|10407,10409
<EOL>|10410,10411
Rivaroxaban|10411,10422
and|10423,10426
wanted|10427,10433
to|10434,10436
avoid|10437,10442
triple|10443,10449
therapy|10450,10457
as|10458,10460
per|10461,10464
her|10465,10468
<EOL>|10469,10470
cardiologist|10470,10482
Dr.|10483,10486
_|10487,10488
_|10488,10489
_|10489,10490
.|10490,10491
<EOL>|10491,10492
<EOL>|10492,10493
Transitional|10493,10505
Issues|10506,10512
:|10512,10513
<EOL>|10513,10514
=|10514,10515
=|10515,10516
=|10516,10517
=|10517,10518
=|10518,10519
=|10519,10520
=|10520,10521
=|10521,10522
=|10522,10523
=|10523,10524
=|10524,10525
=|10525,10526
=|10526,10527
=|10527,10528
=|10528,10529
=|10529,10530
=|10530,10531
=|10531,10532
=|10532,10533
=|10533,10534
=|10534,10535
=|10535,10536
=|10536,10537
=|10537,10538
=|10538,10539
=|10539,10540
=|10540,10541
=|10541,10542
=|10542,10543
=|10543,10544
=|10544,10545
=|10545,10546
=|10546,10547
=|10547,10548
=|10548,10549
=|10549,10550
=|10550,10551
=|10551,10552
=|10552,10553
=|10553,10554
=|10554,10555
=|10555,10556
=|10556,10557
=|10557,10558
=|10558,10559
=|10559,10560
=|10560,10561
=|10561,10562
=|10562,10563
=|10563,10564
=|10564,10565
=|10565,10566
=|10566,10567
=|10567,10568
=|10568,10569
=|10569,10570
=|10570,10571
=|10571,10572
=|10572,10573
=|10573,10574
=|10574,10575
=|10575,10576
<EOL>|10576,10577
1|10577,10578
.|10578,10579
Patient|10580,10587
was|10588,10591
discharged|10592,10602
on|10603,10605
Amiodarone|10606,10616
200|10617,10620
mg|10621,10623
po|10624,10626
twice|10627,10632
daily|10633,10638
<EOL>|10639,10640
for|10640,10643
one|10644,10647
week|10648,10652
until|10653,10658
_|10659,10660
_|10660,10661
_|10661,10662
and|10663,10666
then|10667,10671
200mg|10672,10677
po|10678,10680
daily|10681,10686
thereafter|10687,10697
<EOL>|10698,10699
until|10699,10704
her|10705,10708
EP|10709,10711
appointment|10712,10723
with|10724,10728
Dr.|10729,10732
_|10733,10734
_|10734,10735
_|10735,10736
in|10737,10739
approximately|10740,10753
2|10754,10755
months|10756,10762
.|10762,10763
<EOL>|10763,10764
2.|10764,10766
Pt|10767,10769
was|10770,10773
discharged|10774,10784
on|10785,10787
Rivaroxaban|10788,10799
20|10800,10802
mg|10803,10805
qpm|10806,10809
with|10810,10814
dinner|10815,10821
<EOL>|10821,10822
3.|10822,10824
Pt|10825,10827
discharged|10828,10838
with|10839,10843
outpatient|10844,10854
_|10855,10856
_|10856,10857
_|10857,10858
of|10859,10861
Hearts|10862,10868
monitor|10869,10876
with|10877,10881
<EOL>|10882,10883
results|10883,10890
to|10891,10893
be|10894,10896
interpreted|10897,10908
by|10909,10911
Cardiologist|10912,10924
.|10924,10925
<EOL>|10925,10926
4.|10926,10928
She|10929,10932
presented|10933,10942
with|10943,10947
chest|10948,10953
pain|10954,10958
but|10959,10962
did|10963,10966
not|10967,10970
have|10971,10975
elevated|10976,10984
<EOL>|10985,10986
biomarkers|10986,10996
or|10997,10999
EKG|11000,11003
changes|11004,11011
concerning|11012,11022
for|11023,11026
myocardial|11027,11037
damage|11038,11044
.|11044,11045
<EOL>|11046,11047
Moreover|11047,11055
,|11055,11056
pt|11057,11059
remained|11060,11068
asymptomatic|11069,11081
during|11082,11088
periods|11089,11096
of|11097,11099
<EOL>|11100,11101
supraventricular|11101,11117
tachycardia|11118,11129
while|11130,11135
she|11136,11139
was|11140,11143
hospitalized|11144,11156
.|11156,11157
Patient|11158,11165
<EOL>|11166,11167
may|11167,11170
benefit|11171,11178
from|11179,11183
outpatient|11184,11194
stress|11195,11201
test|11202,11206
if|11207,11209
such|11210,11214
symptoms|11215,11223
return|11224,11230
.|11230,11231
<EOL>|11231,11232
5.|11232,11234
On|11235,11237
day|11238,11241
of|11242,11244
discharge|11245,11254
,|11254,11255
pt|11256,11258
had|11259,11262
significant|11263,11274
R|11275,11276
eye|11277,11280
pain|11281,11285
and|11286,11289
<EOL>|11290,11291
redness|11291,11298
,|11298,11299
was|11300,11303
evaluated|11304,11313
by|11314,11316
Optholmology|11317,11329
,|11329,11330
who|11331,11334
felt|11335,11339
that|11340,11344
it|11345,11347
was|11348,11351
<EOL>|11352,11353
just|11353,11357
dry|11358,11361
eyes|11362,11366
,|11366,11367
treated|11368,11375
with|11376,11380
erythromycin|11381,11393
drops|11394,11399
and|11400,11403
artifiical|11404,11414
<EOL>|11415,11416
tears|11416,11421
.|11421,11422
Patient|11423,11430
already|11431,11438
has|11439,11442
appt|11443,11447
w|11448,11449
/|11449,11450
Opthamology|11451,11462
in|11463,11465
5|11466,11467
days|11468,11472
which|11473,11478
<EOL>|11479,11480
she|11480,11483
will|11484,11488
need|11489,11493
to|11494,11496
attend|11497,11503
.|11503,11504
<EOL>|11504,11505
<EOL>|11505,11506
Full|11506,11510
Code|11511,11515
<EOL>|11515,11516
Contact|11516,11523
:|11523,11524
CONTACT|11525,11532
:|11532,11533
_|11534,11535
_|11535,11536
_|11536,11537
(|11538,11539
husband|11539,11546
)|11546,11547
_|11548,11549
_|11549,11550
_|11550,11551
_|11552,11553
_|11553,11554
_|11554,11555
<EOL>|11556,11557
(|11557,11558
daughter|11558,11566
)|11566,11567
_|11568,11569
_|11569,11570
_|11570,11571
<EOL>|11572,11573
<EOL>|11573,11574
<EOL>|11575,11576
Medications|11576,11587
on|11588,11590
Admission|11591,11600
:|11600,11601
<EOL>|11601,11602
The|11602,11605
Preadmission|11606,11618
Medication|11619,11629
list|11630,11634
is|11635,11637
accurate|11638,11646
and|11647,11650
complete|11651,11659
.|11659,11660
<EOL>|11660,11661
1.|11661,11663
Acetaminophen|11664,11677
325|11678,11681
mg|11682,11684
PO|11685,11687
Q4H|11688,11691
:|11691,11692
PRN|11692,11695
pain|11696,11700
<EOL>|11701,11702
2.|11702,11704
Albuterol|11705,11714
0.083|11715,11720
%|11720,11721
Neb|11722,11725
Soln|11726,11730
1|11731,11732
NEB|11733,11736
IH|11737,11739
Q6H|11740,11743
:|11743,11744
PRN|11744,11747
shortness|11748,11757
of|11758,11760
<EOL>|11761,11762
breath|11762,11768
<EOL>|11769,11770
3.|11770,11772
Aspirin|11773,11780
81|11781,11783
mg|11784,11786
PO|11787,11789
DAILY|11790,11795
<EOL>|11796,11797
4.|11797,11799
Atorvastatin|11800,11812
10|11813,11815
mg|11816,11818
PO|11819,11821
QPM|11822,11825
<EOL>|11826,11827
5.|11827,11829
Clopidogrel|11830,11841
75|11842,11844
mg|11845,11847
PO|11848,11850
DAILY|11851,11856
<EOL>|11857,11858
6.|11858,11860
Diltiazem|11861,11870
Extended|11871,11879
-|11879,11880
Release|11880,11887
180|11888,11891
mg|11892,11894
PO|11895,11897
DAILY|11898,11903
<EOL>|11904,11905
7.|11905,11907
Fluticasone|11908,11919
Propionate|11920,11930
NASAL|11931,11936
2|11937,11938
SPRY|11939,11943
NU|11944,11946
DAILY|11947,11952
:|11952,11953
PRN|11953,11956
nasal|11957,11962
<EOL>|11963,11964
congestion|11964,11974
<EOL>|11975,11976
8.|11976,11978
Fluticasone|11979,11990
-|11990,11991
Salmeterol|11991,12001
Diskus|12002,12008
(|12009,12010
250|12010,12013
/|12013,12014
50|12014,12016
)|12016,12017
1|12019,12020
INH|12021,12024
IH|12025,12027
BID|12028,12031
<EOL>|12032,12033
9.|12033,12035
Hydrochlorothiazide|12036,12055
50|12056,12058
mg|12059,12061
PO|12062,12064
DAILY|12065,12070
<EOL>|12071,12072
10.|12072,12075
Isosorbide|12076,12086
Mononitrate|12087,12098
(|12099,12100
Extended|12100,12108
Release|12109,12116
)|12116,12117
120|12118,12121
mg|12122,12124
PO|12125,12127
DAILY|12128,12133
<EOL>|12134,12135
11.|12135,12138
Latanoprost|12139,12150
0.005|12151,12156
%|12156,12157
Ophth|12158,12163
.|12163,12164
Soln.|12165,12170
1|12171,12172
DROP|12173,12177
LEFT|12178,12182
EYE|12183,12186
HS|12187,12189
<EOL>|12190,12191
12.|12191,12194
Lorazepam|12195,12204
0.5|12205,12208
mg|12209,12211
PO|12212,12214
QHS|12215,12218
:|12218,12219
PRN|12219,12222
insomnia|12223,12231
<EOL>|12232,12233
13.|12233,12236
Multivitamins|12237,12250
W|12251,12252
/|12252,12253
minerals|12253,12261
1|12262,12263
TAB|12264,12267
PO|12268,12270
DAILY|12271,12276
<EOL>|12277,12278
14.|12278,12281
Ranitidine|12282,12292
150|12293,12296
mg|12297,12299
PO|12300,12302
BID|12303,12306
<EOL>|12307,12308
15.|12308,12311
TraMADOL|12312,12320
(|12321,12322
Ultram|12322,12328
)|12328,12329
50|12330,12332
mg|12333,12335
PO|12336,12338
Q6H|12339,12342
:|12342,12343
PRN|12343,12346
pain|12347,12351
<EOL>|12352,12353
16|12353,12355
.|12355,12356
Theophylline|12357,12369
ER|12370,12372
300|12373,12376
mg|12377,12379
PO|12380,12382
BID|12383,12386
<EOL>|12387,12388
17.|12388,12391
Tiotropium|12392,12402
Bromide|12403,12410
1|12411,12412
CAP|12413,12416
IH|12417,12419
DAILY|12420,12425
<EOL>|12426,12427
18.|12427,12430
Guaifenesin|12431,12442
-|12442,12443
CODEINE|12443,12450
Phosphate|12451,12460
5|12461,12462
mL|12463,12465
PO|12466,12468
Q6H|12469,12472
:|12472,12473
PRN|12473,12476
cough|12477,12482
<EOL>|12483,12484
19.|12484,12487
cod|12488,12491
liver|12492,12497
oil|12498,12501
1,250|12502,12507
-|12507,12508
135|12508,12511
unit|12512,12516
oral|12517,12521
BID|12522,12525
<EOL>|12526,12527
20|12527,12529
.|12529,12530
Calcarb|12531,12538
600|12539,12542
With|12543,12547
Vitamin|12548,12555
D|12556,12557
(|12558,12559
calcium|12559,12566
carbonate|12567,12576
-|12576,12577
vitamin|12577,12584
D3|12585,12587
)|12587,12588
<EOL>|12589,12590
315|12590,12593
/|12593,12594
200|12594,12597
mg|12598,12600
oral|12601,12605
daily|12606,12611
<EOL>|12612,12613
<EOL>|12613,12614
<EOL>|12615,12616
Discharge|12616,12625
Medications|12626,12637
:|12637,12638
<EOL>|12638,12639
1.|12639,12641
Amiodarone|12642,12652
200|12653,12656
mg|12657,12659
PO|12660,12662
BID|12663,12666
<EOL>|12667,12668
RX|12668,12670
*|12671,12672
amiodarone|12672,12682
200|12683,12686
mg|12687,12689
1|12690,12691
tablet|12692,12698
(|12698,12699
s|12699,12700
)|12700,12701
by|12702,12704
mouth|12705,12710
twice|12711,12716
a|12717,12718
day|12719,12722
Disp|12723,12727
#|12728,12729
*|12729,12730
60|12730,12732
<EOL>|12733,12734
Tablet|12734,12740
Refills|12741,12748
:|12748,12749
*|12749,12750
1|12750,12751
<EOL>|12751,12752
2.|12752,12754
Rivaroxaban|12755,12766
20|12767,12769
mg|12770,12772
PO|12773,12775
DINNER|12776,12782
<EOL>|12783,12784
RX|12784,12786
*|12787,12788
rivaroxaban|12788,12799
[|12800,12801
Xarelto|12801,12808
]|12808,12809
20|12810,12812
mg|12813,12815
1|12816,12817
tablet|12818,12824
(|12824,12825
s|12825,12826
)|12826,12827
by|12828,12830
mouth|12831,12836
qpm|12837,12840
Disp|12841,12845
<EOL>|12846,12847
#|12847,12848
*|12848,12849
30|12849,12851
Tablet|12852,12858
Refills|12859,12866
:|12866,12867
*|12867,12868
1|12868,12869
<EOL>|12869,12870
3.|12870,12872
Acetaminophen|12873,12886
325|12887,12890
mg|12891,12893
PO|12894,12896
Q4H|12897,12900
:|12900,12901
PRN|12901,12904
pain|12905,12909
<EOL>|12910,12911
4.|12911,12913
Albuterol|12914,12923
0.083|12924,12929
%|12929,12930
Neb|12931,12934
Soln|12935,12939
1|12940,12941
NEB|12942,12945
IH|12946,12948
Q6H|12949,12952
:|12952,12953
PRN|12953,12956
shortness|12957,12966
of|12967,12969
<EOL>|12970,12971
breath|12971,12977
<EOL>|12978,12979
5.|12979,12981
Aspirin|12982,12989
81|12990,12992
mg|12993,12995
PO|12996,12998
DAILY|12999,13004
<EOL>|13005,13006
6.|13006,13008
Atorvastatin|13009,13021
10|13022,13024
mg|13025,13027
PO|13028,13030
QPM|13031,13034
<EOL>|13035,13036
7.|13036,13038
Diltiazem|13039,13048
Extended|13049,13057
-|13057,13058
Release|13058,13065
180|13066,13069
mg|13070,13072
PO|13073,13075
DAILY|13076,13081
<EOL>|13082,13083
8.|13083,13085
Fluticasone|13086,13097
Propionate|13098,13108
NASAL|13109,13114
2|13115,13116
SPRY|13117,13121
NU|13122,13124
DAILY|13125,13130
:|13130,13131
PRN|13131,13134
nasal|13135,13140
<EOL>|13141,13142
congestion|13142,13152
<EOL>|13153,13154
9.|13154,13156
Fluticasone|13157,13168
-|13168,13169
Salmeterol|13169,13179
Diskus|13180,13186
(|13187,13188
250|13188,13191
/|13191,13192
50|13192,13194
)|13194,13195
1|13197,13198
INH|13199,13202
IH|13203,13205
BID|13206,13209
<EOL>|13210,13211
10.|13211,13214
Guaifenesin|13215,13226
-|13226,13227
CODEINE|13227,13234
Phosphate|13235,13244
5|13245,13246
mL|13247,13249
PO|13250,13252
Q6H|13253,13256
:|13256,13257
PRN|13257,13260
cough|13261,13266
<EOL>|13267,13268
11|13268,13270
.|13270,13271
Hydrochlorothiazide|13272,13291
50|13292,13294
mg|13295,13297
PO|13298,13300
DAILY|13301,13306
<EOL>|13307,13308
12.|13308,13311
Isosorbide|13312,13322
Mononitrate|13323,13334
(|13335,13336
Extended|13336,13344
Release|13345,13352
)|13352,13353
120|13354,13357
mg|13358,13360
PO|13361,13363
DAILY|13364,13369
<EOL>|13370,13371
13.|13371,13374
Latanoprost|13375,13386
0.005|13387,13392
%|13392,13393
Ophth|13394,13399
.|13399,13400
Soln.|13401,13406
1|13407,13408
DROP|13409,13413
LEFT|13414,13418
EYE|13419,13422
HS|13423,13425
<EOL>|13426,13427
14.|13427,13430
Lorazepam|13431,13440
0.5|13441,13444
mg|13445,13447
PO|13448,13450
QHS|13451,13454
:|13454,13455
PRN|13455,13458
insomnia|13459,13467
<EOL>|13468,13469
15.|13469,13472
Multivitamins|13473,13486
W|13487,13488
/|13488,13489
minerals|13489,13497
1|13498,13499
TAB|13500,13503
PO|13504,13506
DAILY|13507,13512
<EOL>|13513,13514
16|13514,13516
.|13516,13517
Ranitidine|13518,13528
150|13529,13532
mg|13533,13535
PO|13536,13538
BID|13539,13542
<EOL>|13543,13544
17.|13544,13547
Theophylline|13548,13560
ER|13561,13563
300|13564,13567
mg|13568,13570
PO|13571,13573
BID|13574,13577
<EOL>|13578,13579
18.|13579,13582
Tiotropium|13583,13593
Bromide|13594,13601
1|13602,13603
CAP|13604,13607
IH|13608,13610
DAILY|13611,13616
<EOL>|13617,13618
19|13618,13620
.|13620,13621
TraMADOL|13622,13630
(|13631,13632
Ultram|13632,13638
)|13638,13639
50|13640,13642
mg|13643,13645
PO|13646,13648
Q6H|13649,13652
:|13652,13653
PRN|13653,13656
pain|13657,13661
<EOL>|13662,13663
20|13663,13665
.|13665,13666
Artificial|13667,13677
Tears|13678,13683
Preserv|13684,13691
.|13691,13692
Free|13693,13697
_|13698,13699
_|13699,13700
_|13700,13701
DROP|13702,13706
BOTH|13707,13711
EYES|13712,13716
PRN|13717,13720
eye|13721,13724
<EOL>|13725,13726
irritation|13726,13736
<EOL>|13737,13738
RX|13738,13740
*|13741,13742
dextran|13742,13749
70|13750,13752
-|13752,13753
hypromellose|13753,13765
[|13766,13767
Artificial|13767,13777
Tears|13778,13783
]|13783,13784
1|13786,13787
drop|13788,13792
OPTH|13793,13797
<EOL>|13798,13799
QID|13799,13802
:|13802,13803
prn|13803,13806
Refills|13807,13814
:|13814,13815
*|13815,13816
0|13816,13817
<EOL>|13817,13818
RX|13818,13820
*|13821,13822
dextran|13822,13829
70|13830,13832
-|13832,13833
hypromellose|13833,13845
[|13846,13847
Artificial|13847,13857
Tears|13858,13863
(|13864,13865
PF|13865,13867
)|13867,13868
]|13868,13869
_|13871,13872
_|13872,13873
_|13873,13874
drops|13875,13880
<EOL>|13881,13882
eye|13882,13885
as|13886,13888
needed|13889,13895
Disp|13896,13900
#|13901,13902
*|13902,13903
1|13903,13904
Package|13905,13912
Refills|13913,13920
:|13920,13921
*|13921,13922
1|13922,13923
<EOL>|13923,13924
21|13924,13926
.|13926,13927
Erythromycin|13928,13940
0.5|13941,13944
%|13944,13945
Ophth|13946,13951
Oint|13952,13956
0.5|13957,13960
in|13961,13963
RIGHT|13964,13969
EYE|13970,13973
TID|13974,13977
<EOL>|13978,13979
RX|13979,13981
*|13982,13983
erythromycin|13983,13995
5|13996,13997
mg|13998,14000
/|14000,14001
gram|14001,14005
(|14006,14007
0.5|14007,14010
%|14011,14012
)|14012,14013
0.5|14014,14017
(|14018,14019
One|14019,14022
half|14023,14027
)|14027,14028
inch|14029,14033
OPTH|14034,14038
<EOL>|14039,14040
TID|14040,14043
:|14043,14044
prn|14044,14047
Refills|14048,14055
:|14055,14056
*|14056,14057
0|14057,14058
<EOL>|14058,14059
22.|14059,14062
Calcarb|14063,14070
600|14071,14074
With|14075,14079
Vitamin|14080,14087
D|14088,14089
(|14090,14091
calcium|14091,14098
carbonate|14099,14108
-|14108,14109
vitamin|14109,14116
D3|14117,14119
)|14119,14120
<EOL>|14121,14122
315|14122,14125
/|14125,14126
200|14126,14129
mg|14130,14132
oral|14133,14137
daily|14138,14143
<EOL>|14144,14145
23.|14145,14148
cod|14149,14152
liver|14153,14158
oil|14159,14162
1,250|14163,14168
-|14168,14169
135|14169,14172
unit|14173,14177
oral|14178,14182
BID|14183,14186
<EOL>|14187,14188
<EOL>|14188,14189
<EOL>|14190,14191
Discharge|14191,14200
Disposition|14201,14212
:|14212,14213
<EOL>|14213,14214
Home|14214,14218
<EOL>|14218,14219
<EOL>|14220,14221
Discharge|14221,14230
Diagnosis|14231,14240
:|14240,14241
<EOL>|14241,14242
Rapid|14242,14247
Atrial|14248,14254
Fibrillation|14255,14267
/|14267,14268
Flutter|14268,14275
<EOL>|14275,14276
COPD|14276,14280
<EOL>|14280,14281
<EOL>|14281,14282
<EOL>|14283,14284
Mental|14305,14311
Status|14312,14318
:|14318,14319
Clear|14320,14325
and|14326,14329
coherent|14330,14338
.|14338,14339
<EOL>|14339,14340
Level|14340,14345
of|14346,14348
Consciousness|14349,14362
:|14362,14363
Alert|14364,14369
and|14370,14373
interactive|14374,14385
.|14385,14386
<EOL>|14386,14387
Activity|14387,14395
Status|14396,14402
:|14402,14403
Ambulatory|14404,14414
-|14415,14416
Independent|14417,14428
.|14428,14429
<EOL>|14429,14430
<EOL>|14430,14431
<EOL>|14432,14433
Dear|14457,14461
Ms.|14462,14465
_|14466,14467
_|14467,14468
_|14468,14469
,|14469,14470
<EOL>|14470,14471
<EOL>|14471,14472
You|14472,14475
were|14476,14480
admitted|14481,14489
to|14490,14492
_|14493,14494
_|14494,14495
_|14495,14496
due|14497,14500
to|14501,14503
concerning|14504,14514
chest|14515,14520
pain|14521,14525
symptoms|14526,14534
<EOL>|14535,14536
which|14536,14541
we|14542,14544
think|14545,14550
are|14551,14554
due|14555,14558
to|14559,14561
infrequent|14562,14572
bursts|14573,14579
of|14580,14582
a|14583,14584
rapid|14585,14590
heart|14591,14596
<EOL>|14597,14598
rate|14598,14602
.|14602,14603
Since|14604,14609
the|14610,14613
rapid|14614,14619
rate|14620,14624
makes|14625,14630
you|14631,14634
at|14635,14637
increased|14638,14647
risk|14648,14652
for|14653,14656
<EOL>|14657,14658
stroke|14658,14664
,|14664,14665
you|14666,14669
were|14670,14674
started|14675,14682
on|14683,14685
a|14686,14687
blood|14688,14693
thinning|14694,14702
medication|14703,14713
called|14714,14720
<EOL>|14721,14722
Rivaroxaban|14722,14733
which|14734,14739
you|14740,14743
will|14744,14748
need|14749,14753
to|14754,14756
take|14757,14761
every|14762,14767
day|14768,14771
.|14771,14772
Our|14773,14776
<EOL>|14777,14778
specialized|14778,14789
cardiologists|14790,14803
who|14804,14807
deal|14808,14812
specifically|14813,14825
with|14826,14830
the|14831,14834
<EOL>|14835,14836
electrical|14836,14846
rhythm|14847,14853
of|14854,14856
the|14857,14860
heart|14861,14866
evaluated|14867,14876
you|14877,14880
and|14881,14884
felt|14885,14889
that|14890,14894
you|14895,14898
<EOL>|14899,14900
would|14900,14905
benefit|14906,14913
from|14914,14918
a|14919,14920
medication|14921,14931
called|14932,14938
amiodarone|14939,14949
which|14950,14955
was|14956,14959
also|14960,14964
<EOL>|14965,14966
started|14966,14973
.|14973,14974
You|14975,14978
will|14979,14983
need|14984,14988
to|14989,14991
follow|14992,14998
up|14999,15001
with|15002,15006
them|15007,15011
in|15012,15014
their|15015,15020
clinic|15021,15027
<EOL>|15028,15029
regarding|15029,15038
this|15039,15043
abnormal|15044,15052
rhythm|15053,15059
.|15059,15060
In|15061,15063
the|15064,15067
meantime|15068,15076
,|15076,15077
you|15078,15081
were|15082,15086
<EOL>|15087,15088
outfitted|15088,15097
with|15098,15102
a|15103,15104
Holter|15105,15111
monitor|15112,15119
to|15120,15122
record|15123,15129
your|15130,15134
heart|15135,15140
rate|15141,15145
at|15146,15148
<EOL>|15149,15150
home|15150,15154
.|15154,15155
It|15156,15158
is|15159,15161
very|15162,15166
important|15167,15176
that|15177,15181
you|15182,15185
follow|15186,15192
up|15193,15195
with|15196,15200
Dr.|15201,15204
_|15205,15206
_|15206,15207
_|15207,15208
<EOL>|15209,15210
your|15210,15214
cardiologist|15215,15227
.|15227,15228
<EOL>|15228,15229
<EOL>|15229,15230
We|15230,15232
wish|15233,15237
you|15238,15241
all|15242,15245
the|15246,15249
best|15250,15254
,|15254,15255
<EOL>|15255,15256
<EOL>|15256,15257
Sincerely|15257,15266
,|15266,15267
<EOL>|15267,15268
Your|15268,15272
care|15273,15277
team|15278,15282
at|15283,15285
_|15286,15287
_|15287,15288
_|15288,15289
<EOL>|15289,15290
<EOL>|15291,15292
Followup|15292,15300
Instructions|15301,15313
:|15313,15314
<EOL>|15314,15315
_|15315,15316
_|15316,15317
_|15317,15318
<EOL>|15318,15319

