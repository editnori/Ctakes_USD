 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|176,183|false|false|false|C0591292|Corgard|Corgard
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|176,183|false|false|false|C0591292|Corgard|Corgard
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|186,193|false|false|false|C0728763|Vasotec|Vasotec
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|186,193|false|false|false|C0728763|Vasotec|Vasotec
Event|Event|SIMPLE_SEGMENT|196,205|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|196,205|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|213,228|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|219,228|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|219,228|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|219,228|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|230,233|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|230,239|false|true|false|C0235886|Leg edema|leg edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|234,239|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|234,239|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|234,239|false|false|false|C0013604|Edema|edema
Finding|Classification|SIMPLE_SEGMENT|242,247|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|248,256|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|248,256|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|260,278|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|269,278|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|269,278|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|269,278|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|269,278|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|269,278|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|288,295|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|288,295|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|288,295|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|288,295|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|288,298|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|288,314|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|288,314|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|299,306|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|299,306|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|299,314|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|307,314|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|316,323|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|316,326|false|false|false|C0262926|Medical History|HISTORY OF
Finding|Idea or Concept|SIMPLE_SEGMENT|327,337|true|false|false|C0449450|Presentation|PRESENTING
Event|Event|SIMPLE_SEGMENT|338,345|false|false|false|||ILLNESS
Finding|Sign or Symptom|SIMPLE_SEGMENT|338,345|false|false|false|C0221423|Illness (finding)|ILLNESS
Finding|Idea or Concept|SIMPLE_SEGMENT|368,372|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|368,372|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|373,376|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|392,399|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|392,399|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|392,399|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|392,399|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|392,402|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|403,406|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|403,406|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|403,406|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|403,406|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|403,406|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|403,406|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|403,406|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|403,406|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|416,420|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|416,420|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|429,432|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|429,432|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|429,432|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|429,432|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|429,432|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|429,432|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|438,447|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|438,447|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|438,447|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|448,451|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|448,451|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|453,457|false|false|false|C0004238|Atrial Fibrillation|AFib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|453,457|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Event|Event|SIMPLE_SEGMENT|462,477|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|462,477|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|462,477|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|462,477|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|496,504|false|false|false|||presents
Finding|Intellectual Product|SIMPLE_SEGMENT|510,516|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|510,525|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|517,525|false|false|false|||overload
Finding|Finding|SIMPLE_SEGMENT|531,534|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|531,534|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|535,540|false|false|false|||found
Finding|Finding|SIMPLE_SEGMENT|535,540|false|false|false|C0150312|Present|found
Event|Event|SIMPLE_SEGMENT|544,552|false|false|false|||dilation
Finding|Finding|SIMPLE_SEGMENT|544,552|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Finding|Pathologic Function|SIMPLE_SEGMENT|544,552|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|544,552|false|false|false|C1322279|Dilate procedure|dilation
Finding|Idea or Concept|SIMPLE_SEGMENT|556,562|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|563,577|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|563,577|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Body Substance|SIMPLE_SEGMENT|582,589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|582,589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|582,589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|590,597|false|false|false|||reports
Finding|Mental Process|SIMPLE_SEGMENT|630,637|false|false|false|C1527305|Feelings|feeling
Finding|Sign or Symptom|SIMPLE_SEGMENT|630,645|false|false|false|C0849963|Feeling nervous|feeling nervous
Event|Event|SIMPLE_SEGMENT|638,645|false|false|false|||nervous
Finding|Functional Concept|SIMPLE_SEGMENT|638,645|false|false|false|C0027769;C0599851|Nervous - anatomy qualifier;Nervousness|nervous
Finding|Sign or Symptom|SIMPLE_SEGMENT|638,645|false|false|false|C0027769;C0599851|Nervous - anatomy qualifier;Nervousness|nervous
Event|Event|SIMPLE_SEGMENT|651,658|false|false|false|||jittery
Finding|Mental Process|SIMPLE_SEGMENT|651,658|false|false|false|C2987186|Jittery|jittery
Event|Event|SIMPLE_SEGMENT|668,676|false|false|false|||endorses
Attribute|Clinical Attribute|SIMPLE_SEGMENT|677,683|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|677,683|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|677,683|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|677,683|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|677,683|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|677,688|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Finding|Intellectual Product|SIMPLE_SEGMENT|677,688|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Event|Event|SIMPLE_SEGMENT|684,688|false|false|false|||gain
Finding|Finding|SIMPLE_SEGMENT|694,697|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|694,697|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|694,703|false|false|false|C0746890|new onset|new onset
Anatomy|Body Location or Region|SIMPLE_SEGMENT|704,709|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|704,709|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|711,720|false|false|false|C0015385|Limb structure|extremity
Finding|Sign or Symptom|SIMPLE_SEGMENT|711,729|false|false|false|C0158369|Swelling of limb|extremity swelling
Event|Event|SIMPLE_SEGMENT|721,729|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|721,729|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|721,729|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|746,751|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|746,751|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|746,756|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|746,756|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|752,756|true|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|752,756|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|752,756|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|752,756|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|758,770|true|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|758,770|true|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|773,782|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|773,782|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|773,782|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|787,790|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|787,790|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|787,790|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|SIMPLE_SEGMENT|811,817|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|811,817|true|false|false|C0015967|Fever|fevers
Drug|Organic Chemical|SIMPLE_SEGMENT|819,824|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|819,824|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|819,824|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|819,824|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|826,832|true|false|false|||recent
Event|Event|SIMPLE_SEGMENT|834,840|true|false|false|||travel
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|834,840|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|SIMPLE_SEGMENT|834,840|true|false|false|C1555670|travel charge|travel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|842,852|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|842,852|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|842,852|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Individual Behavior|SIMPLE_SEGMENT|842,867|false|false|false|C3489773|Medication Compliance|medication non compliance
Event|Event|SIMPLE_SEGMENT|857,867|false|false|false|||compliance
Finding|Finding|SIMPLE_SEGMENT|857,867|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|SIMPLE_SEGMENT|857,867|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|SIMPLE_SEGMENT|857,867|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Event|Event|SIMPLE_SEGMENT|869,878|false|false|false|||increased
Drug|Food|SIMPLE_SEGMENT|879,889|false|false|false|C0453862|Salty food|salty food
Drug|Food|SIMPLE_SEGMENT|885,889|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|885,889|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|885,889|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Finding|Organism Function|SIMPLE_SEGMENT|885,896|false|false|false|C0013470|Eating|food intake
Event|Event|SIMPLE_SEGMENT|890,896|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|890,896|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|890,896|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|919,926|true|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|919,926|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|919,926|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|919,938|true|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|SIMPLE_SEGMENT|930,938|true|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|930,938|true|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|943,948|true|false|false|||rides
Event|Event|SIMPLE_SEGMENT|951,956|false|false|false|||miles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|957,960|false|false|false|C0449201|PER (body structure)|per
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|957,960|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|per
Finding|Functional Concept|SIMPLE_SEGMENT|957,960|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Finding|Gene or Genome|SIMPLE_SEGMENT|957,960|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Finding|Intellectual Product|SIMPLE_SEGMENT|957,960|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|per
Finding|Idea or Concept|SIMPLE_SEGMENT|962,965|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|962,965|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|971,981|false|false|false|C3839460||stationary
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|971,986|false|false|false|C2712863|Stationary bike|stationary bike
Event|Event|SIMPLE_SEGMENT|982,986|false|false|false|||bike
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|982,986|false|false|false|C0005377;C1425261|BMP2K gene;Bicycling (recreational activity)|bike
Finding|Gene or Genome|SIMPLE_SEGMENT|982,986|false|false|false|C0005377;C1425261|BMP2K gene;Bicycling (recreational activity)|bike
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1009,1015|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|1009,1015|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|1009,1015|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|1009,1015|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|1009,1015|false|false|false|C1305866|Weighing patient|weight
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1009,1023|false|false|false|C0043095|Weight Lifting|weight lifting
Event|Activity|SIMPLE_SEGMENT|1016,1023|false|false|false|C0206244|Lifting|lifting
Event|Event|SIMPLE_SEGMENT|1016,1023|false|false|false|||lifting
Event|Event|SIMPLE_SEGMENT|1031,1040|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|1062,1072|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|1062,1072|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1062,1072|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|1090,1093|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1090,1093|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|1099,1105|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|1106,1109|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1106,1109|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|1113,1121|false|false|false|||dilation
Finding|Finding|SIMPLE_SEGMENT|1113,1121|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Finding|Pathologic Function|SIMPLE_SEGMENT|1113,1121|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1113,1121|false|false|false|C1322279|Dilate procedure|dilation
Event|Event|SIMPLE_SEGMENT|1130,1138|false|false|false|||referred
Event|Event|SIMPLE_SEGMENT|1151,1153|false|false|false|||ED
Event|Event|SIMPLE_SEGMENT|1166,1176|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|1166,1176|false|true|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1166,1176|false|true|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|1182,1189|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|1182,1189|false|false|true|C2699424|Concern|concern
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1194,1203|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1194,1203|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1194,1203|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|1205,1213|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|1205,1213|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|1205,1213|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Idea or Concept|SIMPLE_SEGMENT|1231,1238|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1239,1245|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1255,1258|false|false|false|||T98
Event|Event|SIMPLE_SEGMENT|1297,1301|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1297,1301|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1297,1301|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|1320,1343|false|false|false|C2237594|bilateral pitting edema|bilateral pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|1330,1337|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|1330,1343|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1338,1343|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1338,1343|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1338,1343|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1347,1352|false|false|false|C0022742|Knee|knees
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1354,1358|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1360,1367|false|false|false|||notable
Finding|Intellectual Product|SIMPLE_SEGMENT|1372,1376|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1377,1389|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|SIMPLE_SEGMENT|1377,1389|false|false|false|||hyponatremia
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1399,1402|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1399,1402|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|1399,1402|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|1399,1402|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|1399,1402|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|1399,1402|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|1399,1402|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1399,1402|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1403,1406|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1403,1406|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1403,1406|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1403,1406|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|1403,1406|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|1403,1406|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|1403,1406|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Event|Event|SIMPLE_SEGMENT|1414,1422|false|false|false|||elevated
Anatomy|Cell|SIMPLE_SEGMENT|1434,1437|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1441,1444|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1441,1444|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|1441,1444|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1441,1444|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1441,1444|false|false|false|C0019029|Hemoglobin concentration|Hgb
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1451,1454|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|1451,1454|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1451,1454|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1451,1454|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1460,1466|false|false|false|C0060323|Fibrin fragment D|DDimer
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1460,1466|false|false|false|C0060323|Fibrin fragment D|DDimer
Event|Event|SIMPLE_SEGMENT|1460,1466|false|false|false|||DDimer
Event|Event|SIMPLE_SEGMENT|1477,1489|false|false|false|||unremarkable
Event|Event|SIMPLE_SEGMENT|1494,1497|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1494,1497|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|1503,1507|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|1508,1520|false|false|false|||cardiomegaly
Finding|Finding|SIMPLE_SEGMENT|1508,1520|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|SIMPLE_SEGMENT|1528,1536|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|1528,1536|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1528,1539|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1540,1553|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|1540,1553|true|false|false|||consolidation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1558,1567|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1558,1567|true|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1558,1567|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|1558,1573|true|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1568,1573|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1568,1573|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1568,1573|true|false|false|C0013604|Edema|edema
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1575,1578|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|1575,1578|true|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|1575,1578|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1575,1578|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|SIMPLE_SEGMENT|1583,1591|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1583,1591|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1583,1591|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1583,1591|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1583,1595|false|false|false|C0205160|Negative|negative for
Event|Event|SIMPLE_SEGMENT|1600,1606|true|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1607,1613|true|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|1607,1613|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1607,1613|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1615,1624|true|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|SIMPLE_SEGMENT|1615,1624|true|false|false|||emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|1615,1624|true|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Finding|Finding|SIMPLE_SEGMENT|1629,1636|false|false|false|C0700124|Dilated|dilated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1629,1653|false|false|false|C0428851|Dilatation of pulmonary artery (disorder)|dilated pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1637,1646|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1637,1646|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1637,1646|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1637,1653|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1647,1653|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|1647,1653|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Body Substance|SIMPLE_SEGMENT|1658,1665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1658,1665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1658,1665|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|1666,1674|false|false|false|||received
Drug|Organic Chemical|SIMPLE_SEGMENT|1684,1689|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1684,1689|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|SIMPLE_SEGMENT|1695,1706|false|false|false|C0750502|Significant|significant
Finding|Body Substance|SIMPLE_SEGMENT|1707,1712|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|1707,1712|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|1707,1712|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1707,1719|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1707,1719|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|SIMPLE_SEGMENT|1713,1719|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|1713,1719|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|1713,1719|false|false|false|C3251815|Measurement of fluid output|output
Finding|Body Substance|SIMPLE_SEGMENT|1725,1732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1725,1732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1725,1732|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1741,1745|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1746,1754|false|false|false|||admitted
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1762,1767|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1762,1767|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1762,1767|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1762,1775|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|1768,1775|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|1768,1775|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|1768,1775|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|1768,1775|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Occupational Activity|SIMPLE_SEGMENT|1776,1783|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|1776,1783|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Finding|Intellectual Product|SIMPLE_SEGMENT|1789,1794|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1789,1808|false|false|false|C0264714|Acute heart failure|acute heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1795,1800|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1795,1800|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1795,1800|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1795,1808|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|1801,1808|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|1801,1808|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|1801,1808|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|1801,1808|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|1809,1821|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|1809,1821|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|SIMPLE_SEGMENT|1834,1840|false|false|false|||workup
Event|Event|SIMPLE_SEGMENT|1848,1856|false|false|false|||dilation
Finding|Finding|SIMPLE_SEGMENT|1848,1856|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Finding|Pathologic Function|SIMPLE_SEGMENT|1848,1856|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1848,1856|false|false|false|C1322279|Dilate procedure|dilation
Event|Event|SIMPLE_SEGMENT|1861,1867|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|1871,1879|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1871,1879|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1871,1879|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1871,1879|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1881,1889|false|false|false|||Afebrile
Finding|Finding|SIMPLE_SEGMENT|1881,1889|false|false|false|C0277797|Apyrexial|Afebrile
Event|Event|SIMPLE_SEGMENT|1931,1937|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|1931,1937|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|1931,1937|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|1931,1940|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1931,1948|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|1931,1948|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|1941,1948|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|1941,1948|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|1953,1959|true|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1970,1977|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1970,1977|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1970,1977|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1970,1977|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1970,1980|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1981,1987|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1981,1987|true|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1981,1987|true|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1990,1993|true|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|SIMPLE_SEGMENT|1990,1993|true|false|false|||TIA
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1995,1999|false|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1995,2017|false|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2000,2006|false|false|false|C0042449|Veins|venous
Finding|Finding|SIMPLE_SEGMENT|2000,2017|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2000,2017|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|SIMPLE_SEGMENT|2007,2017|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2007,2017|false|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2019,2028|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2019,2028|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|2019,2028|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|2019,2037|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|SIMPLE_SEGMENT|2029,2037|false|false|false|||embolism
Finding|Finding|SIMPLE_SEGMENT|2029,2037|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|2029,2037|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|SIMPLE_SEGMENT|2039,2047|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|2039,2047|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|2056,2060|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|2056,2060|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|2056,2060|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|2064,2071|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|2064,2071|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2064,2071|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2064,2071|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2064,2071|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|2073,2081|false|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2073,2081|false|false|false|C0231528|Myalgia|myalgias
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2083,2088|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|SIMPLE_SEGMENT|2083,2088|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|SIMPLE_SEGMENT|2083,2088|false|false|false|C0575044|Joint problem|joint
Finding|Sign or Symptom|SIMPLE_SEGMENT|2083,2094|false|false|false|C0003862|Arthralgia|joint pains
Event|Event|SIMPLE_SEGMENT|2089,2094|false|false|false|||pains
Finding|Sign or Symptom|SIMPLE_SEGMENT|2089,2094|false|false|false|C0030193|Pain|pains
Drug|Organic Chemical|SIMPLE_SEGMENT|2096,2101|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2096,2101|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2096,2101|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2096,2101|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|2103,2113|false|false|false|||hemoptysis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2103,2113|false|false|false|C0019079|Hemoptysis|hemoptysis
Event|Event|SIMPLE_SEGMENT|2115,2120|false|false|false|||black
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2122,2128|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|2122,2128|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|2122,2128|false|false|false|C0015733|Feces|stools
Finding|Finding|SIMPLE_SEGMENT|2132,2135|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|2132,2135|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Sign or Symptom|SIMPLE_SEGMENT|2132,2142|false|false|false|C0278012|Red stools|red stools
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2136,2142|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|2136,2142|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|2136,2142|false|false|false|C0015733|Feces|stools
Event|Event|SIMPLE_SEGMENT|2147,2153|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|2161,2167|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|2161,2167|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|2169,2175|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2169,2175|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|2179,2185|true|false|false|||rigors
Finding|Sign or Symptom|SIMPLE_SEGMENT|2179,2185|true|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Event|Event|SIMPLE_SEGMENT|2191,2197|false|false|false|||denies
Finding|Sign or Symptom|SIMPLE_SEGMENT|2198,2208|true|false|false|C0239313|exercise induced|exertional
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2209,2216|true|false|false|C0006497|Buttocks|buttock
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2220,2224|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2220,2224|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|SIMPLE_SEGMENT|2220,2229|true|false|false|C0236040|Pain in calf|calf pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2225,2229|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2225,2229|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2225,2229|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2225,2229|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2249,2255|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|2249,2255|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|2249,2255|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|2249,2258|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2249,2266|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2249,2266|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|2259,2266|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2259,2266|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|2272,2280|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|2272,2280|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2272,2280|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2272,2280|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2287,2294|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2287,2294|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|SIMPLE_SEGMENT|2295,2301|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|2295,2301|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|2295,2301|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|2295,2304|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2295,2312|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2295,2312|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|2305,2312|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2305,2312|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|2316,2323|false|false|false|||notable
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2328,2335|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|SIMPLE_SEGMENT|2328,2335|false|false|false|||absence
Finding|Functional Concept|SIMPLE_SEGMENT|2328,2335|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|SIMPLE_SEGMENT|2328,2338|false|false|false|C0332197|Absent|absence of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2339,2344|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2339,2344|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2339,2349|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2339,2349|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2345,2349|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2345,2349|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2345,2349|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2345,2349|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2352,2380|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|paroxysmal nocturnal dyspnea
Event|Event|SIMPLE_SEGMENT|2373,2380|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|2373,2380|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2373,2380|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|2382,2391|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|2382,2391|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2382,2391|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|SIMPLE_SEGMENT|2393,2405|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|2393,2405|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|2407,2414|false|false|false|||syncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|2407,2414|false|false|false|C0039070|Syncope|syncope
Event|Event|SIMPLE_SEGMENT|2419,2429|false|false|false|||presyncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|2419,2429|false|false|false|C0700200|Presyncope|presyncope
Finding|Finding|SIMPLE_SEGMENT|2438,2458|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2443,2450|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2443,2450|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2443,2450|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2443,2450|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2443,2450|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2443,2458|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2451,2458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2451,2458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2451,2458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2460,2480|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2465,2472|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2465,2472|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2465,2472|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2465,2472|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2465,2472|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2465,2480|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2473,2480|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2473,2480|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2473,2480|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2492,2500|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Finding|Intellectual Product|SIMPLE_SEGMENT|2492,2500|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2501,2508|false|false|false|C0007272|Carotid Arteries|CAROTID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2501,2516|false|false|false|C0741975|carotid disease|CAROTID DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2509,2516|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|2509,2516|false|false|false|||DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2518,2542|false|false|false|C0018802|Congestive heart failure|CONGESTIVE HEART FAILURE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2529,2534|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2529,2534|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|2529,2534|false|false|false|C0795691|HEART PROBLEM|HEART
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2529,2542|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|HEART FAILURE
Event|Event|SIMPLE_SEGMENT|2535,2542|false|false|false|||FAILURE
Finding|Functional Concept|SIMPLE_SEGMENT|2535,2542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|SIMPLE_SEGMENT|2535,2542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|SIMPLE_SEGMENT|2535,2542|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2544,2552|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2544,2559|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2544,2567|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2553,2559|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|SIMPLE_SEGMENT|2553,2559|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2553,2567|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2560,2567|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|2560,2567|false|false|false|||DISEASE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2569,2585|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2569,2592|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|SIMPLE_SEGMENT|2569,2592|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Event|Event|SIMPLE_SEGMENT|2586,2592|false|false|false|||REFLUX
Finding|Pathologic Function|SIMPLE_SEGMENT|2586,2592|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2594,2606|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|SIMPLE_SEGMENT|2594,2606|false|false|false|||HYPERTENSION
Finding|Finding|SIMPLE_SEGMENT|2608,2614|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Finding|Intellectual Product|SIMPLE_SEGMENT|2608,2614|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2615,2624|false|false|false|C0034067|Pulmonary Emphysema|EMPHYSEMA
Event|Event|SIMPLE_SEGMENT|2615,2624|false|false|false|||EMPHYSEMA
Finding|Pathologic Function|SIMPLE_SEGMENT|2615,2624|false|false|false|C0013990|Pathological accumulation of air in tissues|EMPHYSEMA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2626,2635|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2626,2635|false|false|false|C2707265||PULMONARY
Finding|Finding|SIMPLE_SEGMENT|2626,2635|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Pathologic Function|SIMPLE_SEGMENT|2626,2648|false|false|false|C0020542|Pulmonary Hypertension|PULMONARY HYPERTENSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2636,2648|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|SIMPLE_SEGMENT|2636,2648|false|false|false|||HYPERTENSION
Finding|Functional Concept|SIMPLE_SEGMENT|2650,2655|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2650,2669|false|false|false|C0225916|Structure of right branch of atrioventricular bundle|RIGHT BUNDLE BRANCH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2650,2675|false|false|false|C0085615|Right bundle branch block|RIGHT BUNDLE BRANCH BLOCK
Finding|Finding|SIMPLE_SEGMENT|2650,2675|false|false|false|C0344421||RIGHT BUNDLE BRANCH BLOCK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2656,2675|false|false|false|C0006384;C1879286|Bundle-Branch Block;Hereditary bundle branch system defect|BUNDLE BRANCH BLOCK
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2663,2669|false|false|false|C1881507|Macromolecular Branch|BRANCH
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2670,2675|false|false|false|C1706085|Block Dosage Form|BLOCK
Event|Event|SIMPLE_SEGMENT|2670,2675|false|false|false|||BLOCK
Finding|Body Substance|SIMPLE_SEGMENT|2670,2675|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Finding|SIMPLE_SEGMENT|2670,2675|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Functional Concept|SIMPLE_SEGMENT|2670,2675|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Pathologic Function|SIMPLE_SEGMENT|2677,2705|false|false|false|C1704272|Benign Prostatic Hyperplasia|BENIGN PROSTATIC HYPERTROPHY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2684,2693|false|false|false|C0033572|Prostate|PROSTATIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2684,2705|false|false|false|C1739363|Prostatic Hypertrophy|PROSTATIC HYPERTROPHY
Finding|Pathologic Function|SIMPLE_SEGMENT|2684,2705|false|false|false|C1704272;C2937421|Benign Prostatic Hyperplasia;Prostatic Hyperplasia|PROSTATIC HYPERTROPHY
Event|Event|SIMPLE_SEGMENT|2694,2705|false|false|false|||HYPERTROPHY
Finding|Pathologic Function|SIMPLE_SEGMENT|2694,2705|false|false|false|C0020564|Hypertrophy|HYPERTROPHY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2707,2721|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|SIMPLE_SEGMENT|2707,2721|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|SIMPLE_SEGMENT|2707,2721|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Event|Event|SIMPLE_SEGMENT|2723,2733|false|false|false|||PAROXYSMAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2723,2753|false|false|false|C0235480|Paroxysmal atrial fibrillation|PAROXYSMAL ATRIAL FIBRILLATION
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2734,2740|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2734,2753|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2734,2753|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2734,2753|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2741,2753|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|SIMPLE_SEGMENT|2741,2753|false|false|false|||FIBRILLATION
Finding|Finding|SIMPLE_SEGMENT|2777,2798|false|false|false|C0455610|History of surgery|Past Surgical History
Procedure|Health Care Activity|SIMPLE_SEGMENT|2782,2790|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2782,2790|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Finding|Finding|SIMPLE_SEGMENT|2782,2798|false|false|false|C0744961|history of prior surgery|Surgical History
Event|Event|SIMPLE_SEGMENT|2791,2798|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2791,2798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2791,2798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2791,2798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2800,2813|false|false|false|||CARDIOVERSION
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2800,2813|false|false|false|C0013778|Electric Countershock|CARDIOVERSION
Finding|Functional Concept|SIMPLE_SEGMENT|2819,2824|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2819,2835|false|false|false|C1261075|Structure of right lower lobe of lung|RIGHT LOWER LOBE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2825,2830|false|false|false|C1548802|Body Site Modifier - Lower|LOWER
Event|Activity|SIMPLE_SEGMENT|2825,2830|false|false|false|C2003888|Lower (action)|LOWER
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2825,2835|false|false|false|C0225758|Structure of lower lobe of lung|LOWER LOBE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2831,2835|false|false|false|C0796494|lobe|LOBE
Finding|Gene or Genome|SIMPLE_SEGMENT|2831,2835|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|LOBE
Event|Event|SIMPLE_SEGMENT|2836,2845|false|false|false|||LOBECTOMY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2836,2845|false|true|false|C0023928|Lobectomy|LOBECTOMY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2851,2859|false|false|false|C0018787|Heart|CORONARY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2851,2866|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2851,2874|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS SURGERY
Event|Event|SIMPLE_SEGMENT|2860,2866|false|false|false|||BYPASS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2860,2866|false|false|false|C0813207|Creation of shunt|BYPASS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2860,2874|false|false|false|C1536078|Bypass surgery|BYPASS SURGERY
Event|Event|SIMPLE_SEGMENT|2867,2874|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|2867,2874|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|2867,2874|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|2867,2874|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2867,2874|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|2883,2889|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2883,2897|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2890,2897|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2890,2897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2890,2897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2890,2897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2903,2909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2903,2909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2903,2909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2903,2909|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2903,2917|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2910,2917|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2910,2917|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2910,2917|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2910,2917|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2938,2946|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2938,2946|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2938,2946|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2938,2946|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2938,2951|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2938,2951|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2947,2951|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2947,2951|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2947,2951|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2953,2962|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2994,3000|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|2994,3000|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|2994,3000|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2994,3000|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2994,3000|false|false|false|C1305866|Weighing patient|weight
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3005,3008|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3010,3013|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3010,3013|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3014,3019|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|3014,3019|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|3014,3019|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|3014,3019|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|3024,3031|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3024,3031|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3024,3031|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|3038,3046|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|3038,3046|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|3053,3062|false|false|false|||gentleman
Event|Event|SIMPLE_SEGMENT|3063,3068|false|false|false|||lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3072,3075|false|false|true|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|3072,3075|false|false|true|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|3076,3084|false|false|false|||speaking
Finding|Individual Behavior|SIMPLE_SEGMENT|3076,3084|false|false|false|C0234856|Speaking (function)|speaking
Event|Event|SIMPLE_SEGMENT|3094,3103|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|3094,3103|false|false|false|C0876929|Sentence|sentences
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3107,3110|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3107,3110|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3107,3110|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3107,3110|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3107,3110|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3114,3119|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3121,3126|true|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3121,3126|true|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|3128,3132|true|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3137,3144|true|false|false|C0036410|Sclera|scleral
Finding|Finding|SIMPLE_SEGMENT|3137,3152|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|SIMPLE_SEGMENT|3145,3152|true|false|false|C0022346|Icterus|icterus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3154,3164|true|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|3165,3170|true|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3165,3170|true|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3174,3178|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3174,3178|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3174,3178|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3180,3186|true|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3180,3186|true|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|3188,3191|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3188,3191|true|false|false|C0428897|Jugular venous pressure|JVP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3203,3213|true|false|false|C0497156|Lymphadenopathy|adenopathy
Event|Event|SIMPLE_SEGMENT|3203,3213|true|false|false|||adenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|3203,3213|true|false|false|C4282165|Swollen Lymph Node|adenopathy
Event|Activity|SIMPLE_SEGMENT|3229,3233|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|3229,3233|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3229,3233|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|3238,3244|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|3238,3244|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3238,3244|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Functional Concept|SIMPLE_SEGMENT|3257,3268|false|false|false|C0205463|Physiological|physiologic
Finding|Functional Concept|SIMPLE_SEGMENT|3269,3274|false|false|false|C1534709|Splitting|split
Finding|Finding|SIMPLE_SEGMENT|3269,3277|false|false|false|C0425619|Second heart sound split|split S2
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3284,3292|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|3284,3299|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|SIMPLE_SEGMENT|3293,3299|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3293,3299|false|false|false|C0018808|Heart murmur|murmur
Finding|Finding|SIMPLE_SEGMENT|3293,3307|false|false|false|C2230293|murmur at left lower sternal border|murmur at LLSB
Event|Event|SIMPLE_SEGMENT|3303,3307|false|false|false|||LLSB
Event|Event|SIMPLE_SEGMENT|3312,3316|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|3312,3316|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|3320,3327|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3332,3337|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|3339,3343|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|3339,3343|true|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|3348,3356|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3348,3356|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|3358,3365|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3358,3365|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3370,3377|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3370,3377|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3381,3388|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3381,3388|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|3381,3388|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|3381,3388|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3390,3394|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3390,3394|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3400,3409|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|3400,3409|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3425,3429|false|false|false|C4318566|Deep Resection Margin|deep
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3425,3439|false|false|false|C0278328|Deep palpation|deep palpation
Event|Event|SIMPLE_SEGMENT|3430,3439|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3430,3439|false|false|false|C0030247|Palpation|palpation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3456,3459|true|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3456,3459|true|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|3456,3459|true|false|false|||CVA
Finding|Sign or Symptom|SIMPLE_SEGMENT|3456,3470|true|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|SIMPLE_SEGMENT|3460,3470|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3460,3470|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3460,3470|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|3490,3494|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3490,3494|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3490,3494|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3496,3500|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3501,3509|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3514,3520|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3514,3520|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3514,3520|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3514,3520|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|3524,3530|false|false|false|||radial
Finding|Conceptual Entity|SIMPLE_SEGMENT|3524,3530|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3542,3547|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3542,3547|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3542,3547|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3562,3567|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3562,3567|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3562,3579|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3568,3579|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3583,3588|false|false|false|C0022742|Knee|knees
Finding|Gene or Genome|SIMPLE_SEGMENT|3606,3609|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|SIMPLE_SEGMENT|3621,3627|true|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3621,3627|true|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3629,3635|true|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3642,3653|true|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Intellectual Product|SIMPLE_SEGMENT|3672,3678|true|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|3672,3683|true|false|false|C3266096|Stable gait|stable gait
Event|Event|SIMPLE_SEGMENT|3679,3683|true|false|false|||gait
Finding|Finding|SIMPLE_SEGMENT|3679,3683|true|false|false|C0016928|Gait|gait
Anatomy|Body System|SIMPLE_SEGMENT|3687,3691|true|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3687,3691|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3687,3691|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|SIMPLE_SEGMENT|3687,3691|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|SIMPLE_SEGMENT|3687,3691|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|SIMPLE_SEGMENT|3693,3697|true|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3693,3697|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3693,3697|true|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3699,3703|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3704,3712|true|false|false|||perfused
Event|Event|SIMPLE_SEGMENT|3722,3728|true|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3722,3728|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|3732,3739|true|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|3732,3739|true|false|false|C0221198|Lesion|lesions
Finding|Body Substance|SIMPLE_SEGMENT|3743,3752|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3743,3752|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3743,3752|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3743,3752|true|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3794,3798|false|false|false|||Tele
Finding|Gene or Genome|SIMPLE_SEGMENT|3794,3798|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Finding|Intellectual Product|SIMPLE_SEGMENT|3794,3798|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Event|Event|SIMPLE_SEGMENT|3803,3807|true|false|false|||tele
Finding|Gene or Genome|SIMPLE_SEGMENT|3803,3807|true|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Intellectual Product|SIMPLE_SEGMENT|3803,3807|true|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3859,3865|false|false|false|C0944911||Weight
Event|Event|SIMPLE_SEGMENT|3859,3865|false|false|false|||Weight
Finding|Finding|SIMPLE_SEGMENT|3859,3865|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|3859,3865|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|3859,3865|false|false|false|C1305866|Weighing patient|Weight
Event|Event|SIMPLE_SEGMENT|3869,3878|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3869,3878|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3893,3899|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|3893,3899|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|3893,3899|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|3893,3899|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|3893,3899|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|3907,3914|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3907,3914|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3907,3914|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3925,3928|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3925,3928|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3925,3928|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3925,3928|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3925,3928|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3925,3928|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3925,3928|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3931,3935|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3931,3935|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3931,3935|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3937,3940|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3937,3940|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3944,3948|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3944,3948|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3944,3948|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3944,3948|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|3944,3948|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|3944,3948|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3952,3960|false|false|false|C0008913|Bone structure of clavicle|clavicle
Event|Event|SIMPLE_SEGMENT|3969,3976|false|false|false|||degrees
Finding|Intellectual Product|SIMPLE_SEGMENT|3969,3976|false|false|false|C0542560|Academic degree|degrees
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3977,3982|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|SIMPLE_SEGMENT|3985,3989|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|3985,3989|true|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|3993,4001|true|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3993,4001|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|4006,4009|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|4011,4016|false|false|false|||split
Finding|Finding|SIMPLE_SEGMENT|4011,4019|false|false|false|C0425619|Second heart sound split|split S2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4020,4027|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4020,4027|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|4020,4027|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|4020,4027|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4038,4043|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|4038,4043|false|false|false|||obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4045,4049|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4045,4049|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|4057,4061|false|false|false|||NABS
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4062,4065|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|4062,4065|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|4062,4065|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4070,4075|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4070,4075|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4070,4075|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|SIMPLE_SEGMENT|4097,4106|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4119,4124|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4119,4124|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4119,4124|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4125,4128|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4133,4136|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4133,4136|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4133,4136|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4143,4146|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4143,4146|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4143,4146|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4143,4146|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4153,4156|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4153,4156|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4164,4167|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4164,4167|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4164,4167|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4164,4167|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4164,4167|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4172,4175|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4172,4175|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4172,4175|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4172,4175|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4172,4175|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4172,4175|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4181,4185|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4181,4185|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4213,4216|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4233,4238|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4233,4238|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4233,4238|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4243,4246|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4243,4246|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4243,4246|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4268,4273|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4268,4273|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4268,4273|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4268,4281|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4268,4281|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4268,4281|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4274,4281|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4274,4281|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4274,4281|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4274,4281|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4274,4281|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4274,4281|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4326,4330|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4326,4330|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4326,4330|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4355,4360|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4355,4360|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4355,4360|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4361,4364|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4361,4364|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4361,4364|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4361,4364|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4361,4364|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4361,4364|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4361,4364|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4361,4364|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4369,4372|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4369,4372|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4369,4372|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4369,4372|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4369,4372|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4369,4372|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4369,4372|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4377,4384|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4377,4384|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4412,4417|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4412,4417|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4412,4417|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4418,4423|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4418,4423|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4418,4423|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4418,4423|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|4421,4425|false|false|false|C0602254|MB 3|MB-3
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4440,4446|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|4440,4446|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4465,4470|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4465,4470|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4465,4470|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4465,4478|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4471,4478|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4471,4478|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4471,4478|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|4471,4478|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|4471,4478|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|4471,4478|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4471,4478|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4483,4490|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4483,4490|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4483,4490|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4483,4490|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4483,4490|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4483,4490|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4483,4490|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4483,4490|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4514,4519|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4514,4519|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4514,4519|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4520,4527|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4520,4527|false|false|false|C0060323|Fibrin fragment D|D-Dimer
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4522,4527|false|false|false|C0596448|dimer|Dimer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4545,4550|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4545,4550|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4545,4550|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4551,4554|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4551,4554|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|4551,4554|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4551,4554|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|4551,4554|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4551,4554|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Finding|Body Substance|SIMPLE_SEGMENT|4560,4569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4560,4569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4560,4569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4560,4569|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4582,4587|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4582,4587|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4582,4587|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4588,4591|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4597,4600|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4597,4600|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4597,4600|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4607,4610|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4607,4610|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4607,4610|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4607,4610|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4617,4620|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4617,4620|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4628,4631|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4628,4631|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4628,4631|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4628,4631|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4628,4631|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4636,4639|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4636,4639|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4636,4639|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4636,4639|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4636,4639|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4636,4639|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4645,4649|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4645,4649|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4677,4680|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4697,4702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4697,4702|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4697,4702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4707,4710|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4707,4710|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4707,4710|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4732,4737|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4732,4737|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4732,4737|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4732,4745|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4732,4745|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4732,4745|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4738,4745|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4738,4745|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4738,4745|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4738,4745|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4738,4745|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4738,4745|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4822,4827|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4822,4827|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4822,4827|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4828,4831|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4828,4831|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4828,4831|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4828,4831|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4828,4831|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4828,4831|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4828,4831|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4828,4831|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4836,4839|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4836,4839|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4836,4839|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4836,4839|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4836,4839|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4836,4839|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4836,4839|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4844,4851|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4844,4851|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4879,4884|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4879,4884|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4879,4884|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4879,4892|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4885,4892|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4885,4892|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4885,4892|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4885,4892|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4885,4892|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4885,4892|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4885,4892|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4885,4892|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4915,4919|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|4915,4919|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4915,4919|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|SIMPLE_SEGMENT|4928,4932|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4928,4939|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4933,4939|false|false|false|C0018792|Heart Atrium|atrium
Finding|Finding|SIMPLE_SEGMENT|4943,4953|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Event|Event|SIMPLE_SEGMENT|4954,4961|false|false|false|||dilated
Finding|Functional Concept|SIMPLE_SEGMENT|4967,4972|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4967,4979|false|false|false|C0225844|Right atrial structure|right atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4973,4979|false|false|false|C0018792|Heart Atrium|atrium
Finding|Finding|SIMPLE_SEGMENT|4984,4994|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Event|Event|SIMPLE_SEGMENT|4995,5002|false|false|false|||dilated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5007,5013|true|false|false|C0018792|Heart Atrium|atrial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5007,5027|true|false|false|C0018817|Atrial Septal Defects|atrial septal defect
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5014,5027|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5014,5027|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5021,5027|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|5021,5027|true|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|5021,5027|true|false|false|C1457869|Defect|defect
Event|Event|SIMPLE_SEGMENT|5031,5035|true|false|false|||seen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5046,5051|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5046,5051|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Event|Event|SIMPLE_SEGMENT|5046,5051|false|false|false|||color
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5046,5059|false|false|false|C0474781|Color doppler ultrasound|color Doppler
Event|Event|SIMPLE_SEGMENT|5052,5059|false|false|false|||Doppler
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5052,5059|false|false|false|C0554756|Doppler studies|Doppler
Finding|Functional Concept|SIMPLE_SEGMENT|5061,5065|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5061,5082|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5066,5077|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5066,5082|false|false|false|C0507618|Wall of ventricle|ventricular wall
Event|Event|SIMPLE_SEGMENT|5083,5094|false|false|false|||thicknesses
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5099,5105|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5099,5105|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5099,5105|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5116,5122|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|5133,5137|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|5147,5151|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5152,5163|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|5164,5172|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5164,5172|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5174,5185|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|5174,5185|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|5174,5185|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|5174,5185|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|5174,5185|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|SIMPLE_SEGMENT|5191,5202|false|false|false|||hypokinesis
Finding|Finding|SIMPLE_SEGMENT|5191,5202|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|SIMPLE_SEGMENT|5239,5247|false|false|false|||inferior
Finding|Social Behavior|SIMPLE_SEGMENT|5239,5247|false|false|false|C0678975|inferiority|inferior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5268,5275|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|5268,5275|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Finding|SIMPLE_SEGMENT|5268,5281|false|false|false|C0428776|Cardiac index|cardiac index
Event|Event|SIMPLE_SEGMENT|5276,5281|false|false|false|||index
Finding|Idea or Concept|SIMPLE_SEGMENT|5276,5281|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|SIMPLE_SEGMENT|5276,5281|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Event|Event|SIMPLE_SEGMENT|5285,5291|false|false|false|||normal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5310,5317|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|SIMPLE_SEGMENT|5318,5328|false|false|false|||parameters
Finding|Finding|SIMPLE_SEGMENT|5318,5328|false|false|false|C0449381|Observation parameter|parameters
Event|Event|SIMPLE_SEGMENT|5333,5346|false|false|false|||indeterminate
Event|Event|SIMPLE_SEGMENT|5351,5355|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|5351,5355|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5357,5368|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5369,5378|false|false|false|C0012000|Diastole|diastolic
Event|Event|SIMPLE_SEGMENT|5379,5387|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5379,5387|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5379,5387|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5379,5387|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5379,5387|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5393,5398|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5393,5417|false|false|false|C0503854|Cavity of right ventricle|right ventricular cavity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5399,5410|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5399,5417|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5411,5417|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5411,5417|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5411,5417|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5429,5436|false|false|false|||dilated
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5442,5451|false|false|false|C0344315|Depressed mood|depressed
Event|Event|SIMPLE_SEGMENT|5452,5456|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5452,5456|false|false|false|C0332296|Free of (attribute)|free
Event|Event|SIMPLE_SEGMENT|5462,5475|true|false|false|||contractility
Finding|Finding|SIMPLE_SEGMENT|5462,5475|true|false|false|C5424789|Contractility|contractility
Event|Event|SIMPLE_SEGMENT|5480,5484|true|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5480,5484|true|false|false|C0332296|Free of (attribute)|free
Finding|Finding|SIMPLE_SEGMENT|5498,5502|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5503,5507|true|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5514,5520|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5514,5526|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5521,5526|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5527,5535|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5552,5561|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5566,5572|true|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|SIMPLE_SEGMENT|5566,5581|true|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|SIMPLE_SEGMENT|5573,5581|true|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5573,5581|true|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|5589,5596|true|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|5589,5596|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|5589,5596|true|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5602,5614|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5609,5614|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5616,5624|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5636,5645|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5659,5671|true|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5666,5671|true|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5673,5681|true|false|false|C0033377|Ptosis|prolapse
Event|Event|SIMPLE_SEGMENT|5673,5681|true|false|false|||prolapse
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5691,5711|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|5698,5711|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5698,5711|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5698,5711|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5698,5711|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|5715,5719|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5736,5741|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5742,5750|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5762,5771|false|false|false|||thickened
Finding|Finding|SIMPLE_SEGMENT|5773,5781|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|5773,5781|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|5798,5811|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5798,5811|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5798,5811|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5798,5811|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|5815,5819|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|5830,5838|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|5830,5838|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5839,5848|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5839,5848|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5839,5848|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5839,5855|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5849,5855|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5849,5855|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5857,5865|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5857,5878|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5866,5878|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5866,5878|false|false|false|||hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5884,5898|false|false|false|C0034086|Pulmonary valve structure|pulmonic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5893,5898|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5899,5907|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5913,5922|false|false|false|||thickened
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5936,5947|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5936,5947|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5936,5956|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|5936,5956|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|5948,5956|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5948,5956|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5948,5956|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5948,5956|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5960,5970|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5960,5970|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5960,5970|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5972,5976|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Functional Concept|SIMPLE_SEGMENT|5986,5990|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Pathologic Function|SIMPLE_SEGMENT|5986,6014|false|false|false|C0242698|Ventricular Dysfunction, Left|left ventricular dysfunction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5991,6002|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|SIMPLE_SEGMENT|5991,6014|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6003,6014|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|6003,6014|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|6003,6014|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|6003,6014|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|6003,6014|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6032,6035|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6032,6035|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6032,6035|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6032,6035|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6032,6035|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6032,6035|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6032,6035|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6032,6035|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Intellectual Product|SIMPLE_SEGMENT|6042,6049|false|false|false|C0282416|Overall Publication Type|overall
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6057,6066|false|false|false|C0344315|Depressed mood|depressed
Event|Event|SIMPLE_SEGMENT|6057,6066|false|false|false|||depressed
Event|Event|SIMPLE_SEGMENT|6074,6082|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6074,6082|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|6084,6092|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|6084,6092|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|6084,6092|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|6084,6092|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|6084,6092|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|6101,6108|false|false|false|||dilated
Finding|Functional Concept|SIMPLE_SEGMENT|6109,6114|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6109,6124|false|false|false|C0225883|Right ventricular structure|right ventricle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6115,6124|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6115,6124|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6130,6139|false|false|false|C0344315|Depressed mood|depressed
Event|Event|SIMPLE_SEGMENT|6140,6144|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|6140,6144|false|false|false|C0332296|Free of (attribute)|free
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6151,6159|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|6160,6168|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|6160,6168|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|6160,6168|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|6160,6168|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|6160,6168|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|SIMPLE_SEGMENT|6170,6178|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6170,6178|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Finding|SIMPLE_SEGMENT|6170,6202|false|false|false|C3276922|Tricuspid regurgitation, moderate|Moderate tricuspid regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6179,6202|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|SIMPLE_SEGMENT|6189,6202|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|6189,6202|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|6189,6202|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|6189,6202|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Finding|SIMPLE_SEGMENT|6209,6217|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6209,6217|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Pathologic Function|SIMPLE_SEGMENT|6209,6240|false|false|false|C5395246|Moderate pulmonary hypertension|moderate pulmonary hypertension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6218,6227|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6218,6227|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6218,6227|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|6218,6240|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6228,6240|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|6228,6240|false|false|false|||hypertension
Finding|Intellectual Product|SIMPLE_SEGMENT|6246,6251|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6252,6260|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6252,6267|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6252,6267|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|6287,6291|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|6287,6291|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|6292,6295|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|6311,6318|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6311,6318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6311,6318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6311,6318|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6311,6321|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6322,6325|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6322,6325|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6322,6325|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6322,6325|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6322,6325|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6322,6325|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6322,6325|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6322,6325|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6332,6336|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6332,6336|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6341,6344|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6341,6344|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|SIMPLE_SEGMENT|6341,6344|false|false|false|||PCI
Finding|Gene or Genome|SIMPLE_SEGMENT|6341,6344|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|SIMPLE_SEGMENT|6341,6344|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6341,6344|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6347,6350|false|false|false|C0235480;C0393911|Paroxysmal atrial fibrillation;Pure Autonomic Failure|pAF
Drug|Immunologic Factor|SIMPLE_SEGMENT|6347,6350|false|false|false|C0032172|Platelet Activating Factor|pAF
Drug|Organic Chemical|SIMPLE_SEGMENT|6347,6350|false|false|false|C0032172|Platelet Activating Factor|pAF
Event|Event|SIMPLE_SEGMENT|6347,6350|false|false|false|||pAF
Finding|Gene or Genome|SIMPLE_SEGMENT|6347,6350|false|false|false|C1537443|PCLAF gene|pAF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6347,6350|false|false|false|C0279389|doxorubicin/fluorouracil/melphalan protocol|pAF
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6352,6355|false|false|false|C0265910;C2973725;C3203102|Congenital hypoplasia of pulmonary artery;Idiopathic pulmonary arterial hypertension;Pulmonary arterial hypertension|PAH
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6352,6355|false|false|false|C0265910;C2973725;C3203102|Congenital hypoplasia of pulmonary artery;Idiopathic pulmonary arterial hypertension;Pulmonary arterial hypertension|PAH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6352,6355|false|false|false|C0030123;C0032458;C5890890|4-aminohippuric acid;PAH protein, human;Polycyclic Hydrocarbons, Aromatic|PAH
Drug|Enzyme|SIMPLE_SEGMENT|6352,6355|false|false|false|C0030123;C0032458;C5890890|4-aminohippuric acid;PAH protein, human;Polycyclic Hydrocarbons, Aromatic|PAH
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6352,6355|false|false|false|C0030123;C0032458;C5890890|4-aminohippuric acid;PAH protein, human;Polycyclic Hydrocarbons, Aromatic|PAH
Drug|Organic Chemical|SIMPLE_SEGMENT|6352,6355|false|false|false|C0030123;C0032458;C5890890|4-aminohippuric acid;PAH protein, human;Polycyclic Hydrocarbons, Aromatic|PAH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6352,6355|false|false|false|C0030123;C0032458;C5890890|4-aminohippuric acid;PAH protein, human;Polycyclic Hydrocarbons, Aromatic|PAH
Event|Event|SIMPLE_SEGMENT|6352,6355|false|false|false|||PAH
Finding|Gene or Genome|SIMPLE_SEGMENT|6352,6355|false|false|false|C1418251;C2247505|PAH gene;proclavaminate amidinohydrolase activity|PAH
Finding|Molecular Function|SIMPLE_SEGMENT|6352,6355|false|false|false|C1418251;C2247505|PAH gene;proclavaminate amidinohydrolase activity|PAH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6352,6355|false|false|false|C3540097|PAH gene (lab test)|PAH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6357,6366|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6357,6370|false|false|false|C2183328|diastolic congestive heart failure|diastolic CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6367,6370|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6367,6370|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|6367,6370|false|false|false|||CHF
Event|Event|SIMPLE_SEGMENT|6375,6383|false|false|false|||presents
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6390,6396|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|6390,6396|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|6390,6396|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|6390,6396|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|6390,6396|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|6390,6401|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Finding|Intellectual Product|SIMPLE_SEGMENT|6390,6401|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Event|Event|SIMPLE_SEGMENT|6397,6401|false|false|false|||gain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6403,6406|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|6403,6415|false|false|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|SIMPLE_SEGMENT|6407,6415|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|6407,6415|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|6407,6415|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|SIMPLE_SEGMENT|6420,6423|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6420,6423|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|6424,6432|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|6424,6432|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6424,6435|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|6436,6441|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6436,6451|false|false|false|C0225883|Right ventricular structure|right ventricle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6442,6451|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6442,6451|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Event|Event|SIMPLE_SEGMENT|6453,6461|false|false|false|||dilation
Finding|Finding|SIMPLE_SEGMENT|6453,6461|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Finding|Pathologic Function|SIMPLE_SEGMENT|6453,6461|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6453,6461|false|false|false|C1322279|Dilate procedure|dilation
Finding|Intellectual Product|SIMPLE_SEGMENT|6477,6482|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6477,6507|false|true|false|C4087508|Acute exacerbation of chronic heart failure|acute on chronic heart failure
Finding|Intellectual Product|SIMPLE_SEGMENT|6486,6493|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6486,6493|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6486,6507|false|false|false|C0264716|Chronic heart failure|chronic heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6494,6499|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6494,6499|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6494,6499|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6494,6507|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|6500,6507|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|6500,6507|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|6500,6507|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|6500,6507|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|6509,6521|false|false|false|||exacerbation
Finding|Finding|SIMPLE_SEGMENT|6509,6521|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|SIMPLE_SEGMENT|6527,6532|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6527,6567|false|false|false|C2732749|Acute on chronic diastolic heart failure|Acute on Chronic Diastolic Heart Failure
Finding|Intellectual Product|SIMPLE_SEGMENT|6536,6543|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6536,6543|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6536,6567|false|false|false|C2711480|Chronic diastolic heart failure|Chronic Diastolic Heart Failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6544,6553|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6544,6567|false|false|false|C1135196|Heart Failure, Diastolic|Diastolic Heart Failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6554,6559|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6554,6559|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6554,6559|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6554,6567|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|Heart Failure
Finding|Functional Concept|SIMPLE_SEGMENT|6560,6567|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|6560,6567|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|6560,6567|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Event|Event|SIMPLE_SEGMENT|6568,6580|false|false|false|||Exacerbation
Finding|Finding|SIMPLE_SEGMENT|6568,6580|false|false|false|C4086268|Exacerbation|Exacerbation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6588,6597|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6588,6597|false|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|6588,6597|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|6588,6597|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|6588,6597|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|6588,6597|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|SIMPLE_SEGMENT|6604,6611|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|6604,6611|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|6604,6611|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|6604,6611|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6615,6621|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|6615,6621|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|6615,6621|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|6615,6621|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|6629,6633|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|6629,6633|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6629,6633|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Finding|SIMPLE_SEGMENT|6636,6642|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6636,6642|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6652,6659|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6652,6659|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|6652,6659|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|6652,6659|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6652,6659|false|false|false|C1522240|Process|process
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6663,6667|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6663,6667|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6663,6667|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|6663,6667|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6663,6675|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6668,6675|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6668,6675|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|6676,6683|false|false|false|||causing
Finding|Finding|SIMPLE_SEGMENT|6684,6695|false|false|false|C5539458|Elevated residual volume|elevated RV
Event|Event|SIMPLE_SEGMENT|6696,6705|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|6696,6705|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6696,6705|false|false|false|C0033095||pressures
Finding|Intellectual Product|SIMPLE_SEGMENT|6722,6726|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|6727,6734|false|false|false|||filling
Event|Event|SIMPLE_SEGMENT|6746,6754|false|false|false|||diuresed
Event|Event|SIMPLE_SEGMENT|6761,6765|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|6761,6765|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|6778,6783|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6778,6783|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|6778,6783|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|6793,6803|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6793,6803|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6793,6808|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|6812,6819|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|6812,6819|false|true|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|6812,6819|false|true|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|6812,6819|false|true|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|6822,6829|false|false|false|||Started
Drug|Organic Chemical|SIMPLE_SEGMENT|6834,6843|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6834,6843|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|6834,6843|false|false|false|||torsemide
Finding|Finding|SIMPLE_SEGMENT|6865,6871|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6865,6871|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|6876,6886|false|false|false|||aggressive
Finding|Individual Behavior|SIMPLE_SEGMENT|6876,6886|false|true|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|6876,6886|false|true|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Event|Event|SIMPLE_SEGMENT|6893,6901|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|6905,6909|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|6905,6909|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6905,6909|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|SIMPLE_SEGMENT|6914,6918|false|false|false|||read
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6919,6922|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|6919,6922|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|6919,6922|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Finding|Finding|SIMPLE_SEGMENT|6926,6930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|6926,6930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|6926,6930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|6934,6943|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6934,6943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6934,6943|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|6949,6953|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|6959,6963|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6959,6963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6959,6963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6959,6963|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6969,6977|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|SIMPLE_SEGMENT|6978,6985|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|6978,6985|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6978,6985|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Organic Chemical|SIMPLE_SEGMENT|6989,6998|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6989,6998|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|6989,6998|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|7016,7028|false|false|false|||discontinued
Finding|Idea or Concept|SIMPLE_SEGMENT|7029,7033|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7029,7033|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7029,7033|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7034,7045|false|false|false|C0040869|triamterene|triamterene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7034,7045|false|false|false|C0040869|triamterene|triamterene
Event|Event|SIMPLE_SEGMENT|7034,7045|false|false|false|||triamterene
Drug|Organic Chemical|SIMPLE_SEGMENT|7046,7050|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7046,7050|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|7046,7050|false|false|false|||HCTZ
Finding|Finding|SIMPLE_SEGMENT|7054,7059|false|false|false|C0587267;C3810854|Close;Closed|Close
Finding|Functional Concept|SIMPLE_SEGMENT|7054,7059|false|false|false|C0587267;C3810854|Close;Closed|Close
Finding|Functional Concept|SIMPLE_SEGMENT|7060,7066|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|7060,7066|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|7060,7069|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|7060,7069|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|7067,7069|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|7084,7091|false|false|false|||ensured
Finding|Finding|SIMPLE_SEGMENT|7095,7117|false|false|false|C0438717;C2242708|Hypertransaminasaemia;Transaminases increased|Elevated Transaminases
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7104,7117|false|false|false|C0002594|Transaminases|Transaminases
Drug|Enzyme|SIMPLE_SEGMENT|7104,7117|false|false|false|C0002594|Transaminases|Transaminases
Event|Event|SIMPLE_SEGMENT|7104,7117|false|false|false|||Transaminases
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7104,7117|false|false|false|C0919834|Transaminase Assay|Transaminases
Finding|Body Substance|SIMPLE_SEGMENT|7120,7127|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7120,7127|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7120,7127|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|7140,7152|false|false|false|C0151904|Aspartate Aminotransferase Increased|elevated AST
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7149,7152|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7149,7152|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7149,7152|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7149,7152|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|7149,7152|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|7149,7152|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|7149,7152|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7158,7161|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7158,7161|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|7158,7161|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|7158,7161|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|7158,7161|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|7158,7161|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|7158,7161|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7158,7161|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Finding|Idea or Concept|SIMPLE_SEGMENT|7163,7174|false|false|false|C0750501|most likely|Most likely
Finding|Finding|SIMPLE_SEGMENT|7168,7174|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7168,7174|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|7175,7185|false|false|false|||etiologies
Finding|Functional Concept|SIMPLE_SEGMENT|7175,7185|false|true|false|C0015127|Etiology aspects|etiologies
Finding|Body Substance|SIMPLE_SEGMENT|7194,7201|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7194,7201|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7194,7201|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|7210,7220|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7210,7220|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|7210,7220|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7210,7220|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7222,7230|false|false|false|C0600688|Toxic effect|toxicity
Event|Event|SIMPLE_SEGMENT|7222,7230|false|false|false|||toxicity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7235,7257|false|false|false|C5243996|Congestive hepatopathy|congestive hepatopathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7246,7257|false|false|false|C0023895|Liver diseases|hepatopathy
Event|Event|SIMPLE_SEGMENT|7246,7257|false|false|false|||hepatopathy
Event|Event|SIMPLE_SEGMENT|7271,7281|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|7271,7281|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7271,7281|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|7283,7291|false|false|false|||trending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7296,7305|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7296,7305|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|7296,7305|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7296,7313|false|false|false|C0024115|Lung diseases|Pulmonary disease
Finding|Finding|SIMPLE_SEGMENT|7296,7313|false|false|false|C0455540|History of - respiratory disease|Pulmonary disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7306,7313|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7306,7313|false|false|false|||disease
Finding|Body Substance|SIMPLE_SEGMENT|7315,7322|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7315,7322|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7315,7322|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7338,7347|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|SIMPLE_SEGMENT|7338,7347|false|false|false|||emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|7338,7347|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7351,7354|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|7351,7354|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|7351,7354|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7351,7354|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Body Substance|SIMPLE_SEGMENT|7363,7370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7363,7370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7363,7370|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|7363,7374|true|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|7378,7385|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7378,7385|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7378,7385|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7378,7385|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7378,7388|true|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|7389,7396|true|false|false|||smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|7389,7396|true|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|7389,7396|true|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Event|Event|SIMPLE_SEGMENT|7415,7422|false|false|false|||driving
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7415,7422|false|false|false|C0004379|Automobile Driving|driving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7425,7430|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7425,7430|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|7425,7430|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7425,7438|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|7431,7438|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|7431,7438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|7431,7438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|7431,7438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|7458,7469|false|false|false|||pulmonology
Event|Event|SIMPLE_SEGMENT|7471,7478|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|7471,7478|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|7488,7497|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7488,7497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7488,7497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7488,7497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7488,7497|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|7502,7509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7502,7509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7502,7509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7514,7523|false|false|false|||insistent
Event|Event|SIMPLE_SEGMENT|7527,7534|false|false|false|||leaving
Finding|Classification|SIMPLE_SEGMENT|7556,7566|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7556,7566|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Activity|SIMPLE_SEGMENT|7567,7578|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|7567,7578|false|false|false|||appointment
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7584,7590|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7584,7603|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7584,7603|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7584,7603|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7591,7603|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|SIMPLE_SEGMENT|7591,7603|false|false|false|||Fibrillation
Event|Event|SIMPLE_SEGMENT|7605,7613|false|false|false|||Continue
Finding|Idea or Concept|SIMPLE_SEGMENT|7614,7618|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7614,7618|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7614,7618|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7619,7629|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7619,7629|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|7619,7629|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7619,7629|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|7644,7652|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7644,7652|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7657,7660|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7657,7660|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7657,7660|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7657,7660|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7657,7660|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7665,7668|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7665,7668|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|7665,7668|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|7665,7668|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7665,7668|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7665,7668|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|7665,7668|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7665,7668|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|7670,7678|false|false|false|||Continue
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7679,7682|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|7679,7682|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|7679,7682|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7679,7682|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|7679,7682|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|7679,7682|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|7689,7701|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7689,7701|false|false|false|C0965129|rosuvastatin|rosuvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7715,7718|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|7715,7718|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|7720,7728|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|7729,7733|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7729,7733|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7729,7733|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|7734,7742|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7734,7742|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|7734,7742|false|false|false|||losartan
Event|Event|SIMPLE_SEGMENT|7748,7750|false|false|false|||qD
Finding|Idea or Concept|SIMPLE_SEGMENT|7753,7765|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Finding|SIMPLE_SEGMENT|7776,7779|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|7776,7779|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7780,7790|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|7780,7790|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7780,7790|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|SIMPLE_SEGMENT|7792,7801|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7792,7801|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|SIMPLE_SEGMENT|7829,7840|false|false|false|C0040869|triamterene|triamterene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7829,7840|false|false|false|C0040869|triamterene|triamterene
Event|Event|SIMPLE_SEGMENT|7829,7840|false|false|false|||triamterene
Drug|Organic Chemical|SIMPLE_SEGMENT|7841,7845|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7841,7845|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|7841,7845|false|false|false|||HCTZ
Drug|Organic Chemical|SIMPLE_SEGMENT|7849,7854|false|false|false|C0309049|favor|favor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7849,7854|false|false|false|C0309049|favor|favor
Drug|Vitamin|SIMPLE_SEGMENT|7849,7854|false|false|false|C0309049|favor|favor
Event|Event|SIMPLE_SEGMENT|7849,7854|false|false|false|||favor
Event|Event|SIMPLE_SEGMENT|7858,7863|false|false|false|||above
Finding|Idea or Concept|SIMPLE_SEGMENT|7858,7863|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|7867,7871|false|false|false|||LFTs
Finding|Intellectual Product|SIMPLE_SEGMENT|7872,7876|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|7877,7885|false|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|7896,7904|false|false|false|||consider
Event|Event|SIMPLE_SEGMENT|7905,7913|false|false|false|||possible
Finding|Finding|SIMPLE_SEGMENT|7905,7913|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|7915,7928|false|false|false|||discontinuing
Finding|Functional Concept|SIMPLE_SEGMENT|7929,7937|false|false|false|C0392747|Changing|changing
Drug|Organic Chemical|SIMPLE_SEGMENT|7938,7948|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7938,7948|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|7938,7948|false|false|false|||amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7938,7948|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Event|Event|SIMPLE_SEGMENT|7959,7964|false|false|false|||check
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7965,7968|false|false|false|C5816720|Isolated lipoma of filum terminale|LFT
Finding|Gene or Genome|SIMPLE_SEGMENT|7965,7968|false|false|false|C1537580|LIX1 gene|LFT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7965,7968|false|false|false|C0023901|Liver Function Tests|LFT
Event|Event|SIMPLE_SEGMENT|7965,7970|false|false|false|||LFT's
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7965,7970|false|false|false|C0023901|Liver Function Tests|LFT's
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7975,7985|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7975,7985|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|7975,7985|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7975,7985|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7975,7985|false|false|false|C0201975|Creatinine measurement|Creatinine
Finding|Functional Concept|SIMPLE_SEGMENT|7989,7995|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|7989,7995|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|7989,7998|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|7989,7998|false|false|false|C1522577|follow-up|follow up
Event|Activity|SIMPLE_SEGMENT|7999,8010|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|8026,8034|false|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|8041,8053|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|8057,8063|false|false|false|||Follow
Event|Activity|SIMPLE_SEGMENT|8067,8078|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|8067,8078|false|false|false|||appointment
Anatomy|Body System|SIMPLE_SEGMENT|8084,8094|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|SIMPLE_SEGMENT|8107,8113|false|false|false|||Follow
Event|Activity|SIMPLE_SEGMENT|8117,8128|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|8117,8128|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|8149,8155|false|false|false|||Follow
Event|Activity|SIMPLE_SEGMENT|8159,8170|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|8159,8170|false|false|false|||appointment
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8176,8179|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8176,8179|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8176,8179|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8176,8179|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8176,8179|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8176,8179|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8176,8179|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8176,8179|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|8176,8179|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8176,8179|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8176,8179|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8194,8200|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|8194,8200|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|8194,8200|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|8194,8200|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|8194,8200|false|false|false|C1305866|Weighing patient|weight
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8216,8227|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8216,8227|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8216,8227|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8216,8227|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8216,8240|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8231,8240|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8231,8240|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8259,8269|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8259,8269|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8259,8274|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8270,8274|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8270,8274|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8278,8286|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|8291,8299|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8291,8299|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8291,8299|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|8291,8299|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|8291,8299|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8291,8299|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8304,8314|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8304,8314|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|8304,8314|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8304,8314|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|8335,8343|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8335,8343|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8352,8355|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8352,8355|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8352,8355|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8352,8355|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8352,8355|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8360,8367|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8360,8367|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8387,8395|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8387,8395|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|8387,8395|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|8387,8402|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8387,8402|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8396,8402|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8396,8402|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8396,8402|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|8396,8402|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8396,8402|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8396,8402|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8413,8416|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8413,8416|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8413,8416|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8413,8416|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8413,8416|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8421,8429|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8421,8429|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8421,8429|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|8421,8439|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8421,8439|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8430,8439|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8430,8439|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|8430,8439|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8430,8439|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8430,8439|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|8430,8439|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|8430,8439|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8430,8439|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|8459,8469|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8459,8469|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|8489,8500|false|false|false|C0040869|triamterene|Triamterene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8489,8500|false|false|false|C0040869|triamterene|Triamterene
Drug|Organic Chemical|SIMPLE_SEGMENT|8501,8505|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8501,8505|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|8501,8505|false|false|false|||HCTZ
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8518,8521|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8518,8521|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|SIMPLE_SEGMENT|8518,8521|false|false|false|||CAP
Finding|Gene or Genome|SIMPLE_SEGMENT|8518,8521|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8518,8521|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|SIMPLE_SEGMENT|8535,8540|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8535,8540|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|SIMPLE_SEGMENT|8559,8564|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8559,8564|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8566,8590|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|SIMPLE_SEGMENT|8582,8590|false|false|false|||infantis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8597,8601|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8597,8601|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|8597,8601|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|8597,8601|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|8602,8607|false|false|false|||DAILY
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8613,8621|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|SIMPLE_SEGMENT|8613,8621|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|SIMPLE_SEGMENT|8613,8621|false|false|false|||coenzyme
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8613,8625|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|SIMPLE_SEGMENT|8613,8625|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8613,8625|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|SIMPLE_SEGMENT|8622,8625|false|false|false|||Q10
Finding|Gene or Genome|SIMPLE_SEGMENT|8622,8625|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8633,8637|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8633,8637|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|8633,8637|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|8633,8637|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|8638,8643|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|8649,8661|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8649,8661|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Event|Event|SIMPLE_SEGMENT|8649,8661|false|false|false|||Rosuvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8649,8669|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8649,8669|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8662,8669|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8662,8669|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8662,8669|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8662,8669|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|8662,8669|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|8662,8669|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|8662,8669|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8662,8669|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8662,8672|false|false|false|C0006675|calcium|Calcium 40
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8662,8672|false|false|false|C0006675|calcium|Calcium 40
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8662,8672|false|false|false|C0006675|calcium|Calcium 40
Event|Event|SIMPLE_SEGMENT|8679,8682|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|8688,8695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8688,8695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|8688,8695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|8688,8697|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|8688,8697|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8688,8697|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|8688,8697|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Event|Event|SIMPLE_SEGMENT|8688,8697|false|false|false|||Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8688,8697|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|8708,8710|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|8722,8732|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8722,8732|false|false|false|C0257343|tamsulosin|Tamsulosin
Event|Event|SIMPLE_SEGMENT|8751,8760|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8751,8760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8751,8760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8751,8760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8751,8760|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8751,8772|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8761,8772|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8761,8772|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8761,8772|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8761,8772|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8777,8787|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8777,8787|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|8777,8787|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8777,8787|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|SIMPLE_SEGMENT|8808,8816|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8808,8816|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8825,8828|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8825,8828|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8825,8828|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8825,8828|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8825,8828|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8860,8868|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8860,8868|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|8860,8868|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|8860,8875|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8860,8875|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8869,8875|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8869,8875|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8869,8875|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|8869,8875|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8869,8875|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8869,8875|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8886,8889|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8886,8889|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8886,8889|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8886,8889|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8886,8889|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|8894,8902|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8894,8902|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8894,8902|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|8894,8912|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8894,8912|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8903,8912|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8903,8912|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|8903,8912|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8903,8912|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8903,8912|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|8903,8912|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|8903,8912|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8903,8912|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|8932,8944|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8932,8944|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Event|Event|SIMPLE_SEGMENT|8932,8944|false|false|false|||Rosuvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8932,8952|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8932,8952|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8945,8952|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8945,8952|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8945,8952|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8945,8952|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|8945,8952|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|8945,8952|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|8945,8952|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8945,8952|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8945,8955|false|false|false|C0006675|calcium|Calcium 40
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8945,8955|false|false|false|C0006675|calcium|Calcium 40
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8945,8955|false|false|false|C0006675|calcium|Calcium 40
Event|Event|SIMPLE_SEGMENT|8962,8965|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|8970,8975|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8970,8975|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|SIMPLE_SEGMENT|8995,9005|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8995,9005|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Organic Chemical|SIMPLE_SEGMENT|9007,9012|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9007,9012|false|false|false|C3489575|sennosides, USP|senna
Event|Event|SIMPLE_SEGMENT|9007,9012|false|false|false|||senna
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9023,9030|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|9023,9030|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9023,9030|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|9031,9039|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9034,9039|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9034,9039|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|9040,9044|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9040,9050|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|9047,9050|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9047,9050|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|9051,9055|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|9051,9055|false|false|false|C2828567|PRSS30P gene|Disp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9062,9069|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|9062,9069|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9062,9069|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|9070,9077|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9070,9077|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9084,9091|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9084,9091|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9084,9091|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9084,9093|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9084,9093|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9084,9093|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9084,9093|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9084,9093|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9092,9093|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|9099,9103|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|9117,9126|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9117,9126|false|false|false|C0076840|torsemide|Torsemide
Event|Event|SIMPLE_SEGMENT|9142,9144|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|9146,9155|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9146,9155|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|9146,9155|false|false|false|||torsemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9163,9169|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9173,9181|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9176,9181|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9176,9181|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|SIMPLE_SEGMENT|9182,9186|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9182,9192|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|9189,9192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9189,9192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9204,9210|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9211,9218|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9211,9218|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9226,9231|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9226,9231|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9233,9257|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|SIMPLE_SEGMENT|9249,9257|false|false|false|||infantis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9264,9268|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9264,9268|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9264,9268|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9264,9268|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|9269,9274|false|false|false|||DAILY
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9280,9288|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|SIMPLE_SEGMENT|9280,9288|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|SIMPLE_SEGMENT|9280,9288|false|false|false|||coenzyme
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9280,9292|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|SIMPLE_SEGMENT|9280,9292|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9280,9292|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|SIMPLE_SEGMENT|9289,9292|false|false|false|||Q10
Finding|Gene or Genome|SIMPLE_SEGMENT|9289,9292|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9300,9304|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9300,9304|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9300,9304|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9300,9304|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|9305,9310|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|9316,9326|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9316,9326|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|9347,9357|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9347,9357|false|false|false|C0257343|tamsulosin|Tamsulosin
Event|Event|SIMPLE_SEGMENT|9376,9385|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9376,9385|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9376,9385|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9376,9385|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9376,9385|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9376,9397|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|9376,9397|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9386,9397|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|9386,9397|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|9386,9397|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|9399,9403|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9399,9403|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9399,9403|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9399,9403|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|9406,9415|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9406,9415|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9406,9415|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9406,9415|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9406,9415|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9406,9425|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9416,9425|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9416,9425|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9416,9425|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9416,9425|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9416,9425|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|9436,9441|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9436,9487|false|false|false|C2732749|Acute on chronic diastolic heart failure|Acute on chronic diastolic congestive heart failure
Finding|Intellectual Product|SIMPLE_SEGMENT|9445,9452|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|9445,9452|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9445,9487|false|false|false|C2711480|Chronic diastolic heart failure|chronic diastolic congestive heart failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9453,9462|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9453,9487|false|false|false|C2183328|diastolic congestive heart failure|diastolic congestive heart failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9463,9487|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9474,9479|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9474,9479|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9474,9479|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9474,9487|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|9480,9487|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|9480,9487|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|9480,9487|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|9480,9487|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9488,9491|false|false|false|C0018787|Heart|Cor
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|9488,9491|false|false|false|C0056331|cordycepin|Cor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9488,9491|false|false|false|C0056331|cordycepin|Cor
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9488,9501|false|false|false|C0034072;C0238074|Chronic pulmonary heart disease;Cor pulmonale|Cor pulmonale
Event|Event|SIMPLE_SEGMENT|9492,9501|false|false|false|||pulmonale
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9503,9512|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|9503,9512|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|9503,9512|false|false|false|C1522484|metastatic qualifier|Secondary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9514,9523|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9514,9523|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|9514,9523|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|9514,9536|false|false|false|C0020542|Pulmonary Hypertension|Pulmonary hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9524,9536|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|9524,9536|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9537,9567|false|false|false|C0235480|Paroxysmal atrial fibrillation|Paroxysmal atrial fibrillation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9548,9554|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9548,9567|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9548,9567|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9548,9567|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9555,9567|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|9555,9567|false|false|false|||fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9568,9580|false|false|false|C0020625|Hyponatremia|Hyponatremia
Event|Event|SIMPLE_SEGMENT|9568,9580|false|false|false|||Hyponatremia
Event|Event|SIMPLE_SEGMENT|9584,9593|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9584,9593|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9584,9593|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9584,9593|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9584,9593|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9594,9603|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9594,9603|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9594,9603|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9594,9603|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9605,9611|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9605,9618|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9605,9618|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9612,9618|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9612,9618|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9620,9625|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9620,9625|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|9630,9638|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|9630,9638|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|9640,9645|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9640,9662|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9640,9662|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9649,9662|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9649,9662|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9649,9662|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9664,9669|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|9664,9669|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9664,9669|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|9664,9669|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|9664,9669|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|9664,9669|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|9664,9669|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|9674,9685|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|9674,9685|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|9687,9695|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9687,9695|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9687,9695|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9696,9702|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9696,9702|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9696,9702|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9704,9714|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|9704,9714|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9704,9714|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9704,9714|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9704,9714|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9717,9728|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|9717,9728|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|9717,9728|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|9733,9742|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9733,9742|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9733,9742|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9733,9742|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9733,9742|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9733,9755|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9733,9755|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9733,9755|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9743,9755|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9743,9755|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9743,9755|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|9757,9761|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|9781,9793|false|false|false|||hospitalized
Finding|Functional Concept|SIMPLE_SEGMENT|9798,9809|false|false|false|C0205329|Progressive|progressive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9810,9813|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|9810,9822|false|false|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|SIMPLE_SEGMENT|9814,9822|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|9814,9822|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|9814,9822|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Intellectual Product|SIMPLE_SEGMENT|9838,9842|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|9859,9866|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|9876,9879|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|9876,9879|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9880,9890|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9880,9890|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9880,9890|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9909,9913|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|9914,9921|false|false|false|||prevent
Event|Event|SIMPLE_SEGMENT|9966,9975|false|false|false|||concerned
Drug|Organic Chemical|SIMPLE_SEGMENT|9984,9988|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9984,9988|false|false|false|C0009074|clotrimazole|clot
Event|Event|SIMPLE_SEGMENT|9984,9988|false|false|false|||clot
Finding|Pathologic Function|SIMPLE_SEGMENT|9984,9988|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9997,10002|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|10012,10017|true|false|false|||scans
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10012,10017|true|false|false|C0441633|Scanning|scans
Event|Event|SIMPLE_SEGMENT|10018,10024|true|false|false|||showed
Drug|Organic Chemical|SIMPLE_SEGMENT|10029,10033|true|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10029,10033|true|false|false|C0009074|clotrimazole|clot
Event|Event|SIMPLE_SEGMENT|10029,10033|true|false|false|||clot
Finding|Pathologic Function|SIMPLE_SEGMENT|10029,10033|true|false|false|C0302148|Blood Clot|clot
Finding|Intellectual Product|SIMPLE_SEGMENT|10046,10050|false|false|false|C0282425|News (Publication Type)|news
Event|Event|SIMPLE_SEGMENT|10061,10071|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|10072,10076|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10072,10076|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10072,10076|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10072,10076|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10082,10085|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10082,10085|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10082,10085|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10082,10085|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|10082,10085|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10082,10085|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|10082,10085|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10082,10085|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|10082,10085|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|10082,10085|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|10082,10085|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Anatomy|Body System|SIMPLE_SEGMENT|10091,10101|false|false|false|C0007226|Cardiovascular system|cardiology
Finding|Functional Concept|SIMPLE_SEGMENT|10102,10108|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|10102,10108|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|10102,10111|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|10102,10111|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|10109,10111|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|10121,10129|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|10133,10137|false|false|false|||take
Drug|Organic Chemical|SIMPLE_SEGMENT|10143,10152|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10143,10152|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|10143,10152|false|false|false|||torsemide
Event|Activity|SIMPLE_SEGMENT|10156,10161|false|false|false|C1705178|Order (action)|order
Finding|Classification|SIMPLE_SEGMENT|10156,10161|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Idea or Concept|SIMPLE_SEGMENT|10156,10161|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Intellectual Product|SIMPLE_SEGMENT|10156,10161|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10156,10161|false|false|false|C1373200|Order [PK]|order
Event|Event|SIMPLE_SEGMENT|10165,10173|false|false|false|||maintain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10180,10186|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|10180,10186|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|10180,10186|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|10180,10186|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|10180,10186|false|false|false|C1305866|Weighing patient|weight
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10195,10201|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|10195,10201|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|10195,10201|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|10195,10201|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|10195,10201|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|10224,10228|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|10235,10247|false|false|false|||cardiologist
Finding|Finding|SIMPLE_SEGMENT|10255,10269|false|false|false|C0005911|Body Weight Changes|weight changes
Event|Event|SIMPLE_SEGMENT|10262,10269|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|10262,10269|false|false|false|C0392747|Changing|changes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10303,10312|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10303,10312|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10303,10312|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10303,10325|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10313,10325|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|10313,10325|false|false|false|||hypertension
Event|Event|SIMPLE_SEGMENT|10341,10344|false|false|false|||due
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10365,10369|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10365,10369|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10365,10369|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|10365,10369|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10365,10377|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10370,10377|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10370,10377|false|false|false|||disease
Drug|Organic Chemical|SIMPLE_SEGMENT|10379,10389|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10379,10389|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|10379,10389|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10379,10389|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Event|Event|SIMPLE_SEGMENT|10399,10404|false|false|false|||cause
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10405,10409|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10405,10409|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10405,10409|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|10405,10409|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|10410,10417|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|10410,10417|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|10426,10435|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|10436,10445|false|false|false|||following
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10458,10462|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10458,10462|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10458,10462|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|10458,10462|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|10463,10470|false|false|false|||doctors
Event|Event|SIMPLE_SEGMENT|10479,10489|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|10479,10489|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|10479,10489|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|10493,10496|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|10512,10524|false|false|false|||contributing
Event|Event|SIMPLE_SEGMENT|10537,10545|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|10537,10545|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|10537,10545|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|10553,10557|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10553,10557|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10553,10557|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10553,10557|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10553,10560|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|SIMPLE_SEGMENT|10582,10590|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10591,10603|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10591,10603|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10591,10603|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

