 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
PODIATRY|156,164
<EOL>|164,165
<EOL>|166,167
Patient|179,186
recorded|187,195
as|196,198
having|199,205
No|206,208
Known|209,214
Allergies|215,224
to|225,227
Drugs|228,233
<EOL>|233,234
<EOL>|235,236
Attending|236,245
:|245,246
_|247,248
_|248,249
_|249,250
.|250,251
<EOL>|251,252
<EOL>|253,254
L|271,272
posterior|273,282
tibial|283,289
tendonitis|290,300
/|300,301
tear|301,305
<EOL>|305,306
L|306,307
tarsal|308,314
tunnel|315,321
release|322,329
<EOL>|329,330
<EOL>|331,332
Major|332,337
Surgical|338,346
or|347,349
Invasive|350,358
Procedure|359,368
:|368,369
<EOL>|369,370
L|370,371
_|372,373
_|373,374
_|374,375
tendon|376,382
repair|383,389
<EOL>|389,390
L|390,391
tarsal|392,398
tunnel|399,405
release|406,413
<EOL>|413,414
<EOL>|414,415
<EOL>|416,417
_|445,446
_|446,447
_|447,448
with|449,453
DM|454,456
,|456,457
CAD|458,461
,|461,462
HTN|463,466
admitted|467,475
post-operatively|476,492
following|493,502
<EOL>|502,503
correction|503,513
of|514,516
her|517,520
left|521,525
posterior|526,535
tibial|536,542
tendon|543,549
and|550,553
a|554,555
tarsal|556,562
<EOL>|562,563
tunnel|563,569
release|570,577
.|577,578
Pt|580,582
has|583,586
had|587,590
pain|591,595
in|596,598
her|599,602
left|603,607
foot|608,612
for|613,616
quite|617,622
some|623,627
<EOL>|627,628
time|628,632
,|632,633
an|634,636
MRI|637,640
revealed|641,649
a|650,651
possible|652,660
tear|661,665
,|665,666
intra-operatively|667,684
there|685,690
<EOL>|690,691
was|691,694
a|695,696
large|697,702
posterior|703,712
tear|713,717
to|718,720
the|721,724
_|725,726
_|726,727
_|727,728
tendon|729,735
.|735,736
Also|738,742
,|742,743
a|744,745
tarsal|746,752
<EOL>|752,753
tunnel|753,759
release|760,767
was|768,771
done|772,776
and|777,780
scar|781,785
tissue|786,792
removed|793,800
along|801,806
the|807,810
tibial|811,817
<EOL>|817,818
nerve|818,823
.|823,824
Pt|826,828
has|829,832
a|833,834
history|835,842
of|843,845
pulmonary|846,855
issues|856,862
,|862,863
will|864,868
want|869,873
to|874,876
<EOL>|876,877
observe|877,884
patient|885,892
post-operatively|893,909
as|910,912
she|913,916
underwent|917,926
GA|927,929
to|930,932
make|933,937
<EOL>|938,939
sure|939,943
<EOL>|943,944
she|944,947
does|948,952
not|953,956
have|957,961
problems|962,970
.|970,971
<EOL>|973,974
<EOL>|974,975
<EOL>|976,977
asthma|999,1005
,|1005,1006
emphysema|1007,1016
,|1016,1017
chronic|1018,1025
bronchitis|1026,1036
,|1036,1037
HTN|1038,1041
,|1041,1042
CAD|1043,1046
(|1047,1048
MIx2|1048,1052
,|1052,1053
2|1054,1055
<EOL>|1055,1056
cardiac|1056,1063
stents|1064,1070
_|1071,1072
_|1072,1073
_|1073,1074
,|1074,1075
migraines|1076,1085
,|1085,1086
GERD|1087,1091
,|1091,1092
DM|1093,1095
(|1096,1097
takes|1097,1102
pills|1103,1108
and|1109,1112
<EOL>|1112,1113
insulin|1113,1120
)|1120,1121
,|1121,1122
Anemia|1123,1129
,|1129,1130
neuropathy|1131,1141
,|1141,1142
anxiety|1143,1150
<EOL>|1150,1151
<EOL>|1151,1152
<EOL>|1153,1154
:|1168,1169
<EOL>|1169,1170
_|1170,1171
_|1171,1172
_|1172,1173
<EOL>|1173,1174
:|1188,1189
<EOL>|1189,1190
parents|1190,1197
not|1198,1201
known|1202,1207
.|1207,1208
daughter|1209,1217
htn|1218,1221
<EOL>|1223,1224
<EOL>|1224,1225
<EOL>|1226,1227
Physical|1227,1235
_|1236,1237
_|1237,1238
_|1238,1239
:|1239,1240
<EOL>|1240,1241
Appearance|1241,1251
:|1251,1252
NAD|1253,1256
<EOL>|1256,1257
HEENT|1257,1262
:|1262,1263
PERLA|1264,1269
<EOL>|1269,1270
Heart|1270,1275
:|1275,1276
RRR|1277,1280
<EOL>|1280,1281
Lungs|1281,1286
:|1286,1287
faint|1288,1293
wheezes|1294,1301
otherwise|1302,1311
clear|1312,1317
<EOL>|1317,1318
Abdomen|1318,1325
:|1325,1326
obese|1327,1332
,|1332,1333
NT|1334,1336
/|1336,1337
ND|1337,1339
<EOL>|1339,1340
VASCULAR|1340,1348
<EOL>|1348,1349
Pedal|1349,1354
Pulses|1355,1361
:|1361,1362
[|1368,1369
x|1369,1370
]|1370,1371
Palpable|1372,1380
[|1382,1383
]|1383,1384
Non-palpable|1385,1397
<EOL>|1397,1398
Sub-Papillary|1398,1411
VFT|1412,1415
:|1415,1416
[|1417,1418
x|1418,1419
]|1419,1420
<|1421,1422
3|1423,1424
sec|1425,1428
.|1428,1429
[|1431,1432
]|1432,1433
>|1434,1435
3|1436,1437
sec|1438,1441
.|1441,1442
[|1443,1444
]|1444,1445
Immediate|1446,1455
<EOL>|1455,1456
NEUROLOGICAL|1456,1468
Sensation|1475,1484
:|1484,1485
[|1491,1492
x|1492,1493
]|1493,1494
Intact|1495,1501
[|1503,1504
]|1504,1505
Absent|1506,1512
<EOL>|1512,1513
Proprioception|1532,1546
:|1546,1547
[|1548,1549
]|1549,1550
Intact|1551,1557
[|1559,1560
x|1560,1561
]|1561,1562
Absent|1563,1569
<EOL>|1569,1570
<EOL>|1570,1571
<EOL>|1572,1573
Pertinent|1573,1582
Results|1583,1590
:|1590,1591
<EOL>|1591,1592
Admission|1592,1601
Labs|1602,1606
:|1606,1607
<EOL>|1607,1608
_|1608,1609
_|1609,1610
_|1610,1611
02|1612,1614
:|1614,1615
07PM|1615,1619
BLOOD|1620,1625
WBC|1626,1629
-|1629,1630
9.6|1630,1633
RBC|1634,1637
-|1637,1638
3|1638,1639
.|1639,1640
64|1640,1642
*|1642,1643
Hgb|1644,1647
-|1647,1648
12.3|1648,1652
Hct|1653,1656
-|1656,1657
33|1657,1659
.|1659,1660
1|1660,1661
*|1661,1662
<EOL>|1663,1664
MCV|1664,1667
-|1667,1668
91|1668,1670
MCH|1671,1674
-|1674,1675
33|1675,1677
.|1677,1678
7|1678,1679
*|1679,1680
MCHC|1681,1685
-|1685,1686
37|1686,1688
.|1688,1689
0|1689,1690
*|1690,1691
#|1691,1692
RDW|1693,1696
-|1696,1697
12.9|1697,1701
Plt|1702,1705
_|1706,1707
_|1707,1708
_|1708,1709
<EOL>|1709,1710
_|1710,1711
_|1711,1712
_|1712,1713
11|1714,1716
:|1716,1717
10AM|1717,1721
BLOOD|1722,1727
UreaN|1728,1733
-|1733,1734
15|1734,1736
Creat|1737,1742
-|1742,1743
0.7|1743,1746
Na|1747,1749
-|1749,1750
140|1750,1753
K|1754,1755
-|1755,1756
3.7|1756,1759
Cl|1760,1762
-|1762,1763
98|1763,1765
<EOL>|1766,1767
HCO3|1767,1771
-|1771,1772
28|1772,1774
AnGap|1775,1780
-|1780,1781
18|1781,1783
<EOL>|1783,1784
_|1784,1785
_|1785,1786
_|1786,1787
11|1788,1790
:|1790,1791
10AM|1791,1795
BLOOD|1796,1801
ALT|1802,1805
-|1805,1806
17|1806,1808
AST|1809,1812
-|1812,1813
19|1813,1815
<EOL>|1815,1816
_|1816,1817
_|1817,1818
_|1818,1819
11|1820,1822
:|1822,1823
10AM|1823,1827
BLOOD|1828,1833
Cholest|1834,1841
-|1841,1842
187|1842,1845
<EOL>|1845,1846
_|1846,1847
_|1847,1848
_|1848,1849
11|1850,1852
:|1852,1853
10AM|1853,1857
BLOOD|1858,1863
%|1864,1865
HbA1c|1865,1870
-|1870,1871
10|1871,1873
.|1873,1874
0|1874,1875
*|1875,1876
<EOL>|1876,1877
_|1877,1878
_|1878,1879
_|1879,1880
11|1881,1883
:|1883,1884
10AM|1884,1888
BLOOD|1889,1894
Triglyc|1895,1902
-|1902,1903
185|1903,1906
*|1906,1907
HDL|1908,1911
-|1911,1912
54|1912,1914
CHOL|1915,1919
/|1919,1920
HD|1920,1922
-|1922,1923
3.5|1923,1926
<EOL>|1927,1928
LDLcalc|1928,1935
-|1935,1936
96|1936,1938
<EOL>|1938,1939
<EOL>|1939,1940
<EOL>|1941,1942
The|1965,1968
patient|1969,1976
was|1977,1980
admitted|1981,1989
post-operatively|1990,2006
for|2007,2010
L|2011,2012
_|2013,2014
_|2014,2015
_|2015,2016
repair|2017,2023
and|2024,2027
L|2028,2029
<EOL>|2030,2031
tarsal|2031,2037
tunnel|2038,2044
release|2045,2052
.|2052,2053
The|2055,2058
patient|2059,2066
was|2067,2070
placed|2071,2077
in|2078,2080
a|2081,2082
BK|2083,2085
cast|2086,2090
<EOL>|2091,2092
following|2092,2101
the|2102,2105
completion|2106,2116
of|2117,2119
the|2120,2123
case|2124,2128
.|2128,2129
The|2131,2134
patient|2135,2142
tolerated|2143,2152
the|2153,2156
<EOL>|2157,2158
procedure|2158,2167
and|2168,2171
anesthesia|2172,2182
well|2183,2187
without|2188,2195
apparent|2196,2204
complications|2205,2218
<EOL>|2219,2220
(|2220,2221
see|2221,2224
op|2225,2227
report|2228,2234
for|2235,2238
full|2239,2243
details|2244,2251
)|2251,2252
.|2252,2253
On|2255,2257
POD1|2258,2262
Pt|2263,2265
given|2266,2271
25mg|2272,2276
PO|2277,2279
<EOL>|2280,2281
benadryl|2281,2289
for|2290,2293
RUE|2294,2297
rash|2298,2302
and|2303,2306
shortly|2307,2314
after|2315,2320
,|2320,2321
Pt|2322,2324
triggered|2325,2334
for|2335,2338
<EOL>|2339,2340
hypotension|2340,2351
with|2352,2356
SBP|2357,2360
into|2361,2365
80's|2366,2370
.|2370,2371
Pt|2373,2375
asymptomatic|2376,2388
with|2389,2393
other|2394,2399
<EOL>|2400,2401
vital|2401,2406
signs|2407,2412
stable|2413,2419
,|2419,2420
saturating|2421,2431
well|2432,2436
on|2437,2439
room|2440,2444
air|2445,2448
.|2448,2449
Pt|2451,2453
given|2454,2459
<EOL>|2460,2461
several|2461,2468
500cc|2469,2474
boluses|2475,2482
of|2483,2485
NS|2486,2488
with|2489,2493
return|2494,2500
to|2501,2503
normal|2504,2510
pressures|2511,2520
of|2521,2523
<EOL>|2524,2525
110's|2525,2530
systolic|2531,2539
.|2539,2540
Effects|2542,2549
of|2550,2552
Benadryl|2553,2561
likely|2562,2568
exacerbated|2569,2580
by|2581,2583
Pt|2584,2586
<EOL>|2587,2588
concomitantly|2588,2601
on|2602,2604
narcotics|2605,2614
for|2615,2618
LLE|2619,2622
surgery|2623,2630
.|2630,2631
<EOL>|2633,2634
.|2634,2635
<EOL>|2635,2636
The|2636,2639
patient|2640,2647
was|2648,2651
seen|2652,2656
by|2657,2659
_|2660,2661
_|2661,2662
_|2662,2663
for|2664,2667
NWB|2668,2671
status|2672,2678
and|2679,2682
was|2683,2686
cleared|2687,2694
for|2695,2698
<EOL>|2699,2700
discharge|2700,2709
home|2710,2714
.|2714,2715
The|2716,2719
patient|2720,2727
's|2727,2729
LLE|2730,2733
cast|2734,2738
was|2739,2742
bivalved|2743,2751
and|2752,2755
wrapped|2756,2763
<EOL>|2764,2765
in|2765,2767
ACE|2768,2771
.|2771,2772
The|2773,2776
patient|2777,2784
was|2785,2788
given|2789,2794
strict|2795,2801
instructions|2802,2814
for|2815,2818
_|2819,2820
_|2820,2821
_|2821,2822
LLE|2823,2826
.|2826,2827
<EOL>|2828,2829
Please|2829,2835
see|2836,2839
discharge|2840,2849
intructions|2850,2861
for|2862,2865
full|2866,2870
details|2871,2878
.|2878,2879
<EOL>|2879,2880
.|2880,2881
<EOL>|2881,2882
Advised|2882,2889
to|2890,2892
follow|2893,2899
up|2900,2902
with|2903,2907
Dr.|2908,2911
_|2912,2913
_|2913,2914
_|2914,2915
.|2915,2916
<EOL>|2916,2917
.|2917,2918
<EOL>|2918,2919
Discharged|2919,2929
in|2930,2932
good|2933,2937
condition|2938,2947
with|2948,2952
VSS|2953,2956
.|2956,2957
<EOL>|2957,2958
<EOL>|2958,2959
<EOL>|2960,2961
Medications|2961,2972
on|2973,2975
Admission|2976,2985
:|2985,2986
<EOL>|2986,2987
Advair250|2987,2996
/|2996,2997
50|2997,2999
daily|3000,3005
,|3005,3006
Albuterol|3007,3016
Aerosol|3017,3024
prn|3025,3028
,|3028,3029
EC|3030,3032
ASA|3033,3036
,|3036,3037
Atenolol|3038,3046
100|3047,3050
<EOL>|3051,3052
Insulin|3052,3059
levimir|3060,3067
30|3068,3070
units|3071,3076
AM|3077,3079
;|3079,3080
60|3081,3083
units|3084,3089
_|3090,3091
_|3091,3092
_|3092,3093
,|3093,3094
Isosorbide|3095,3105
Mononitrate|3106,3117
<EOL>|3118,3119
120|3119,3122
,|3122,3123
<EOL>|3123,3124
Lisinopril|3124,3134
10|3135,3137
,|3137,3138
Metformin|3139,3148
[|3149,3150
Glucophage|3150,3160
]|3160,3161
500|3162,3165
mg|3166,3168
TID|3169,3172
,|3172,3173
Nitroglycerin|3174,3187
<EOL>|3188,3189
SL|3189,3191
,|3191,3192
Omeprazole|3193,3203
40|3204,3206
mg|3207,3209
daily|3210,3215
,|3215,3216
Plavix|3217,3223
75|3224,3226
mg|3227,3229
daily|3230,3235
,|3235,3236
Potassium|3237,3246
<EOL>|3247,3248
chloride|3248,3256
20|3258,3260
mEq|3261,3264
,|3264,3265
Simvastatin|3266,3277
80|3278,3280
mg|3281,3283
<EOL>|3283,3284
<EOL>|3285,3286
Discharge|3286,3295
Medications|3296,3307
:|3307,3308
<EOL>|3308,3309
1.|3309,3311
Albuterol|3312,3321
90|3322,3324
mcg|3325,3328
/|3328,3329
Actuation|3329,3338
Aerosol|3339,3346
Sig|3347,3350
:|3350,3351
_|3352,3353
_|3353,3354
_|3354,3355
Puffs|3356,3361
Inhalation|3362,3372
<EOL>|3373,3374
Q4H|3374,3377
(|3378,3379
every|3379,3384
4|3385,3386
hours|3387,3392
)|3392,3393
as|3394,3396
needed|3397,3403
for|3404,3407
wheeze|3408,3414
.|3414,3415
<EOL>|3417,3418
2.|3418,3420
Aspirin|3421,3428
325|3429,3432
mg|3433,3435
Tablet|3436,3442
,|3442,3443
Delayed|3444,3451
Release|3452,3459
(|3460,3461
E.C|3461,3464
.|3464,3465
)|3465,3466
Sig|3467,3470
:|3470,3471
One|3472,3475
(|3476,3477
1|3477,3478
)|3478,3479
<EOL>|3480,3481
Tablet|3481,3487
,|3487,3488
Delayed|3489,3496
Release|3497,3504
(|3505,3506
E.C|3506,3509
.|3509,3510
)|3510,3511
PO|3512,3514
DAILY|3515,3520
(|3521,3522
Daily|3522,3527
)|3527,3528
.|3528,3529
<EOL>|3531,3532
3.|3532,3534
Atenolol|3535,3543
50|3544,3546
mg|3547,3549
Tablet|3550,3556
Sig|3557,3560
:|3560,3561
Two|3562,3565
(|3566,3567
2|3567,3568
)|3568,3569
Tablet|3570,3576
PO|3577,3579
DAILY|3580,3585
(|3586,3587
Daily|3587,3592
)|3592,3593
.|3593,3594
<EOL>|3596,3597
4.|3597,3599
Isosorbide|3600,3610
Mononitrate|3611,3622
60|3623,3625
mg|3626,3628
Tablet|3629,3635
Sustained|3636,3645
Release|3646,3653
24|3654,3656
hr|3657,3659
<EOL>|3660,3661
Sig|3661,3664
:|3664,3665
Two|3666,3669
(|3670,3671
2|3671,3672
)|3672,3673
Tablet|3674,3680
Sustained|3681,3690
Release|3691,3698
24|3699,3701
hr|3702,3704
PO|3705,3707
DAILY|3708,3713
(|3714,3715
Daily|3715,3720
)|3720,3721
.|3721,3722
<EOL>|3724,3725
5.|3725,3727
Lisinopril|3728,3738
10|3739,3741
mg|3742,3744
Tablet|3745,3751
Sig|3752,3755
:|3755,3756
One|3757,3760
(|3761,3762
1|3762,3763
)|3763,3764
Tablet|3765,3771
PO|3772,3774
DAILY|3775,3780
(|3781,3782
Daily|3782,3787
)|3787,3788
.|3788,3789
<EOL>|3790,3791
<EOL>|3792,3793
6.|3793,3795
Metformin|3796,3805
500|3806,3809
mg|3810,3812
Tablet|3813,3819
Sig|3820,3823
:|3823,3824
One|3825,3828
(|3829,3830
1|3830,3831
)|3831,3832
Tablet|3833,3839
PO|3840,3842
TID|3843,3846
(|3847,3848
3|3848,3849
times|3850,3855
a|3856,3857
<EOL>|3858,3859
day|3859,3862
)|3862,3863
.|3863,3864
<EOL>|3866,3867
7.|3867,3869
Nitroglycerin|3870,3883
0.3|3884,3887
mg|3888,3890
Tablet|3891,3897
,|3897,3898
Sublingual|3899,3909
Sig|3910,3913
:|3913,3914
One|3915,3918
(|3919,3920
1|3920,3921
)|3921,3922
Tablet|3923,3929
,|3929,3930
<EOL>|3931,3932
Sublingual|3932,3942
Sublingual|3943,3953
PRN|3954,3957
(|3958,3959
as|3959,3961
needed|3962,3968
)|3968,3969
.|3969,3970
<EOL>|3972,3973
8.|3973,3975
Omeprazole|3976,3986
20|3987,3989
mg|3990,3992
Capsule|3993,4000
,|4000,4001
Delayed|4002,4009
Release|4010,4017
(|4017,4018
E.C|4018,4021
.|4021,4022
)|4022,4023
Sig|4024,4027
:|4027,4028
Two|4029,4032
(|4033,4034
2|4034,4035
)|4035,4036
<EOL>|4037,4038
Capsule|4038,4045
,|4045,4046
Delayed|4047,4054
Release|4055,4062
(|4062,4063
E.C|4063,4066
.|4066,4067
)|4067,4068
PO|4069,4071
DAILY|4072,4077
(|4078,4079
Daily|4079,4084
)|4084,4085
.|4085,4086
<EOL>|4088,4089
9.|4089,4091
Clopidogrel|4092,4103
75|4104,4106
mg|4107,4109
Tablet|4110,4116
Sig|4117,4120
:|4120,4121
One|4122,4125
(|4126,4127
1|4127,4128
)|4128,4129
Tablet|4130,4136
PO|4137,4139
DAILY|4140,4145
<EOL>|4146,4147
(|4147,4148
Daily|4148,4153
)|4153,4154
.|4154,4155
<EOL>|4157,4158
10.|4158,4161
Potassium|4162,4171
Chloride|4172,4180
20|4181,4183
mEq|4184,4187
Tab|4188,4191
Sust|4192,4196
.|4196,4197
Rel|4197,4200
.|4200,4201
Particle|4202,4210
/|4210,4211
Crystal|4211,4218
<EOL>|4219,4220
Sig|4220,4223
:|4223,4224
One|4225,4228
(|4229,4230
1|4230,4231
)|4231,4232
Tab|4233,4236
Sust|4237,4241
.|4241,4242
Rel|4242,4245
.|4245,4246
Particle|4247,4255
/|4255,4256
Crystal|4256,4263
PO|4264,4266
DAILY|4267,4272
(|4273,4274
Daily|4274,4279
)|4279,4280
.|4280,4281
<EOL>|4283,4284
11|4284,4286
.|4286,4287
Simvastatin|4288,4299
40|4300,4302
mg|4303,4305
Tablet|4306,4312
Sig|4313,4316
:|4316,4317
Two|4318,4321
(|4322,4323
2|4323,4324
)|4324,4325
Tablet|4326,4332
PO|4333,4335
DAILY|4336,4341
<EOL>|4342,4343
(|4343,4344
Daily|4344,4349
)|4349,4350
.|4350,4351
<EOL>|4353,4354
12.|4354,4357
Fluticasone|4358,4369
-|4369,4370
Salmeterol|4370,4380
250|4381,4384
-|4384,4385
50|4385,4387
mcg|4388,4391
/|4391,4392
Dose|4392,4396
Disk|4397,4401
with|4402,4406
Device|4407,4413
Sig|4414,4417
:|4417,4418
<EOL>|4419,4420
One|4420,4423
(|4424,4425
1|4425,4426
)|4426,4427
Disk|4428,4432
with|4433,4437
Device|4438,4444
Inhalation|4445,4455
BID|4456,4459
(|4460,4461
2|4461,4462
times|4463,4468
a|4469,4470
day|4471,4474
)|4474,4475
.|4475,4476
<EOL>|4478,4479
13.|4479,4482
Insulin|4483,4490
<EOL>|4490,4491
levimir|4491,4498
30|4499,4501
units|4502,4507
qAM|4508,4511
and|4512,4515
60|4516,4518
units|4519,4524
qPM|4525,4528
<EOL>|4528,4529
14.|4529,4532
Compazine|4533,4542
10|4543,4545
mg|4546,4548
Tablet|4549,4555
Sig|4556,4559
:|4559,4560
One|4561,4564
(|4565,4566
1|4566,4567
)|4567,4568
Tablet|4569,4575
PO|4576,4578
every|4579,4584
six|4585,4588
(|4589,4590
6|4590,4591
)|4591,4592
<EOL>|4593,4594
hours|4594,4599
as|4600,4602
needed|4603,4609
for|4610,4613
nausea|4614,4620
.|4620,4621
<EOL>|4621,4622
Disp|4622,4626
:|4626,4627
*|4627,4628
30|4628,4630
Tablet|4631,4637
(|4637,4638
s|4638,4639
)|4639,4640
*|4640,4641
Refills|4642,4649
:|4649,4650
*|4650,4651
0|4651,4652
*|4652,4653
<EOL>|4653,4654
15.|4654,4657
Oxycodone|4658,4667
-|4667,4668
Acetaminophen|4668,4681
_|4682,4683
_|4683,4684
_|4684,4685
mg|4686,4688
Tablet|4689,4695
Sig|4696,4699
:|4699,4700
_|4701,4702
_|4702,4703
_|4703,4704
Tablets|4705,4712
PO|4713,4715
<EOL>|4716,4717
Q4H|4717,4720
(|4721,4722
every|4722,4727
4|4728,4729
hours|4730,4735
)|4735,4736
as|4737,4739
needed|4740,4746
for|4747,4750
pain|4751,4755
.|4755,4756
<EOL>|4756,4757
Disp|4757,4761
:|4761,4762
*|4762,4763
50|4763,4765
Tablet|4766,4772
(|4772,4773
s|4773,4774
)|4774,4775
*|4775,4776
Refills|4777,4784
:|4784,4785
*|4785,4786
0|4786,4787
*|4787,4788
<EOL>|4788,4789
16|4789,4791
.|4791,4792
Oxycodone|4793,4802
10|4803,4805
mg|4806,4808
Tablet|4809,4815
Sustained|4816,4825
Release|4826,4833
12|4834,4836
hr|4837,4839
Sig|4840,4843
:|4843,4844
_|4845,4846
_|4846,4847
_|4847,4848
<EOL>|4849,4850
Tablet|4850,4856
Sustained|4857,4866
Release|4867,4874
12|4875,4877
hrs|4878,4881
PO|4882,4884
Q12H|4885,4889
(|4890,4891
every|4891,4896
12|4897,4899
hours|4900,4905
)|4905,4906
.|4906,4907
<EOL>|4907,4908
Disp|4908,4912
:|4912,4913
*|4913,4914
40|4914,4916
Tablet|4917,4923
Sustained|4924,4933
Release|4934,4941
12|4942,4944
hr|4945,4947
(|4947,4948
s|4948,4949
)|4949,4950
*|4950,4951
Refills|4952,4959
:|4959,4960
*|4960,4961
1|4961,4962
*|4962,4963
<EOL>|4963,4964
17.|4964,4967
Docusate|4968,4976
Sodium|4977,4983
100|4984,4987
mg|4988,4990
Tablet|4991,4997
Sig|4998,5001
:|5001,5002
Two|5003,5006
(|5007,5008
2|5008,5009
)|5009,5010
Tablet|5011,5017
PO|5018,5020
twice|5021,5026
a|5027,5028
<EOL>|5029,5030
day|5030,5033
.|5033,5034
<EOL>|5034,5035
Disp|5035,5039
:|5039,5040
*|5040,5041
60|5041,5043
Tablet|5044,5050
(|5050,5051
s|5051,5052
)|5052,5053
*|5053,5054
Refills|5055,5062
:|5062,5063
*|5063,5064
2|5064,5065
*|5065,5066
<EOL>|5066,5067
<EOL>|5067,5068
<EOL>|5069,5070
Discharge|5070,5079
Disposition|5080,5091
:|5091,5092
<EOL>|5092,5093
Home|5093,5097
<EOL>|5097,5098
<EOL>|5099,5100
Discharge|5100,5109
Diagnosis|5110,5119
:|5119,5120
<EOL>|5120,5121
Left|5121,5125
posterior|5126,5135
tibialis|5136,5144
tendonitis|5145,5155
<EOL>|5155,5156
Left|5156,5160
tarsal|5161,5167
tunnel|5168,5174
<EOL>|5174,5175
<EOL>|5175,5176
<EOL>|5177,5178
Good|5199,5203
<EOL>|5203,5204
<EOL>|5204,5205
<EOL>|5206,5207
Please|5231,5237
resume|5238,5244
all|5245,5248
pre-admission|5249,5262
medications|5263,5274
.|5274,5275
You|5277,5280
were|5281,5285
given|5286,5291
new|5292,5295
<EOL>|5296,5297
prescriptions|5297,5310
,|5310,5311
please|5312,5318
take|5319,5323
as|5324,5326
directed|5327,5335
.|5335,5336
<EOL>|5336,5337
.|5337,5338
<EOL>|5338,5339
Keep|5339,5343
your|5344,5348
dressing|5349,5357
/|5357,5358
cast|5358,5362
clean|5363,5368
and|5369,5372
dry|5373,5376
at|5377,5379
all|5380,5383
times|5384,5389
.|5389,5390
You|5392,5395
will|5396,5400
<EOL>|5401,5402
not|5402,5405
have|5406,5410
any|5411,5414
dressing|5415,5423
changes|5424,5431
.|5431,5432
<EOL>|5432,5433
.|5433,5434
<EOL>|5434,5435
You|5435,5438
are|5439,5442
to|5443,5445
remain|5446,5452
NON|5453,5456
WEIGHT|5457,5463
BEARING|5464,5471
on|5472,5474
your|5475,5479
left|5480,5484
foot|5485,5489
in|5490,5492
a|5493,5494
cast|5495,5499
<EOL>|5500,5501
with|5501,5505
crutches|5506,5514
/|5514,5515
walker|5515,5521
/|5521,5522
wheelchair|5522,5532
at|5533,5535
all|5536,5539
times|5540,5545
.|5545,5546
Keep|5548,5552
your|5553,5557
left|5558,5562
<EOL>|5563,5564
foot|5564,5568
elevated|5569,5577
to|5578,5580
prevent|5581,5588
swelling|5589,5597
.|5597,5598
<EOL>|5598,5599
.|5599,5600
<EOL>|5600,5601
Call|5601,5605
your|5606,5610
doctor|5611,5617
or|5618,5620
go|5621,5623
to|5624,5626
the|5627,5630
ED|5631,5633
for|5634,5637
any|5638,5641
increase|5642,5650
in|5651,5653
left|5654,5658
foot|5659,5663
<EOL>|5664,5665
redness|5665,5672
,|5672,5673
swelling|5674,5682
or|5683,5685
purulent|5686,5694
drainage|5695,5703
from|5704,5708
your|5709,5713
wound|5714,5719
,|5719,5720
for|5721,5724
any|5725,5728
<EOL>|5729,5730
nausea|5730,5736
,|5736,5737
vomiting|5738,5746
,|5746,5747
fevers|5748,5754
greater|5755,5762
than|5763,5767
101.5|5768,5773
,|5773,5774
chills|5775,5781
,|5781,5782
night|5783,5788
<EOL>|5789,5790
sweats|5790,5796
or|5797,5799
any|5800,5803
worsening|5804,5813
symptoms|5814,5822
.|5822,5823
<EOL>|5823,5824
<EOL>|5825,5826
Followup|5826,5834
Instructions|5835,5847
:|5847,5848
<EOL>|5848,5849
_|5849,5850
_|5850,5851
_|5851,5852
<EOL>|5852,5853

