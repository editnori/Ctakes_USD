CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|tramadol|Drug|false|false||Tramadol
null|tramadol|Drug|false|false||Tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||Tramadolnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Abdomen distended|Finding|false|false||Abdominal distentionnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Distention|Finding|false|false||distention
null|Pathological Dilatation|Finding|false|false||distentionnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Paracentesis|Procedure|false|false||Paracentesisnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Alcohol abuse|Disorder|false|false||ETOH abusenull|ethanol|Drug|false|false||ETOH
null|ethanol|Drug|false|false||ETOHnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Abdomen distended|Finding|false|false||abdominal distentionnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Distention|Finding|false|false||distention
null|Pathological Dilatation|Finding|false|false||distentionnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|Clinic|Device|false|false||Clinic
null|Ambulatory Care Facilities|Device|false|false||Clinicnull|Clinic|Entity|false|false||Clinic
null|Ambulatory Care Facilities|Entity|false|false||Clinicnull|Patient location type - Clinic|Modifier|false|false||Clinic
null|Person location type - Clinic|Modifier|false|false||Clinicnull|Recent|Time|false|false||recentlynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Combined diagnostic and therapeutic intent|Finding|false|false||diagnostic and therapeuticnull|Diagnostic agents|Drug|false|false||diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||diagnostic
null|Diagnostic|Finding|false|false||diagnosticnull|Diagnostic dental procedure|Procedure|false|false||diagnostic
null|Diagnosis|Procedure|false|false||diagnosticnull|Therapeutic abdominal paracentesis|Procedure|false|false||therapeutic paracentesisnull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Paracentesis|Procedure|false|false||paracentesisnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|Clinic|Device|false|false||Clinic
null|Ambulatory Care Facilities|Device|false|false||Clinicnull|Clinic|Entity|false|false||Clinic
null|Ambulatory Care Facilities|Entity|false|false||Clinicnull|Patient location type - Clinic|Modifier|false|false||Clinic
null|Person location type - Clinic|Modifier|false|false||Clinicnull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Presentation|Finding|false|false||presentationnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Fever|Finding|false|false||feversnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Alcohol abuse|Disorder|false|false||Alcohol abusenull|Alcohols|Drug|false|false||Alcohol
null|Alcohols|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||Alcoholnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Chronic back pain|Finding|false|false||Chronic back painnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Malignant neoplasm of breast|Disorder|false|false||Breast cancer
null|Breast Carcinoma|Disorder|false|false||Breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||Breastnull|Breast problem|Finding|false|false||Breastnull|Procedures on breast|Procedure|false|false||Breastnull|Breast|Anatomy|false|false||Breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|ibudilast|Drug|true|false||IBD
null|ibudilast|Drug|true|false||IBDnull|Inflammatory Bowel Diseases|Disorder|true|false||IBD
null|Irritable Bowel Syndrome|Disorder|true|false||IBDnull|ACAD8 wt Allele|Finding|true|false||IBDnull|Liver Failure|Disorder|true|false||liver failurenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Failure (biologic function)|Finding|true|false||failure
null|Failure|Finding|true|false||failure
null|Personal failure|Finding|true|false||failurenull|Numerous|LabModifier|false|false||Multiplenull|Relative (related person)|Subject|false|false||relativesnull|Alcoholic Intoxication, Chronic|Disorder|false|false||alcoholismnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|Pleasant|Finding|false|false||pleasantnull|Appropriate|Modifier|false|false||appropriatenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|HEENT|Anatomy|false|false||HEENTnull|Facial wasting|Disorder|true|false||temporal wastingnull|Temporal wasting|Finding|true|false||temporal wastingnull|Temporal - Temporal Qualifier|Time|false|false||temporalnull|Temporal Anatomic Qualifier|Modifier|false|false||temporalnull|Wasting|Disorder|true|false||wastingnull|Cachexia|Finding|true|false||wastingnull|Jugular venous engorgement|Finding|true|false||JVDnull|Neck>Neck veins|Anatomy|false|false||neck veins
null|Structure of vein of neck|Anatomy|false|false||neck veinsnull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Fill|Event|false|false||fillnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|MAS1L gene|Finding|true|false||MRGnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|cetrimonium bromide|Drug|false|false||CTABnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Dilated|Finding|false|false||Distendednull|Distended|Modifier|false|false||Distendednull|Tights|Device|false|false||tightnull|Tightness sensation quality|Modifier|false|false||tightnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Flatulence|Finding|false|false||flatulencenull|Limb structure|Anatomy|false|false||LIMBSnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Lewis Blood-Group System|Finding|false|false||LEsnull|Inferior esophageal sphincter structure|Anatomy|false|false||LEsnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Asterixis|Finding|true|false||asterixisnull|Very mild|Finding|true|false||very mildnull|Very|Modifier|false|false||verynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||generalnull|General medical service|Procedure|false|false||generalnull|Generalized|Modifier|false|false||generalnull|Tremor|Finding|false|false||tremornull|Laboratory test finding|Lab|false|false||Labsnull|at admission|Finding|false|false||at Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bands|Device|false|false||Bandsnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood ethanol|Procedure|false|false||BLOOD Ethanolnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CNS depressants ethanol|Drug|false|false||Ethanol
null|CNS depressants ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanolnull|Toxic effect of ethyl alcohol|Disorder|false|false||Ethanolnull|Ethanol measurement|Procedure|false|false||Ethanolnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Laboratory test finding|Lab|false|false||Labsnull|At discharge|Time|false|false||at Dischargenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Micro (prefix)|Finding|false|false||Micro
null|Microbiology - Laboratory Class|Finding|false|false||Micronull|Microbiology procedure|Procedure|false|false||Micronull|Unit Of Measure Prefix - micro|LabModifier|false|false||Micronull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|peritoneal fluid Gram stain|Procedure|false|false||PERITONEAL FLUID GRAM STAINnull|Peritoneal fluid (substance)|Finding|true|false||PERITONEAL FLUIDnull|Peritoneal fluid analysis|Procedure|true|false||PERITONEAL FLUIDnull|peritoneal|Anatomy|false|false||PERITONEAL
null|Peritoneum|Anatomy|false|false||PERITONEALnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|true|false||STAINnull|Staining method|Procedure|true|false||STAINnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Pending - Allergy Clinical Status|Finding|false|false||PENDING
null|Pending - referral status|Finding|false|false||PENDINGnull|Pending - status|Time|false|false||PENDINGnull|pending - ManagedParticipationStatus|Modifier|false|false||PENDING
null|pending - RoleStatus|Modifier|false|false||PENDING
null|Pending - Day type|Modifier|false|false||PENDINGnull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Feces|Finding|false|false||STOOLnull|Stool seat|Device|false|false||STOOLnull|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN Anull|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXINnull|Clostridioides difficile|Entity|false|false||CLOSTRIDIUM DIFFICILEnull|Genus Clostridium (organism)|Entity|false|false||CLOSTRIDIUMnull|Toxin|Drug|false|false||TOXIN
null|Toxin|Drug|false|false||TOXINnull|Toxin (disposition)|Modifier|false|false||TOXINnull|Tests (qualifier value)|Finding|false|false||TEST
null|Testing|Finding|false|false||TESTnull|Laboratory Procedures|Procedure|false|false||TESTnull|Test - temporal region|Anatomy|false|false||TESTnull|Test Result|Lab|false|false||TESTnull|Test Dosing Unit|LabModifier|false|false||TESTnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Swab Dosage Form|Drug|false|false||SWAB
null|Swab specimen|Drug|false|false||SWABnull|Taking of swab|Procedure|false|false||SWABnull|Swab|Device|false|false||SWABnull|Swab Dosing Unit|LabModifier|false|false||SWABnull|Vancomycin-Resistant Enterococci|Entity|false|false||VANCOMYCIN RESISTANT ENTEROCOCCUSnull|vancomycin|Drug|false|false||VANCOMYCIN
null|vancomycin|Drug|false|false||VANCOMYCINnull|Vancomycin measurement|Procedure|false|false||VANCOMYCINnull|resistant - Observation Interpretation Susceptibility|Finding|false|false||RESISTANT
null|Resistant (qualifier value)|Finding|false|false||RESISTANTnull|Antimicrobial Resistance Result|Lab|false|false||RESISTANTnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Feces|Finding|false|false||STOOLnull|Stool seat|Device|false|false||STOOLnull|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN Anull|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXINnull|Clostridioides difficile|Entity|false|false||CLOSTRIDIUM DIFFICILEnull|Genus Clostridium (organism)|Entity|false|false||CLOSTRIDIUMnull|Toxin|Drug|false|false||TOXIN
null|Toxin|Drug|false|false||TOXINnull|Toxin (disposition)|Modifier|false|false||TOXINnull|Tests (qualifier value)|Finding|false|false||TEST
null|Testing|Finding|false|false||TESTnull|Laboratory Procedures|Procedure|false|false||TESTnull|Test - temporal region|Anatomy|false|false||TESTnull|Test Result|Lab|false|false||TESTnull|Test Dosing Unit|LabModifier|false|false||TESTnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|In Blood|Finding|false|false||IN BLOODnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|In Blood|Finding|false|false||BLOOD
null|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOODnull|Culture Bottles|Device|false|false||CULTURE BOTTLESnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|null|Device|false|false||BOTTLESnull|Bottle Dosing Unit|LabModifier|false|false||BOTTLESnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|null|Device|false|false||Bottlesnull|Bottle Dosing Unit|LabModifier|false|false||Bottlesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|peritoneal fluid Gram stain|Procedure|false|false||PERITONEAL FLUID GRAM STAINnull|Peritoneal fluid (substance)|Finding|false|false||PERITONEAL FLUIDnull|Peritoneal fluid analysis|Procedure|false|false||PERITONEAL FLUIDnull|peritoneal|Anatomy|false|false||PERITONEAL
null|Peritoneum|Anatomy|false|false||PERITONEALnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood culture|Procedure|false|false||CULTURE Bloodnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood culture|Procedure|false|false||CULTURE Bloodnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|gram|LabModifier|false|false||GRAMnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|bacteria aspects|Finding|false|false||BACTERIAnull|Bacteria <walking sticks>|Entity|false|false||BACTERIA
null|Bacteria|Entity|false|false||BACTERIAnull|Referral category - Inpatient|Finding|false|false||INPATIENT
null|Patient Class - Inpatient|Finding|false|false||INPATIENTnull|inpatient encounter|Procedure|false|false||INPATIENTnull|inpatient|Subject|false|false||INPATIENTnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|In Blood|Finding|false|false||IN BLOODnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|In Blood|Finding|false|false||BLOOD
null|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOODnull|Culture Bottles|Device|false|false||CULTURE BOTTLESnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|null|Device|false|false||BOTTLESnull|Bottle Dosing Unit|LabModifier|false|false||BOTTLESnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Pulmonary Embolism|Finding|true|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|true|false||embolism
null|Embolus|Finding|true|false||embolismnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Atelectasis|Finding|false|false||atelectasisnull|Structure of base of right lung|Anatomy|false|false||right lung basenull|Right lung|Anatomy|false|false||right lungnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Basal segment of lung|Anatomy|false|false||lung basenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Small|LabModifier|false|false||smallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Hepatomegaly|Finding|false|false||Hepatomegalynull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hepatic|Anatomy|false|false||portalnull|Venous thrombosis after immobility|Finding|true|false||venous thrombosis
null|Venous Thrombosis|Finding|true|false||venous thrombosisnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|true|false||thrombosisnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|null|Time|false|false||priornull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Extreme|Modifier|false|false||extremelynull|Slow|Modifier|false|false||slownull|Undetectable|Attribute|false|false||undetectablenull|Flow|Phenomenon|false|false||flownull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Small|LabModifier|false|false||smallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Basilar atelectasis|Finding|false|false||basilar atelectasisnull|Basilar|Modifier|false|false||basilarnull|Atelectasis|Finding|false|false||atelectasisnull|Replaced by|Finding|false|false||Replaced
null|Replacement|Finding|false|false||Replacednull|Structure of right branch of hepatic artery|Anatomy|false|false||right hepatic artery
null|null|Anatomy|false|false||right hepatic arterynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Abdomen>Hepatic artery|Anatomy|false|false||hepatic artery
null|Hepatic artery|Anatomy|false|false||hepatic arterynull|Hepatic|Anatomy|false|false||hepaticnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|SNRPF protein, human|Drug|false|false||SMA
null|SNRPF protein, human|Drug|false|false||SMAnull|Minor Salivary Gland Sclerosing Microcystic Adenocarcinoma|Disorder|false|false||SMA
null|Proximal spinal muscular atrophy|Disorder|false|false||SMA
null|Spinal Muscular Atrophy|Disorder|false|false||SMAnull|SMN1 wt Allele|Finding|false|false||SMA
null|SMN1 gene|Finding|false|false||SMAnull|Southern Sami Language|Entity|false|false||SMAnull|Conventional|Modifier|false|false||conventionalnull|Arteries|Anatomy|false|false||arterialnull|Arterial|Modifier|false|false||arterialnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Anatomical structure|Anatomy|false|false||anatomynull|Science of Anatomy|Title|false|false||anatomynull|Anatomy aspects|Modifier|false|false||anatomynull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Fever|Finding|false|false||feversnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Ascites|Disorder|false|false||ASCITESnull|Peritoneal Effusion|Finding|false|false||ASCITESnull|ALLC gene|Finding|false|false||ALCnull|Absolute Blood Lymphocyte Count|Procedure|false|false||ALCnull|area LC of Bonin|Anatomy|false|false||ALCnull|Hepatitis A|Disorder|false|false||HEPATITIS
null|Hepatitis|Disorder|false|false||HEPATITISnull|Leukocytosis|Disorder|false|false||LEUKOCYTOSISnull|Blood leukocyte number above reference range|Finding|false|false||LEUKOCYTOSISnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Fatty Liver|Disorder|false|false||fatty liver
null|Steatohepatitis|Disorder|false|false||fatty livernull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Extensive|Modifier|false|false||extensivenull|Drinking (function)|Finding|false|false||drinking
null|Alcohol consumption|Finding|false|false||drinkingnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Paracentesis|Procedure|false|false||paracentesisnull|Peritoneal fluid (substance)|Finding|false|false||peritoneal fluidnull|Peritoneal fluid analysis|Procedure|false|false||peritoneal fluidnull|peritoneal|Anatomy|false|false||peritoneal
null|Peritoneum|Anatomy|false|false||peritonealnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Androgen Binding Protein|Drug|true|false||SBP
null|Androgen Binding Protein|Drug|true|false||SBPnull|CCHCR1 wt Allele|Finding|true|false||SBP
null|SHBG wt Allele|Finding|true|false||SBPnull|Systolic blood pressure measurement|Procedure|true|false||SBPnull|Systolic Pressure|Attribute|true|false||SBPnull|Diuretics|Drug|false|false||Diureticsnull|Initially|Time|false|false||initiallynull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Hyponatremia|Disorder|false|false||hyponatremianull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|BRIEF Health Literacy Screening Tool|Finding|false|false||brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|day|Time|false|false||daysnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Paracentesis|Procedure|false|false||paracentesesnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Leukocytes|Anatomy|false|false||white cellnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Cell Count|Procedure|false|false||cell countnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Bilirubin|Drug|false|false||total bilirubin
null|Bilirubin|Drug|false|false||total bilirubinnull|Total bilirubin metabolic function|Finding|false|false||total bilirubinnull|Bilirubin, total measurement|Procedure|false|false||total bilirubinnull|Total bilirubin level|Lab|false|false||total bilirubinnull|Total|Modifier|false|false||totalnull|bilirubin preparation|Drug|false|false||bilirubin
null|bilirubin preparation|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubinnull|Bilirubin, total measurement|Procedure|false|false||bilirubin
null|blood bilirubin level test|Procedure|false|false||bilirubinnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Ambulatory Care Facilities|Device|false|false||clinic
null|Clinic|Device|false|false||clinicnull|Ambulatory Care Facilities|Entity|false|false||clinic
null|Clinic|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Primary Care Provider - Provider role|Finding|false|false||primary care providernull|null|Attribute|false|false||primary care providernull|Primary care provider|Subject|false|false||primary care providernull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|Two weeks|Time|false|false||two weeksnull|week|Time|false|false||weeksnull|Hyponatremia|Disorder|false|false||HYPONATREMIAnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Hypovolemic|Lab|false|false||hypovolemicnull|Hyponatremia|Disorder|false|false||hyponatremianull|Protein Component|Drug|false|false||component
null|Protein Component|Drug|false|false||componentnull|Specimen Child Role - Component|Finding|false|false||component
null|Component (part)|Finding|false|false||component
null|Component, LOINC Axis 1|Finding|false|false||componentnull|Component object|Device|false|false||componentnull|Hyponatremia|Disorder|false|false||hyponatremianull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Discretion|Finding|false|false||discretionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Team|Subject|false|false||teamnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Sodium decreased|Finding|false|false||low sodiumnull|Low sodium diet|Procedure|false|false||low sodiumnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Free water|Drug|false|false||free waternull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Restricted|Finding|false|false||restrictionnull|Daily|Time|false|false||dailynull|Alcoholic Intoxication, Chronic|Disorder|false|false||ALCOHOLISMnull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Recent|Time|false|false||recentlynull|Report (document)|Finding|false|false||reportsnull|Reporting|Procedure|false|false||reportsnull|Daily|Time|false|false||dailynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Alcohol consumption|Finding|false|false||alcohol intakenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|year|Time|false|false||yearsnull|Withdrawal Symptoms|Finding|false|false||withdrawal symptomsnull|Withdrawal (dysfunction)|Disorder|false|false||withdrawalnull|Withdrawal - birth control|Procedure|false|false||withdrawalnull|Withdraw (activity)|Event|false|false||withdrawalnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Seizures|Finding|true|false||seizuresnull|Shakes|Finding|false|false||Shakes
null|Tremor|Finding|false|false||Shakesnull|Hallucinations|Disorder|false|false||hallucinationsnull|Report (document)|Finding|false|false||Reportsnull|Reporting|Procedure|false|false||Reportsnull|sobriety|Finding|false|false||sobrietynull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Urinary tract infection|Disorder|false|false||URINARY TRACT INFECTIONnull|Urinary tract|Anatomy|false|false||URINARY TRACT
null|Urinary system|Anatomy|false|false||URINARY TRACTnull|Urinary tract|Anatomy|false|false||URINARYnull|urinary|Modifier|false|false||URINARYnull|Tract|Anatomy|false|false||TRACTnull|Communicable Diseases|Disorder|false|false||INFECTIONnull|Infection|Finding|false|false||INFECTIONnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Empiric|Modifier|false|false||empiricnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Concern|Finding|false|false||concernnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Back Pain|Finding|false|false||BACK PAINnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Abdominal Pain|Finding|false|false||ABDOMINAL PAINnull|Abdomen|Anatomy|false|false||ABDOMINALnull|Abdominal (qualifier value)|Modifier|false|false||ABDOMINALnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch Dosage Form|Device|false|false||patchesnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Course|Time|false|false||coursenull|tramadol|Drug|false|false||Tramadol
null|tramadol|Drug|false|false||Tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||Tramadolnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Primary Care Provider - Provider role|Finding|false|false||primary care providernull|null|Attribute|false|false||primary care providernull|Primary care provider|Subject|false|false||primary care providernull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|EntityNameUseR2 - temporary|Finding|false|false||temporary
null|Job Status - Temporary|Finding|false|false||temporarynull|Transitory|Time|false|false||temporarynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Acute hepatitis|Disorder|false|false||acute hepatitisnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Prophylactic treatment|Procedure|false|false||Prophylaxisnull|prevention & control|Modifier|false|false||Prophylaxisnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|PPP4C gene|Finding|false|false||ppxnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Bowel Regimen|Procedure|false|false||Bowel regimennull|Intestines|Anatomy|false|false||Bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|lactulose|Drug|false|false||lactulose
null|lactulose|Drug|false|false||lactulosenull|Proton Pump Inhibitors|Drug|true|false||PPInull|Prepulse Inhibition|Finding|true|false||PPInull|Pain management (procedure)|Procedure|false|false||Pain managementnull|Pain Management (specialty)|Title|false|false||Pain managementnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Lidocaine Patch|Drug|false|false||lidocaine patchnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Communication|Finding|false|false||Communicationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||fullnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Thiamine Drug Class|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|thiamine|Drug|false|false||thiamine
null|Thiamine Drug Class|Drug|false|false||thiaminenull|Thiamine measurement|Procedure|false|false||thiaminenull|folate|Drug|false|false||folate
null|folate|Drug|false|false||folate
null|folate|Drug|false|false||folatenull|Folic acid measurement|Procedure|false|false||folatenull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Daily|Time|false|false||dailynull|Lidocaine Patch|Drug|false|false||lidocaine patchnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Nicotine Transdermal Patch|Drug|false|false||nicotine patchnull|nicotine|Drug|false|false||nicotine
null|nicotine|Drug|false|false||nicotinenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Multivitamin tablet|Drug|false|false||Multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HClnull|Thiamine Drug Class|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|Thiamine Drug Class|Drug|false|false||Thiaminenull|Thiamine measurement|Procedure|false|false||Thiaminenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acidnull|Folic acid measurement|Procedure|false|false||Folic Acidnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|nicotine|Drug|false|false||Nicotine
null|nicotine|Drug|false|false||Nicotinenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Transdermal Route of Administration|Finding|false|false||Transdermal
null|transdermal|Finding|false|false||Transdermal
null|Transdermal (intended site)|Finding|false|false||Transdermalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|ADHESIVE PATCH, MEDICATED|Device|false|false||Adhesive Patch, Medicatednull|Adhesives|Device|false|false||Adhesivenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Medicated|Drug|false|false||Medicatednull|Medicated (finding)|Finding|false|false||Medicatednull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|ADHESIVE PATCH, MEDICATED|Device|false|false||Adhesive Patch, Medicatednull|Adhesives|Device|false|false||Adhesivenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Medicated|Drug|false|false||Medicatednull|Medicated (finding)|Finding|false|false||Medicatednull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|tramadol|Drug|false|false||Tramadol
null|tramadol|Drug|false|false||Tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||Tramadolnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary diagnosisnull|Principal diagnosis|Modifier|false|false||Primary diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Hepatitis, Alcoholic|Disorder|false|false||Alcoholic hepatitisnull|Alcoholics|Subject|false|false||Alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Excessive (qualifier value)|Modifier|false|false||excessivenull|Alcohol consumption|Finding|false|false||alcohol intakenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocytes|Anatomy|false|false||white cellnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Cell Count|Procedure|false|false||cell countnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Sometimes|Time|false|false||sometimesnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Behavior Rating Inventory of Executive Function|Finding|false|false||brief
null|BRIEF Health Literacy Screening Tool|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Course|Time|false|false||coursenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Urinary tract infection|Disorder|false|false||urinary tract infectionnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Peritoneal fluid (substance)|Finding|false|false||peritoneal fluidnull|Peritoneal fluid analysis|Procedure|false|false||peritoneal fluidnull|peritoneal|Anatomy|false|false||peritoneal
null|Peritoneum|Anatomy|false|false||peritonealnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Blood sodium|Procedure|false|false||blood sodiumnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Too low|Finding|false|false||too lownull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|tramadol|Drug|false|false||Tramadol
null|tramadol|Drug|false|false||Tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||Tramadolnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions