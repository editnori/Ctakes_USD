 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Chief|210,215
Complaint|216,225
:|225,226
<EOL>|226,227
Back|227,231
Pain|232,236
<EOL>|236,237
<EOL>|238,239
Major|239,244
Surgical|245,253
or|254,256
Invasive|257,265
Procedure|266,275
:|275,276
<EOL>|276,277
None|277,281
<EOL>|281,282
<EOL>|282,283
<EOL>|284,285
History|285,292
of|293,295
Present|296,303
Illness|304,311
:|311,312
<EOL>|312,313
The|313,316
patient|317,324
is|325,327
a|328,329
_|330,331
_|331,332
_|332,333
y|334,335
/|335,336
o|336,337
F|338,339
with|340,344
pMHx|345,349
significant|350,361
for|362,365
HTN|366,369
,|369,370
GERD|371,375
,|375,376
<EOL>|377,378
CAD|378,381
s|382,383
/|383,384
p|384,385
CABG|386,390
and|391,394
stenting|395,403
,|403,404
IDDM|405,409
with|410,414
periperal|415,424
neuropathy|425,435
who|436,439
<EOL>|440,441
presents|441,449
with|450,454
R|455,456
flank|457,462
pain|463,467
.|467,468
<EOL>|470,471
Per|471,474
patient|475,482
,|482,483
this|484,488
pain|489,493
has|494,497
been|498,502
going|503,508
on|509,511
for|512,515
the|516,519
past|520,524
3|525,526
weeks|527,532
<EOL>|533,534
but|534,537
has|538,541
worsened|542,550
over|551,555
the|556,559
past|560,564
2|565,566
days|567,571
.|571,572
It|573,575
is|576,578
worsened|579,587
with|588,592
<EOL>|593,594
coughing|594,602
and|603,606
moving|607,613
.|613,614
She|615,618
otherwise|619,628
denies|629,635
any|636,639
dysuria|640,647
,|647,648
urinary|649,656
<EOL>|657,658
frequency|658,667
,|667,668
abdominal|669,678
pain|679,683
,|683,684
n|685,686
/|686,687
v|687,688
,|688,689
chest|690,695
pain|696,700
,|700,701
shortness|702,711
of|712,714
breath|715,721
<EOL>|722,723
or|723,725
dizziness|726,735
.|735,736
She|737,740
endorses|741,749
4|750,751
episodes|752,760
of|761,763
diarrhea|764,772
today|773,778
.|778,779
<EOL>|781,782
In|782,784
the|785,788
ED|789,791
initial|792,799
vitals|800,806
were|807,811
:|811,812
10|813,815
98.2|816,820
106|821,824
167|825,828
/|828,829
84|829,831
16|832,834
99|835,837
%|837,838
RA|839,841
.|841,842
RR|843,845
<EOL>|846,847
later|847,852
trended|853,860
up|861,863
to|864,866
20|867,869
,|869,870
HR|871,873
down|874,878
to|879,881
89|882,884
.|884,885
Labs|886,890
were|891,895
significant|896,907
for|908,911
<EOL>|912,913
positive|913,921
UA|922,924
(|925,926
WBC|926,929
19|930,932
)|932,933
,|933,934
lactate|935,942
3.0|943,946
,|946,947
WBC|948,951
9.4|952,955
%|955,956
(|957,958
70|958,960
%|960,961
PMN|962,965
)|965,966
,|966,967
AST|968,971
53|972,974
,|974,975
<EOL>|976,977
ALT|977,980
16|981,983
,|983,984
Lip|985,988
70|989,991
,|991,992
trop|993,997
-|997,998
T|998,999
<|1000,1001
0.01|1002,1006
,|1006,1007
Chem|1008,1012
hemolyzed|1013,1022
but|1023,1026
Cr|1027,1029
1.4|1030,1033
<EOL>|1034,1035
(|1035,1036
baseline|1036,1044
1.0|1045,1048
in|1049,1051
_|1052,1053
_|1053,1054
_|1054,1055
,|1055,1056
repeat|1057,1063
K|1064,1065
3.6|1066,1069
.|1069,1070
Hyperglycemic|1071,1084
to|1085,1087
446|1088,1091
,|1091,1092
340|1093,1096
<EOL>|1097,1098
on|1098,1100
repeat|1101,1107
.|1107,1108
CXR|1109,1112
showed|1113,1119
no|1120,1122
acute|1123,1128
process|1129,1136
.|1136,1137
Patient|1138,1145
was|1146,1149
given|1150,1155
1L|1156,1158
NS|1159,1161
,|1161,1162
<EOL>|1163,1164
1g|1164,1166
CTX|1167,1170
,|1170,1171
14|1172,1174
units|1175,1180
insulin|1181,1188
.|1188,1189
Unclear|1190,1197
if|1198,1200
she|1201,1204
received|1205,1213
her|1214,1217
home|1218,1222
<EOL>|1223,1224
long|1224,1228
-|1228,1229
acting|1229,1235
insulin|1236,1243
.|1243,1244
UCx|1245,1248
and|1249,1252
BCx|1253,1256
's|1256,1258
were|1259,1263
sent|1264,1268
after|1269,1274
antibiotics|1275,1286
<EOL>|1287,1288
initiated.|1288,1298
Vitals|1299,1305
prior|1306,1311
to|1312,1314
transfer|1315,1323
were|1324,1328
:|1328,1329
3|1330,1331
98.4|1332,1336
89|1337,1339
152|1340,1343
/|1343,1344
80|1344,1346
20|1347,1349
<EOL>|1350,1351
100|1351,1354
%|1354,1355
RA|1356,1358
.|1358,1359
<EOL>|1361,1362
<EOL>|1362,1363
<EOL>|1364,1365
Past|1365,1369
Medical|1370,1377
History|1378,1385
:|1385,1386
<EOL>|1386,1387
COPD|1387,1391
<EOL>|1393,1394
CAD|1394,1397
s|1398,1399
/|1399,1400
p|1400,1401
CABG|1402,1406
and|1407,1410
stenting|1411,1419
<EOL>|1421,1422
Depression|1422,1432
<EOL>|1434,1435
DM|1435,1437
<EOL>|1439,1440
GERD|1440,1444
<EOL>|1446,1447
HTN|1447,1450
<EOL>|1452,1453
Migraines|1453,1462
<EOL>|1464,1465
Chronic|1465,1472
shoulder|1473,1481
pain|1482,1486
on|1487,1489
narcotics|1490,1499
<EOL>|1501,1502
OSA|1502,1505
<EOL>|1507,1508
Peripheral|1508,1518
neuropathy|1519,1529
<EOL>|1531,1532
Restless|1532,1540
leg|1541,1544
<EOL>|1546,1547
<EOL>|1547,1548
<EOL>|1549,1550
Social|1550,1556
History|1557,1564
:|1564,1565
<EOL>|1565,1566
_|1566,1567
_|1567,1568
_|1568,1569
<EOL>|1569,1570
Family|1570,1576
History|1577,1584
:|1584,1585
<EOL>|1585,1586
Mother|1586,1592
Unknown|1593,1600
ALCOHOL|1601,1608
ABUSE|1609,1614
pt|1615,1617
was|1618,1621
ward|1622,1626
of|1627,1629
state|1630,1635
,|1635,1636
does|1637,1641
n't|1641,1644
know|1645,1649
<EOL>|1650,1651
full|1651,1655
details|1656,1663
of|1664,1666
family|1667,1673
hx|1674,1676
<EOL>|1678,1679
Father|1679,1685
_|1686,1687
_|1687,1688
_|1688,1689
_|1690,1691
_|1691,1692
_|1692,1693
HODGKIN|1694,1701
'S|1701,1703
DISEASE|1704,1711
per|1712,1715
old|1716,1719
records|1720,1727
<EOL>|1729,1730
<EOL>|1730,1731
<EOL>|1732,1733
Physical|1733,1741
Exam|1742,1746
:|1746,1747
<EOL>|1747,1748
Admission|1748,1757
Physical|1758,1766
Exam|1767,1771
:|1771,1772
<EOL>|1772,1773
Vitals|1773,1779
-|1780,1781
98.3|1782,1786
155|1787,1790
/|1790,1791
88|1791,1793
92|1794,1796
20|1797,1799
99|1800,1802
%|1802,1803
on|1804,1806
RA|1807,1809
<EOL>|1811,1812
GENERAL|1812,1819
:|1819,1820
NAD|1821,1824
<EOL>|1826,1827
HEENT|1827,1832
:|1832,1833
NCAT|1834,1838
<EOL>|1840,1841
CARDIAC|1841,1848
:|1848,1849
RRR|1850,1853
,|1853,1854
S1|1855,1857
/|1857,1858
S2|1858,1860
,|1860,1861
no|1862,1864
murmurs|1865,1872
,|1872,1873
gallops|1874,1881
,|1881,1882
or|1883,1885
rubs|1886,1890
<EOL>|1892,1893
LUNG|1893,1897
:|1897,1898
CTAB|1899,1903
,|1903,1904
no|1905,1907
wheezes|1908,1915
,|1915,1916
rales|1917,1922
,|1922,1923
rhonchi|1924,1931
,|1931,1932
breathing|1933,1942
comfortably|1943,1954
<EOL>|1955,1956
without|1956,1963
use|1964,1967
of|1968,1970
accessory|1971,1980
muscles|1981,1988
<EOL>|1990,1991
ABDOMEN|1991,1998
:|1998,1999
nondistended|2000,2012
,|2012,2013
+|2014,2015
BS|2015,2017
,|2017,2018
nontender|2019,2028
in|2029,2031
all|2032,2035
quadrants|2036,2045
,|2045,2046
no|2047,2049
<EOL>|2050,2051
rebound|2051,2058
/|2058,2059
guarding|2059,2067
<EOL>|2069,2070
EXTREMITIES|2070,2081
:|2081,2082
no|2083,2085
cyanosis|2086,2094
,|2094,2095
clubbing|2096,2104
or|2105,2107
edema|2108,2113
,|2113,2114
moving|2115,2121
all|2122,2125
4|2126,2127
<EOL>|2128,2129
extremities|2129,2140
with|2141,2145
purpose|2146,2153
<EOL>|2155,2156
BACK|2156,2160
:|2160,2161
no|2162,2164
tenderness|2165,2175
to|2176,2178
spinal|2179,2185
processes|2186,2195
,|2195,2196
no|2197,2199
pain|2200,2204
the|2205,2208
left|2209,2213
side|2214,2218
,|2218,2219
<EOL>|2220,2221
+|2221,2222
CVA|2222,2225
tenderness|2226,2236
,|2236,2237
tenderness|2238,2248
to|2249,2251
palpation|2252,2261
of|2262,2264
the|2265,2268
R|2269,2270
sided|2271,2276
<EOL>|2277,2278
paraspinal|2278,2288
muscles|2289,2296
along|2297,2302
entire|2303,2309
length|2310,2316
of|2317,2319
spinal|2320,2326
cord|2327,2331
<EOL>|2333,2334
<EOL>|2334,2335
Discharge|2335,2344
Physical|2345,2353
Exam|2354,2358
:|2358,2359
<EOL>|2359,2360
Vitals|2360,2366
:|2366,2367
97.8|2368,2372
107|2373,2376
/|2376,2377
59|2377,2379
78|2380,2382
18|2383,2385
97|2386,2388
/|2388,2389
RA|2389,2391
<EOL>|2391,2392
General|2392,2399
:|2399,2400
awake|2401,2406
,|2406,2407
alert|2408,2413
,|2413,2414
NAD|2415,2418
<EOL>|2418,2419
HEENT|2419,2424
:|2424,2425
NCAT|2426,2430
EOMI|2431,2435
MMM|2436,2439
grossly|2440,2447
normal|2448,2454
oropharynx|2455,2465
<EOL>|2465,2466
CV|2466,2468
:|2468,2469
RRR|2470,2473
nl|2474,2476
S1|2477,2479
+|2479,2480
S2|2480,2482
no|2483,2485
g|2486,2487
/|2487,2488
r|2488,2489
/|2489,2490
m|2490,2491
no|2492,2494
JVD|2495,2498
/|2498,2499
HJR|2499,2502
.|2502,2503
<EOL>|2504,2505
Lungs|2505,2510
:|2510,2511
CTAB|2512,2516
no|2517,2519
w|2520,2521
/|2521,2522
r|2522,2523
/|2523,2524
r|2524,2525
,|2525,2526
good|2527,2531
movement|2532,2540
in|2541,2543
all|2544,2547
fields|2548,2554
<EOL>|2554,2555
Abdomen|2555,2562
:|2562,2563
obese|2564,2569
,|2569,2570
soft|2571,2575
nt|2576,2578
/|2578,2579
nd|2579,2581
normoactive|2582,2593
BS|2594,2596
<EOL>|2596,2597
Back|2597,2601
:|2601,2602
ttp|2603,2606
along|2607,2612
right|2613,2618
paraspinal|2619,2629
region|2630,2636
from|2637,2641
sacrum|2642,2648
to|2649,2651
shoulder|2652,2660
.|2660,2661
<EOL>|2662,2663
+|2663,2664
CVA|2665,2668
tenderness|2669,2679
.|2679,2680
<EOL>|2680,2681
Ext|2681,2684
:|2684,2685
dry|2686,2689
and|2690,2693
WWP|2694,2697
.|2697,2698
no|2699,2701
c|2702,2703
/|2703,2704
c|2704,2705
/|2705,2706
e|2706,2707
<EOL>|2707,2708
Neuro|2708,2713
:|2713,2714
AAOx3|2715,2720
,|2720,2721
moving|2722,2728
all|2729,2732
extrem|2733,2739
with|2740,2744
purpose|2745,2752
,|2752,2753
facial|2754,2760
movements|2761,2770
<EOL>|2771,2772
symmetric|2772,2781
,|2781,2782
no|2783,2785
focal|2786,2791
deficits|2792,2800
.|2800,2801
<EOL>|2801,2802
Skin|2802,2806
:|2806,2807
no|2808,2810
rashes|2811,2817
,|2817,2818
lesions|2819,2826
,|2826,2827
excoriations|2828,2840
<EOL>|2840,2841
<EOL>|2841,2842
<EOL>|2843,2844
Pertinent|2844,2853
Results|2854,2861
:|2861,2862
<EOL>|2862,2863
CT|2863,2865
ABD|2866,2869
/|2869,2870
PELVIS|2870,2876
_|2877,2878
_|2878,2879
_|2879,2880
:|2880,2881
<EOL>|2881,2882
Noncontrast|2882,2893
imaging|2894,2901
of|2902,2904
the|2905,2908
abdomen|2909,2916
and|2917,2920
pelvis|2921,2927
demonstrates|2928,2940
a|2941,2942
<EOL>|2943,2944
punctate|2944,2952
<EOL>|2953,2954
nonobstructing|2954,2968
calculus|2969,2977
in|2978,2980
the|2981,2984
right|2985,2990
collecting|2991,3001
system|3002,3008
(|3009,3010
02|3010,3012
:|3012,3013
31|3013,3015
)|3015,3016
.|3016,3017
<EOL>|3018,3019
There|3019,3024
is|3025,3027
no|3028,3030
left|3031,3035
renal|3036,3041
calculus|3042,3050
.|3050,3051
There|3052,3057
is|3058,3060
no|3061,3063
evidence|3064,3072
of|3073,3075
<EOL>|3076,3077
ureteral|3077,3085
or|3086,3088
urinary|3089,3096
bladder|3097,3104
calculus|3105,3113
.|3113,3114
There|3115,3120
is|3121,3123
symmetric|3124,3133
renal|3134,3139
<EOL>|3140,3141
enhancement|3141,3152
and|3153,3156
excretion|3157,3166
of|3167,3169
intravenous|3170,3181
contrast|3182,3190
.|3190,3191
Subcentimeter|3192,3205
<EOL>|3206,3207
cortically|3207,3217
based|3218,3223
hypodensity|3224,3235
in|3236,3238
the|3239,3242
left|3243,3247
interpolar|3248,3258
region|3259,3265
<EOL>|3266,3267
(|3267,3268
06|3268,3270
:|3270,3271
30|3271,3273
)|3273,3274
is|3275,3277
too|3278,3281
small|3282,3287
to|3288,3290
accurately|3291,3301
characterize|3302,3314
but|3315,3318
likely|3319,3325
<EOL>|3326,3327
represents|3327,3337
renal|3338,3343
cyst|3344,3348
.|3348,3349
There|3350,3355
is|3356,3358
no|3359,3361
evidence|3362,3370
of|3371,3373
collecting|3374,3384
system|3385,3391
<EOL>|3392,3393
filling|3393,3400
defect|3401,3407
.|3407,3408
There|3409,3414
are|3415,3418
segments|3419,3427
of|3428,3430
the|3431,3434
mid|3435,3438
to|3439,3441
distal|3442,3448
ureters|3449,3456
<EOL>|3457,3458
are|3458,3461
not|3462,3465
well|3466,3470
opacified|3471,3480
,|3480,3481
possibly|3482,3490
secondary|3491,3500
to|3501,3503
peristalsis|3504,3515
,|3515,3516
<EOL>|3517,3518
however|3518,3525
there|3526,3531
is|3532,3534
no|3535,3537
evidence|3538,3546
of|3547,3549
inflammatory|3550,3562
change|3563,3569
or|3570,3572
mass|3573,3577
<EOL>|3578,3579
about|3579,3584
the|3585,3588
ureters|3589,3596
.|3596,3597
The|3598,3601
adrenal|3602,3609
glands|3610,3616
are|3617,3620
unremarkable|3621,3633
.|3633,3634
<EOL>|3635,3636
<EOL>|3638,3639
Low|3639,3642
hepatic|3643,3650
attenuation|3651,3662
on|3663,3665
noncontrast|3666,3677
imaging|3678,3685
is|3686,3688
consistent|3689,3699
<EOL>|3700,3701
with|3701,3705
hepatic|3706,3713
<EOL>|3714,3715
steatosis|3715,3724
.|3724,3725
There|3726,3731
is|3732,3734
no|3735,3737
evidence|3738,3746
of|3747,3749
focal|3750,3755
hepatic|3756,3763
mass|3764,3768
.|3768,3769
There|3770,3775
is|3776,3778
<EOL>|3779,3780
no|3780,3782
<EOL>|3783,3784
intrahepatic|3784,3796
or|3797,3799
extrahepatic|3800,3812
biliary|3813,3820
ductal|3821,3827
dilatation|3828,3838
.|3838,3839
There|3840,3845
<EOL>|3846,3847
are|3847,3850
numerous|3851,3859
gallstones|3860,3870
within|3871,3877
the|3878,3881
gallbladder|3882,3893
without|3894,3901
evidence|3902,3910
<EOL>|3911,3912
of|3912,3914
acute|3915,3920
cholecystitis|3921,3934
.|3934,3935
<EOL>|3936,3937
<EOL>|3939,3940
The|3940,3943
spleen|3944,3950
is|3951,3953
not|3954,3957
enlarged|3958,3966
.|3966,3967
There|3968,3973
is|3974,3976
no|3977,3979
pancreatic|3980,3990
ductal|3991,3997
<EOL>|3998,3999
dilatation|3999,4009
or|4010,4012
<EOL>|4013,4014
evidence|4014,4022
of|4023,4025
pancreatic|4026,4036
mass|4037,4041
.|4041,4042
<EOL>|4043,4044
<EOL>|4046,4047
There|4047,4052
are|4053,4056
no|4057,4059
dilated|4060,4067
loops|4068,4073
of|4074,4076
bowel|4077,4082
.|4082,4083
There|4084,4089
is|4090,4092
no|4093,4095
evidence|4096,4104
of|4105,4107
<EOL>|4108,4109
bowel|4109,4114
wall|4115,4119
<EOL>|4120,4121
thickening|4121,4131
.|4131,4132
There|4133,4138
is|4139,4141
no|4142,4144
intraperitoneal|4145,4160
free|4161,4165
air|4166,4169
or|4170,4172
free|4173,4177
fluid|4178,4183
.|4183,4184
<EOL>|4185,4186
<EOL>|4188,4189
There|4189,4194
are|4195,4198
no|4199,4201
enlarged|4202,4210
inguinal|4211,4219
,|4219,4220
iliac|4221,4226
chain|4227,4232
,|4232,4233
retrocrural|4234,4245
,|4245,4246
or|4247,4249
<EOL>|4250,4251
retroperitoneal|4251,4266
lymph|4267,4272
nodes|4273,4278
.|4278,4279
Abdominal|4280,4289
aorta|4290,4295
has|4296,4299
a|4300,4301
normal|4302,4308
course|4309,4315
<EOL>|4316,4317
and|4317,4320
caliber|4321,4328
with|4329,4333
moderate|4334,4342
atherosclerotic|4343,4358
calcification|4359,4372
.|4372,4373
There|4374,4379
<EOL>|4380,4381
is|4381,4383
atherosclerotic|4384,4399
calcification|4400,4413
of|4414,4416
the|4417,4420
superior|4421,4429
mesenteric|4430,4440
<EOL>|4441,4442
artery|4442,4448
origin|4449,4455
.|4455,4456
There|4457,4462
is|4463,4465
no|4466,4468
suspicious|4469,4479
osseous|4480,4487
lesion|4488,4494
.|4494,4495
<EOL>|4496,4497
<EOL>|4499,4500
IMPRESSION|4500,4510
:|4510,4511
<EOL>|4512,4513
1.|4513,4515
Tiny|4516,4520
nonobstructing|4521,4535
right|4536,4541
collecting|4542,4552
system|4553,4559
calculus|4560,4568
.|4568,4569
<EOL>|4570,4571
2.|4571,4573
Hepatic|4574,4581
steatosis|4582,4591
.|4591,4592
<EOL>|4593,4594
3.|4594,4596
3|4597,4598
nodular|4599,4606
pulmonary|4607,4616
densities|4617,4626
in|4627,4629
the|4630,4633
left|4634,4638
basilar|4639,4646
region|4647,4653
<EOL>|4654,4655
measuring|4655,4664
up|4665,4667
to|4668,4670
8|4671,4672
x|4673,4674
8|4675,4676
mm|4677,4679
.|4679,4680
These|4681,4686
findings|4687,4695
may|4696,4699
may|4700,4703
represent|4704,4713
areas|4714,4719
<EOL>|4720,4721
of|4721,4723
rounded|4724,4731
atelectasis|4732,4743
,|4743,4744
however|4745,4752
short|4753,4758
-|4758,4759
term|4759,4763
followup|4764,4772
with|4773,4777
<EOL>|4778,4779
nonemergent|4779,4790
CT|4791,4793
chest|4794,4799
is|4800,4802
recommended|4803,4814
.|4814,4815
<EOL>|4816,4817
<EOL>|4817,4818
ADMISSION|4818,4827
LABS|4828,4832
:|4832,4833
<EOL>|4833,4834
_|4834,4835
_|4835,4836
_|4836,4837
08|4838,4840
:|4840,4841
30PM|4841,4845
BLOOD|4846,4851
WBC|4852,4855
-|4855,4856
9.4|4856,4859
RBC|4860,4863
-|4863,4864
3|4864,4865
.|4865,4866
95|4866,4868
*|4868,4869
Hgb|4870,4873
-|4873,4874
13.3|4874,4878
Hct|4879,4882
-|4882,4883
37.4|4883,4887
<EOL>|4888,4889
MCV|4889,4892
-|4892,4893
95|4893,4895
MCH|4896,4899
-|4899,4900
33|4900,4902
.|4902,4903
7|4903,4904
*|4904,4905
MCHC|4906,4910
-|4910,4911
35|4911,4913
.|4913,4914
5|4914,4915
*|4915,4916
RDW|4917,4920
-|4920,4921
13.5|4921,4925
Plt|4926,4929
_|4930,4931
_|4931,4932
_|4932,4933
<EOL>|4933,4934
_|4934,4935
_|4935,4936
_|4936,4937
08|4938,4940
:|4940,4941
30PM|4941,4945
BLOOD|4946,4951
Neuts|4952,4957
-|4957,4958
70|4958,4960
.|4960,4961
1|4961,4962
*|4962,4963
_|4964,4965
_|4965,4966
_|4966,4967
Monos|4968,4973
-|4973,4974
5.2|4974,4977
Eos|4978,4981
-|4981,4982
1.6|4982,4985
<EOL>|4986,4987
Baso|4987,4991
-|4991,4992
0.7|4992,4995
<EOL>|4995,4996
_|4996,4997
_|4997,4998
_|4998,4999
08|5000,5002
:|5002,5003
30PM|5003,5007
BLOOD|5008,5013
Glucose|5014,5021
-|5021,5022
446|5022,5025
*|5025,5026
UreaN|5027,5032
-|5032,5033
18|5033,5035
Creat|5036,5041
-|5041,5042
1|5042,5043
.|5043,5044
4|5044,5045
*|5045,5046
Na|5047,5049
-|5049,5050
133|5050,5053
<EOL>|5054,5055
K|5055,5056
-|5056,5057
5|5057,5058
.|5058,5059
6|5059,5060
*|5060,5061
Cl|5062,5064
-|5064,5065
97|5065,5067
HCO3|5068,5072
-|5072,5073
21|5073,5075
*|5075,5076
AnGap|5077,5082
-|5082,5083
21|5083,5085
*|5085,5086
<EOL>|5086,5087
_|5087,5088
_|5088,5089
_|5089,5090
08|5091,5093
:|5093,5094
30PM|5094,5098
BLOOD|5099,5104
ALT|5105,5108
-|5108,5109
16|5109,5111
AST|5112,5115
-|5115,5116
54|5116,5118
*|5118,5119
AlkPhos|5120,5127
-|5127,5128
65|5128,5130
TotBili|5131,5138
-|5138,5139
0.4|5139,5142
<EOL>|5142,5143
_|5143,5144
_|5144,5145
_|5145,5146
08|5147,5149
:|5149,5150
30PM|5150,5154
BLOOD|5155,5160
Albumin|5161,5168
-|5168,5169
4.1|5169,5172
Calcium|5173,5180
-|5180,5181
9.1|5181,5184
Phos|5185,5189
-|5189,5190
3.9|5190,5193
Mg|5194,5196
-|5196,5197
1.8|5197,5200
<EOL>|5200,5201
_|5201,5202
_|5202,5203
_|5203,5204
08|5205,5207
:|5207,5208
30PM|5208,5212
BLOOD|5213,5218
cTropnT|5219,5226
-|5226,5227
<|5227,5228
0|5228,5229
.|5229,5230
01|5230,5232
<EOL>|5232,5233
_|5233,5234
_|5234,5235
_|5235,5236
08|5237,5239
:|5239,5240
30PM|5240,5244
BLOOD|5245,5250
Lipase|5251,5257
-|5257,5258
70|5258,5260
*|5260,5261
<EOL>|5261,5262
_|5262,5263
_|5263,5264
_|5264,5265
10|5266,5268
:|5268,5269
53PM|5269,5273
BLOOD|5274,5279
_|5280,5281
_|5281,5282
_|5282,5283
pO2|5284,5287
-|5287,5288
38|5288,5290
*|5290,5291
pCO2|5292,5296
-|5296,5297
45|5297,5299
pH|5300,5302
-|5302,5303
7.37|5303,5307
<EOL>|5308,5309
calTCO2|5309,5316
-|5316,5317
27|5317,5319
Base|5320,5324
XS|5325,5327
-|5327,5328
0|5328,5329
<EOL>|5329,5330
_|5330,5331
_|5331,5332
_|5332,5333
10|5334,5336
:|5336,5337
53PM|5337,5341
BLOOD|5342,5347
Lactate|5348,5355
-|5355,5356
3|5356,5357
.|5357,5358
0|5358,5359
*|5359,5360
K|5361,5362
-|5362,5363
3.6|5363,5366
<EOL>|5366,5367
_|5367,5368
_|5368,5369
_|5369,5370
10|5371,5373
:|5373,5374
53PM|5374,5378
BLOOD|5379,5384
O2|5385,5387
Sat|5388,5391
-|5391,5392
69|5392,5394
<EOL>|5394,5395
_|5395,5396
_|5396,5397
_|5397,5398
10|5399,5401
:|5401,5402
40PM|5402,5406
URINE|5407,5412
Blood|5413,5418
-|5418,5419
NEG|5419,5422
Nitrite|5423,5430
-|5430,5431
POS|5431,5434
Protein|5435,5442
-|5442,5443
NEG|5443,5446
<EOL>|5447,5448
Glucose|5448,5455
-|5455,5456
1000|5456,5460
Ketone|5461,5467
-|5467,5468
TR|5468,5470
Bilirub|5471,5478
-|5478,5479
NEG|5479,5482
Urobiln|5483,5490
-|5490,5491
NEG|5491,5494
pH|5495,5497
-|5497,5498
6.0|5498,5501
Leuks|5502,5507
-|5507,5508
MOD|5508,5511
<EOL>|5511,5512
_|5512,5513
_|5513,5514
_|5514,5515
10|5516,5518
:|5518,5519
40PM|5519,5523
URINE|5524,5529
RBC|5530,5533
-|5533,5534
3|5534,5535
*|5535,5536
WBC|5537,5540
-|5540,5541
19|5541,5543
*|5543,5544
Bacteri|5545,5552
-|5552,5553
FEW|5553,5556
Yeast|5557,5562
-|5562,5563
NONE|5563,5567
<EOL>|5568,5569
Epi|5569,5572
-|5572,5573
1|5573,5574
TransE|5575,5581
-|5581,5582
<|5582,5583
1|5583,5584
<EOL>|5584,5585
_|5585,5586
_|5586,5587
_|5587,5588
10|5589,5591
:|5591,5592
40PM|5592,5596
URINE|5597,5602
Color|5603,5608
-|5608,5609
Straw|5609,5614
Appear|5615,5621
-|5621,5622
Clear|5622,5627
Sp|5628,5630
_|5631,5632
_|5632,5633
_|5633,5634
<EOL>|5634,5635
<EOL>|5635,5636
DISHCARGE|5636,5645
LABS|5646,5650
:|5650,5651
<EOL>|5651,5652
_|5652,5653
_|5653,5654
_|5654,5655
07|5656,5658
:|5658,5659
00AM|5659,5663
BLOOD|5664,5669
WBC|5670,5673
-|5673,5674
7.0|5674,5677
RBC|5678,5681
-|5681,5682
3|5682,5683
.|5683,5684
37|5684,5686
*|5686,5687
Hgb|5688,5691
-|5691,5692
11|5692,5694
.|5694,5695
2|5695,5696
*|5696,5697
Hct|5698,5701
-|5701,5702
31|5702,5704
.|5704,5705
8|5705,5706
*|5706,5707
<EOL>|5708,5709
MCV|5709,5712
-|5712,5713
94|5713,5715
MCH|5716,5719
-|5719,5720
33|5720,5722
.|5722,5723
2|5723,5724
*|5724,5725
MCHC|5726,5730
-|5730,5731
35|5731,5733
.|5733,5734
2|5734,5735
*|5735,5736
RDW|5737,5740
-|5740,5741
12.9|5741,5745
Plt|5746,5749
_|5750,5751
_|5751,5752
_|5752,5753
<EOL>|5753,5754
_|5754,5755
_|5755,5756
_|5756,5757
06|5758,5760
:|5760,5761
23AM|5761,5765
BLOOD|5766,5771
Neuts|5772,5777
-|5777,5778
53.5|5778,5782
_|5783,5784
_|5784,5785
_|5785,5786
Monos|5787,5792
-|5792,5793
5.0|5793,5796
Eos|5797,5800
-|5800,5801
1.8|5801,5804
<EOL>|5805,5806
Baso|5806,5810
-|5810,5811
0.6|5811,5814
<EOL>|5814,5815
_|5815,5816
_|5816,5817
_|5817,5818
07|5819,5821
:|5821,5822
00AM|5822,5826
BLOOD|5827,5832
Glucose|5833,5840
-|5840,5841
254|5841,5844
*|5844,5845
UreaN|5846,5851
-|5851,5852
13|5852,5854
Creat|5855,5860
-|5860,5861
1.0|5861,5864
Na|5865,5867
-|5867,5868
136|5868,5871
<EOL>|5872,5873
K|5873,5874
-|5874,5875
3.9|5875,5878
Cl|5879,5881
-|5881,5882
101|5882,5885
HCO3|5886,5890
-|5890,5891
24|5891,5893
AnGap|5894,5899
-|5899,5900
15|5900,5902
<EOL>|5902,5903
_|5903,5904
_|5904,5905
_|5905,5906
07|5907,5909
:|5909,5910
00AM|5910,5914
BLOOD|5915,5920
ALT|5921,5924
-|5924,5925
14|5925,5927
AST|5928,5931
-|5931,5932
17|5932,5934
AlkPhos|5935,5942
-|5942,5943
50|5943,5945
<EOL>|5945,5946
_|5946,5947
_|5947,5948
_|5948,5949
07|5950,5952
:|5952,5953
00AM|5953,5957
BLOOD|5958,5963
Calcium|5964,5971
-|5971,5972
8.5|5972,5975
Phos|5976,5980
-|5980,5981
3.5|5981,5984
Mg|5985,5987
-|5987,5988
1|5988,5989
.|5989,5990
5|5990,5991
*|5991,5992
<EOL>|5992,5993
<EOL>|5993,5994
<EOL>|5995,5996
Brief|5996,6001
Hospital|6002,6010
Course|6011,6017
:|6017,6018
<EOL>|6018,6019
_|6019,6020
_|6020,6021
_|6021,6022
PMH|6023,6026
with|6027,6031
HTN|6032,6035
,|6035,6036
GERD|6037,6041
,|6041,6042
CAD|6043,6046
s|6047,6048
/|6048,6049
p|6049,6050
CABG|6051,6055
and|6056,6059
stenting|6060,6068
,|6068,6069
IDDM|6070,6074
with|6075,6079
R|6080,6081
<EOL>|6082,6083
flank|6083,6088
pain|6089,6093
presumed|6094,6102
to|6103,6105
musculoskeletal|6106,6121
in|6122,6124
nature|6125,6131
due|6132,6135
to|6136,6138
negative|6139,6147
<EOL>|6148,6149
workup|6149,6155
.|6155,6156
Incidental|6157,6167
UTI|6168,6171
/|6172,6173
asymptomatic|6174,6186
bacturia|6187,6195
.|6195,6196
<EOL>|6196,6197
<EOL>|6197,6198
ACUTE|6198,6203
ISSUES|6204,6210
:|6210,6211
<EOL>|6212,6213
#|6213,6214
UTI|6215,6218
/|6219,6220
Bacturia|6221,6229
:|6229,6230
Patient|6231,6238
presented|6239,6248
without|6249,6256
any|6257,6260
history|6261,6268
of|6269,6271
<EOL>|6272,6273
urinary|6273,6280
or|6281,6283
systemic|6284,6292
symptoms|6293,6301
,|6301,6302
but|6303,6306
was|6307,6310
started|6311,6318
on|6319,6321
ceftriaxone|6322,6333
in|6334,6336
<EOL>|6337,6338
the|6338,6341
ED|6342,6344
after|6345,6350
U|6351,6352
/|6352,6353
A|6353,6354
with|6355,6359
_|6360,6361
_|6361,6362
_|6362,6363
positive|6364,6372
and|6373,6376
19|6377,6379
WBCs|6380,6384
.|6384,6385
<EOL>|6386,6387
Antibiotics|6387,6398
were|6399,6403
taken|6404,6409
prior|6410,6415
to|6416,6418
drawing|6419,6426
urinary|6427,6434
or|6435,6437
blood|6438,6443
<EOL>|6444,6445
cultures|6445,6453
,|6453,6454
and|6455,6458
there|6459,6464
was|6465,6468
no|6469,6471
yield|6472,6477
.|6477,6478
Patient|6479,6486
switched|6487,6495
to|6496,6498
<EOL>|6499,6500
ciprofloxacin|6500,6513
and|6514,6517
received|6518,6526
a|6527,6528
three|6529,6534
day|6535,6538
total|6539,6544
antibiotic|6545,6555
course|6556,6562
.|6562,6563
<EOL>|6564,6565
CT|6565,6567
scan|6568,6572
performed|6573,6582
did|6583,6586
not|6587,6590
have|6591,6595
any|6596,6599
evidence|6600,6608
of|6609,6611
pyelonephritis|6612,6626
.|6626,6627
<EOL>|6628,6629
Antibiotics|6629,6640
were|6641,6645
discontinued|6646,6658
at|6659,6661
time|6662,6666
of|6667,6669
discharge|6670,6679
.|6679,6680
<EOL>|6680,6681
<EOL>|6681,6682
#|6682,6683
Flank|6684,6689
Pain|6690,6694
:|6694,6695
<EOL>|6696,6697
Patient|6697,6704
reported|6705,6713
3|6714,6715
weeks|6716,6721
of|6722,6724
back|6725,6729
/|6729,6730
flank|6730,6735
pain|6736,6740
,|6740,6741
constant|6742,6750
and|6751,6754
achy|6755,6759
<EOL>|6760,6761
in|6761,6763
nature|6764,6770
and|6771,6774
worsened|6775,6783
by|6784,6786
movement|6787,6795
.|6795,6796
Treated|6797,6804
with|6805,6809
<EOL>|6810,6811
anti-inflammatories|6811,6830
with|6831,6835
minimal|6836,6843
effect|6844,6850
.|6850,6851
CT|6852,6854
scan|6855,6859
demonstrated|6860,6872
no|6873,6875
<EOL>|6876,6877
nephrolithiasis|6877,6892
.|6892,6893
CXR|6894,6897
showed|6898,6904
no|6905,6907
bony|6908,6912
abnormality|6913,6924
,|6924,6925
but|6926,6929
could|6930,6935
not|6936,6939
<EOL>|6940,6941
totally|6941,6948
exclude|6949,6956
multiple|6957,6965
rib|6966,6969
fractures|6970,6979
.|6979,6980
Patient|6981,6988
's|6988,6990
pain|6991,6995
was|6996,6999
well|7000,7004
<EOL>|7005,7006
controlled|7006,7016
and|7017,7020
tolerating|7021,7031
PO|7032,7034
medications|7035,7046
,|7046,7047
so|7048,7050
she|7051,7054
was|7055,7058
discharged|7059,7069
<EOL>|7070,7071
with|7071,7075
PCP|7076,7079
following|7080,7089
for|7090,7093
further|7094,7101
workup|7102,7108
.|7108,7109
<EOL>|7109,7110
<EOL>|7110,7111
#|7111,7112
Diabetes|7113,7121
/|7122,7123
Hyperglycemia|7124,7137
:|7137,7138
<EOL>|7138,7139
Patient|7139,7146
had|7147,7150
persistently|7151,7163
<EOL>|7164,7165
<EOL>|7165,7166
#|7166,7167
IDDM|7168,7172
:|7172,7173
Last|7174,7178
A1C|7179,7182
(|7183,7184
_|7184,7185
_|7185,7186
_|7186,7187
)|7187,7188
8.0|7189,7192
.|7192,7193
Serum|7194,7199
glucose|7200,7207
initially|7208,7217
in|7218,7220
the|7221,7224
400s|7225,7229
<EOL>|7230,7231
and|7231,7234
Chem|7235,7239
-|7239,7240
7|7240,7241
with|7242,7246
gap|7247,7250
;|7250,7251
however|7252,7259
,|7259,7260
this|7261,7265
was|7266,7269
likely|7270,7276
_|7277,7278
_|7278,7279
_|7279,7280
lactate|7281,7288
and|7289,7292
<EOL>|7293,7294
unlikely|7294,7302
to|7303,7305
be|7306,7308
DKA|7309,7312
given|7313,7318
normal|7319,7325
pH|7326,7328
on|7329,7331
ABG|7332,7335
.|7335,7336
AM|7337,7339
glucose|7340,7347
218|7348,7351
.|7351,7352
<EOL>|7352,7353
-|7353,7354
continue|7355,7363
home|7364,7368
dose|7369,7373
lantus|7374,7380
90|7381,7383
units|7384,7389
qPM|7390,7393
<EOL>|7395,7396
-|7396,7397
per|7398,7401
_|7402,7403
_|7403,7404
_|7404,7405
records|7406,7413
,|7413,7414
is|7415,7417
on|7418,7420
a|7421,7422
very|7423,7427
aggressive|7428,7438
ISS|7439,7442
,|7442,7443
will|7444,7448
decrease|7449,7457
<EOL>|7458,7459
for|7459,7462
now|7463,7466
and|7467,7470
uptitrate|7471,7480
as|7481,7483
necessary|7484,7493
depending|7494,7503
on|7504,7506
_|7507,7508
_|7508,7509
_|7509,7510
<EOL>|7512,7513
<EOL>|7513,7514
#|7514,7515
_|7516,7517
_|7517,7518
_|7518,7519
on|7520,7522
CKD|7523,7526
:|7526,7527
Cr|7528,7530
elevated|7531,7539
at|7540,7542
1.4|7543,7546
from|7547,7551
baseline|7552,7560
1.0|7561,7564
.|7564,7565
Most|7566,7570
likely|7571,7577
<EOL>|7578,7579
pre-renal|7579,7588
in|7589,7591
the|7592,7595
setting|7596,7603
of|7604,7606
infection|7607,7616
.|7616,7617
Now|7618,7621
s|7622,7623
/|7623,7624
p|7624,7625
2L|7626,7628
IVF|7629,7632
in|7633,7635
the|7636,7639
ED|7640,7642
<EOL>|7643,7644
and|7644,7647
creatinine|7648,7658
has|7659,7662
corrected|7663,7672
to|7673,7675
1.0|7676,7679
.|7679,7680
Appears|7681,7688
euvolemic|7689,7698
,|7698,7699
maybe|7700,7705
<EOL>|7706,7707
slightly|7707,7715
up|7716,7718
.|7718,7719
<EOL>|7720,7721
-|7721,7722
consider|7723,7731
further|7732,7739
workup|7740,7746
if|7747,7749
no|7750,7752
improvement|7753,7764
(|7765,7766
urine|7766,7771
lytes|7772,7777
,|7777,7778
<EOL>|7779,7780
spinning|7780,7788
urine|7789,7794
,|7794,7795
renal|7796,7801
u|7802,7803
/|7803,7804
s|7804,7805
)|7805,7806
<EOL>|7808,7809
-|7809,7810
renally|7811,7818
dose|7819,7823
medications|7824,7835
for|7836,7839
now|7840,7843
<EOL>|7845,7846
<EOL>|7846,7847
CHRONIC|7847,7854
ISSUES|7855,7861
:|7861,7862
<EOL>|7862,7863
#|7863,7864
HF|7865,7867
with|7868,7872
pEF|7873,7876
/|7876,7877
CAD|7877,7880
s|7881,7882
/|7882,7883
p|7883,7884
CABG|7885,7889
and|7890,7893
stents|7894,7900
:|7900,7901
Was|7902,7905
not|7906,7909
an|7910,7912
active|7913,7919
issue|7920,7925
<EOL>|7926,7927
whil|7927,7931
inpatient|7932,7941
.|7941,7942
Fluid|7943,7948
use|7949,7952
was|7953,7956
judicious|7957,7966
.|7966,7967
Metoprolo|7968,7977
converted|7978,7987
to|7988,7990
<EOL>|7991,7992
short|7992,7997
acting|7998,8004
while|8005,8010
in|8011,8013
house|8014,8019
,|8019,8020
isosorbide|8021,8031
,|8031,8032
aspirin|8033,8040
and|8041,8044
<EOL>|8045,8046
atorvastatin|8046,8058
were|8059,8063
continued|8064,8073
.|8073,8074
Losartan|8075,8083
held|8084,8088
as|8089,8091
below|8092,8097
.|8097,8098
<EOL>|8100,8101
#|8101,8102
HTN|8103,8106
:|8106,8107
home|8108,8112
metoprolol|8113,8123
and|8124,8127
isosorbide|8128,8138
continued|8139,8148
,|8148,8149
losartan|8150,8158
held|8159,8163
<EOL>|8164,8165
while|8165,8170
inpt|8171,8175
as|8176,8178
pressures|8179,8188
were|8189,8193
soft|8194,8198
and|8199,8202
within|8203,8209
normal|8210,8216
range|8217,8222
.|8222,8223
<EOL>|8224,8225
Discharged|8225,8235
home|8236,8240
off|8241,8244
losartan|8245,8253
.|8253,8254
<EOL>|8254,8255
#|8255,8256
Restless|8257,8265
leg|8266,8269
syndrome|8270,8278
:|8278,8279
home|8280,8284
ropinarole|8285,8295
continued|8296,8305
<EOL>|8305,8306
#|8306,8307
Shoulder|8308,8316
pain|8317,8321
:|8321,8322
oxycodone|8323,8332
and|8333,8336
tylenol|8337,8344
seperately|8345,8355
dose|8356,8360
while|8361,8366
<EOL>|8367,8368
inpatient|8368,8377
<EOL>|8379,8380
#|8380,8381
COPD|8382,8386
:|8386,8387
home|8388,8392
advair|8393,8399
and|8400,8403
PRN|8404,8407
albuterol|8408,8417
nebs|8418,8422
were|8423,8427
continued|8428,8437
<EOL>|8439,8440
#|8440,8441
GERD|8442,8446
:|8446,8447
home|8448,8452
pantoprazole|8453,8465
continued|8466,8475
<EOL>|8476,8477
#|8477,8478
Insomnia|8479,8487
:|8487,8488
home|8489,8493
trazodone|8494,8503
continued|8504,8513
<EOL>|8515,8516
<EOL>|8516,8517
TRANSITIONAL|8517,8529
ISSUES|8530,8536
:|8536,8537
<EOL>|8537,8538
-|8538,8539
Losartan|8540,8548
held|8549,8553
inpatient|8554,8563
and|8564,8567
at|8568,8570
discharge|8571,8580
andpatient|8581,8591
blood|8592,8597
<EOL>|8598,8599
pressures|8599,8608
were|8609,8613
low|8614,8617
-|8617,8618
normal|8618,8624
.|8624,8625
PCP|8626,8629
to|8630,8632
determine|8633,8642
restart|8643,8650
.|8650,8651
<EOL>|8651,8652
-|8652,8653
Patient|8654,8661
to|8662,8664
follow|8665,8671
up|8672,8674
with|8675,8679
PCP|8680,8683
for|8684,8687
resolution|8688,8698
of|8699,8701
UTI|8702,8705
and|8706,8709
back|8710,8714
<EOL>|8715,8716
pain|8716,8720
symptoms|8721,8729
<EOL>|8729,8730
-|8730,8731
Patient|8732,8739
should|8740,8746
have|8747,8751
insulin|8752,8759
regiment|8760,8768
adjustments|8769,8780
for|8781,8784
optimal|8785,8792
<EOL>|8793,8794
glycemic|8794,8802
control|8803,8810
-|8811,8812
no|8813,8815
changes|8816,8823
to|8824,8826
regimen|8827,8834
were|8835,8839
made|8840,8844
at|8845,8847
discharge|8848,8857
.|8857,8858
<EOL>|8858,8859
<EOL>|8860,8861
Medications|8861,8872
on|8873,8875
Admission|8876,8885
:|8885,8886
<EOL>|8886,8887
The|8887,8890
Preadmission|8891,8903
Medication|8904,8914
list|8915,8919
may|8920,8923
be|8924,8926
inaccurate|8927,8937
and|8938,8941
requires|8942,8950
<EOL>|8951,8952
futher|8952,8958
investigation|8959,8972
.|8972,8973
<EOL>|8973,8974
1.|8974,8976
Losartan|8977,8985
Potassium|8986,8995
25|8996,8998
mg|8999,9001
PO|9002,9004
DAILY|9005,9010
<EOL>|9011,9012
2.|9012,9014
Metoprolol|9015,9025
Succinate|9026,9035
XL|9036,9038
200|9039,9042
mg|9043,9045
PO|9046,9048
DAILY|9049,9054
<EOL>|9055,9056
3.|9056,9058
Atorvastatin|9059,9071
80|9072,9074
mg|9075,9077
PO|9078,9080
HS|9081,9083
<EOL>|9084,9085
4.|9085,9087
Isosorbide|9088,9098
Mononitrate|9099,9110
(|9111,9112
Extended|9112,9120
Release|9121,9128
)|9128,9129
120|9130,9133
mg|9134,9136
PO|9137,9139
DAILY|9140,9145
<EOL>|9146,9147
5.|9147,9149
Nitroglycerin|9150,9163
SL|9164,9166
0.3|9167,9170
mg|9171,9173
SL|9174,9176
Q5MIN|9177,9182
:|9182,9183
PRN|9183,9186
pain|9187,9191
<EOL>|9192,9193
6.|9193,9195
Ropinirole|9196,9206
0.5|9207,9210
mg|9211,9213
PO|9214,9216
QPM|9217,9220
<EOL>|9221,9222
7.|9222,9224
Oxycodone|9225,9234
-|9234,9235
Acetaminophen|9235,9248
(|9249,9250
5mg|9250,9253
-|9253,9254
325mg|9254,9259
)|9259,9260
1|9261,9262
TAB|9263,9266
PO|9267,9269
Q8H|9270,9273
:|9273,9274
PRN|9274,9277
pain|9278,9282
<EOL>|9283,9284
8.|9284,9286
Fluticasone|9287,9298
Propionate|9299,9309
110mcg|9310,9316
2|9317,9318
PUFF|9319,9323
IH|9324,9326
BID|9327,9330
<EOL>|9331,9332
9.|9332,9334
Pantoprazole|9335,9347
40|9348,9350
mg|9351,9353
PO|9354,9356
Q12H|9357,9361
<EOL>|9362,9363
10.|9363,9366
Aspirin|9367,9374
325|9375,9378
mg|9379,9381
PO|9382,9384
DAILY|9385,9390
<EOL>|9391,9392
11.|9392,9395
albuterol|9396,9405
sulfate|9406,9413
90|9414,9416
mcg|9417,9420
/|9420,9421
actuation|9421,9430
inhalation|9431,9441
q4hrs|9442,9447
wheezing|9448,9456
<EOL>|9457,9458
<EOL>|9458,9459
12.|9459,9462
TraZODone|9463,9472
150|9473,9476
mg|9477,9479
PO|9480,9482
HS|9483,9485
<EOL>|9486,9487
13|9487,9489
.|9489,9490
Vitamin|9491,9498
D|9499,9500
1000|9501,9505
UNIT|9506,9510
PO|9511,9513
DAILY|9514,9519
<EOL>|9520,9521
14.|9521,9524
Levemir|9525,9532
Flexpen|9533,9540
(|9541,9542
insulin|9542,9549
detemir|9550,9557
)|9557,9558
90|9559,9561
units|9562,9567
subcutaneous|9568,9580
in|9581,9583
<EOL>|9584,9585
the|9585,9588
evening|9589,9596
<EOL>|9597,9598
15.|9598,9601
HumaLOG|9602,9609
KwikPen|9610,9617
(|9618,9619
insulin|9619,9626
lispro|9627,9633
)|9633,9634
per|9635,9638
sliding|9639,9646
scale|9647,9652
<EOL>|9654,9655
subcutaneous|9655,9667
as|9668,9670
directed|9671,9679
<EOL>|9680,9681
<EOL>|9681,9682
<EOL>|9683,9684
Discharge|9684,9693
Medications|9694,9705
:|9705,9706
<EOL>|9706,9707
1.|9707,9709
Oxycodone|9710,9719
-|9719,9720
Acetaminophen|9720,9733
(|9734,9735
5mg|9735,9738
-|9738,9739
325mg|9739,9744
)|9744,9745
1|9746,9747
TAB|9748,9751
PO|9752,9754
Q8H|9755,9758
:|9758,9759
PRN|9759,9762
pain|9763,9767
<EOL>|9768,9769
2.|9769,9771
Nitroglycerin|9772,9785
SL|9786,9788
0.3|9789,9792
mg|9793,9795
SL|9796,9798
Q5MIN|9799,9804
:|9804,9805
PRN|9805,9808
pain|9809,9813
<EOL>|9814,9815
3.|9815,9817
Metoprolol|9818,9828
Succinate|9829,9838
XL|9839,9841
200|9842,9845
mg|9846,9848
PO|9849,9851
DAILY|9852,9857
<EOL>|9858,9859
4.|9859,9861
Levemir|9862,9869
Flexpen|9870,9877
(|9878,9879
insulin|9879,9886
detemir|9887,9894
)|9894,9895
90|9896,9898
units|9899,9904
subcutaneous|9905,9917
in|9918,9920
<EOL>|9921,9922
the|9922,9925
evening|9926,9933
<EOL>|9934,9935
5.|9935,9937
HumaLOG|9938,9945
KwikPen|9946,9953
(|9954,9955
insulin|9955,9962
lispro|9963,9969
)|9969,9970
0|9971,9972
SUBCUTANEOUS|9975,9987
AS|9988,9990
DIRECTED|9991,9999
<EOL>|10000,10001
<EOL>|10001,10002
6.|10002,10004
albuterol|10005,10014
sulfate|10015,10022
90|10023,10025
mcg|10026,10029
/|10029,10030
actuation|10030,10039
inhalation|10040,10050
q4hrs|10051,10056
wheezing|10057,10065
<EOL>|10066,10067
7.|10067,10069
Ciprofloxacin|10070,10083
HCl|10084,10087
500|10088,10091
mg|10092,10094
PO|10095,10097
Q12H|10098,10102
Duration|10103,10111
:|10111,10112
7|10113,10114
Days|10115,10119
<EOL>|10120,10121
RX|10121,10123
*|10124,10125
ciprofloxacin|10125,10138
[|10139,10140
Cipro|10140,10145
]|10145,10146
500|10147,10150
mg|10151,10153
1|10154,10155
tablet|10156,10162
(|10162,10163
s|10163,10164
)|10164,10165
by|10166,10168
mouth|10169,10174
twice|10175,10180
a|10181,10182
<EOL>|10183,10184
day|10184,10187
Disp|10188,10192
#|10193,10194
*|10194,10195
11|10195,10197
Tablet|10198,10204
Refills|10205,10212
:|10212,10213
*|10213,10214
0|10214,10215
<EOL>|10215,10216
8.|10216,10218
Vitamin|10219,10226
D|10227,10228
1000|10229,10233
UNIT|10234,10238
PO|10239,10241
DAILY|10242,10247
<EOL>|10248,10249
9.|10249,10251
TraZODone|10252,10261
150|10262,10265
mg|10266,10268
PO|10269,10271
HS|10272,10274
<EOL>|10275,10276
10.|10276,10279
Isosorbide|10280,10290
Mononitrate|10291,10302
(|10303,10304
Extended|10304,10312
Release|10313,10320
)|10320,10321
120|10322,10325
mg|10326,10328
PO|10329,10331
DAILY|10332,10337
<EOL>|10338,10339
11.|10339,10342
Aspirin|10343,10350
325|10351,10354
mg|10355,10357
PO|10358,10360
DAILY|10361,10366
<EOL>|10367,10368
12.|10368,10371
Atorvastatin|10372,10384
80|10385,10387
mg|10388,10390
PO|10391,10393
HS|10394,10396
<EOL>|10397,10398
13.|10398,10401
Fluticasone|10402,10413
Propionate|10414,10424
110mcg|10425,10431
2|10432,10433
PUFF|10434,10438
IH|10439,10441
BID|10442,10445
<EOL>|10446,10447
14.|10447,10450
Pantoprazole|10451,10463
40|10464,10466
mg|10467,10469
PO|10470,10472
Q12H|10473,10477
<EOL>|10478,10479
15.|10479,10482
Ropinirole|10483,10493
0.5|10494,10497
mg|10498,10500
PO|10501,10503
QPM|10504,10507
<EOL>|10508,10509
<EOL>|10509,10510
<EOL>|10511,10512
Discharge|10512,10521
Disposition|10522,10533
:|10533,10534
<EOL>|10534,10535
Home|10535,10539
<EOL>|10539,10540
<EOL>|10541,10542
Discharge|10542,10551
Diagnosis|10552,10561
:|10561,10562
<EOL>|10562,10563
Primary|10563,10570
Diagnosis|10571,10580
:|10580,10581
<EOL>|10581,10582
UTI|10582,10585
<EOL>|10585,10586
<EOL>|10586,10587
Secondary|10587,10596
Diagnosis|10597,10606
:|10606,10607
<EOL>|10607,10608
Back|10608,10612
Pain|10613,10617
<EOL>|10617,10618
Diabetes|10618,10626
<EOL>|10626,10627
<EOL>|10627,10628
<EOL>|10629,10630
Discharge|10630,10639
Condition|10640,10649
:|10649,10650
<EOL>|10650,10651
Mental|10651,10657
Status|10658,10664
:|10664,10665
Clear|10666,10671
and|10672,10675
coherent|10676,10684
.|10684,10685
<EOL>|10685,10686
Level|10686,10691
of|10692,10694
Consciousness|10695,10708
:|10708,10709
Alert|10710,10715
and|10716,10719
interactive|10720,10731
.|10731,10732
<EOL>|10732,10733
Activity|10733,10741
Status|10742,10748
:|10748,10749
Ambulatory|10750,10760
-|10761,10762
Independent|10763,10774
.|10774,10775
<EOL>|10775,10776
<EOL>|10776,10777
<EOL>|10778,10779
Discharge|10779,10788
Instructions|10789,10801
:|10801,10802
<EOL>|10802,10803
Dear|10803,10807
_|10808,10809
_|10809,10810
_|10810,10811
,|10811,10812
<EOL>|10812,10813
<EOL>|10813,10814
_|10814,10815
_|10815,10816
_|10816,10817
were|10818,10822
seen|10823,10827
in|10828,10830
the|10831,10834
emergency|10835,10844
department|10845,10855
for|10856,10859
back|10860,10864
pain|10865,10869
.|10869,10870
_|10871,10872
_|10872,10873
_|10873,10874
<EOL>|10875,10876
were|10876,10880
admitted|10881,10889
to|10890,10892
the|10893,10896
hospital|10897,10905
where|10906,10911
_|10912,10913
_|10913,10914
_|10914,10915
were|10916,10920
also|10921,10925
diagnosed|10926,10935
with|10936,10940
<EOL>|10941,10942
a|10942,10943
urinary|10944,10951
tract|10952,10957
infection|10958,10967
.|10967,10968
_|10969,10970
_|10970,10971
_|10971,10972
were|10973,10977
treated|10978,10985
with|10986,10990
antibiotics|10991,11002
,|11002,11003
IV|11004,11006
<EOL>|11007,11008
fluids|11008,11014
and|11015,11018
pain|11019,11023
medication|11024,11034
.|11034,11035
Due|11036,11039
to|11040,11042
the|11043,11046
concern|11047,11054
of|11055,11057
your|11058,11062
back|11063,11067
<EOL>|11068,11069
pain|11069,11073
,|11073,11074
a|11075,11076
CT|11077,11079
scan|11080,11084
was|11085,11088
as|11089,11091
performed|11092,11101
and|11102,11105
it|11106,11108
was|11109,11112
determined|11113,11123
that|11124,11128
_|11129,11130
_|11130,11131
_|11131,11132
<EOL>|11133,11134
did|11134,11137
not|11138,11141
have|11142,11146
a|11147,11148
kidney|11149,11155
stone|11156,11161
or|11162,11164
an|11165,11167
infection|11168,11177
.|11177,11178
Your|11179,11183
diabetes|11184,11192
was|11193,11196
<EOL>|11197,11198
controlled|11198,11208
with|11209,11213
an|11214,11216
insulin|11217,11224
scale|11225,11230
while|11231,11236
_|11237,11238
_|11238,11239
_|11239,11240
were|11241,11245
an|11246,11248
inpatient|11249,11258
.|11258,11259
<EOL>|11260,11261
_|11261,11262
_|11262,11263
_|11263,11264
will|11265,11269
be|11270,11272
discharged|11273,11283
home|11284,11288
on|11289,11291
antibiotics|11292,11303
and|11304,11307
intent|11308,11314
to|11315,11317
follow|11318,11324
<EOL>|11325,11326
up|11326,11328
with|11329,11333
your|11334,11338
primary|11339,11346
care|11347,11351
provider|11352,11360
,|11360,11361
Dr.|11362,11365
_|11366,11367
_|11367,11368
_|11368,11369
.|11369,11370
Please|11371,11377
take|11378,11382
all|11383,11386
<EOL>|11387,11388
medications|11388,11399
as|11400,11402
prescribed|11403,11413
and|11414,11417
keep|11418,11422
all|11423,11426
scheduled|11427,11436
appointments|11437,11449
.|11449,11450
<EOL>|11451,11452
Weigh|11452,11457
yourself|11458,11466
every|11467,11472
morning|11473,11480
,|11480,11481
call|11482,11486
MD|11487,11489
if|11490,11492
weight|11493,11499
goes|11500,11504
up|11505,11507
more|11508,11512
<EOL>|11513,11514
than|11514,11518
3|11519,11520
lbs|11521,11524
.|11524,11525
<EOL>|11525,11526
<EOL>|11526,11527
It|11527,11529
was|11530,11533
a|11534,11535
pleasure|11536,11544
taking|11545,11551
care|11552,11556
of|11557,11559
_|11560,11561
_|11561,11562
_|11562,11563
!|11563,11564
<EOL>|11564,11565
Your|11565,11569
_|11570,11571
_|11571,11572
_|11572,11573
Care|11574,11578
Team|11579,11583
<EOL>|11583,11584
<EOL>|11585,11586
Followup|11586,11594
Instructions|11595,11607
:|11607,11608
<EOL>|11608,11609
_|11609,11610
_|11610,11611
_|11611,11612
<EOL>|11612,11613

