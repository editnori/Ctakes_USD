 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
Chief|240,245
Complaint|246,255
:|255,256
<EOL>|256,257
Syncope|257,264
<EOL>|264,265
<EOL>|266,267
Major|267,272
Surgical|273,281
or|282,284
Invasive|285,293
Procedure|294,303
:|303,304
<EOL>|304,305
None|305,309
<EOL>|309,310
<EOL>|311,312
History|312,319
of|320,322
Present|323,330
Illness|331,338
:|338,339
<EOL>|339,340
Ms.|340,343
_|344,345
_|345,346
_|346,347
is|348,350
a|351,352
_|353,354
_|354,355
_|355,356
w|357,358
/|358,359
hx|359,361
of|362,364
AR|365,367
,|367,368
hypothyroidism|369,383
,|383,384
Sjogrens|385,393
,|393,394
HTN|395,398
,|398,399
<EOL>|400,401
PNA|401,404
who|405,408
presents|409,417
as|418,420
a|421,422
transfer|423,431
from|432,436
_|437,438
_|438,439
_|439,440
after|441,446
a|447,448
syncopal|449,457
<EOL>|458,459
episode|459,466
on|467,469
_|470,471
_|471,472
_|472,473
AM|474,476
.|476,477
She|478,481
was|482,485
standing|486,494
and|495,498
speaking|499,507
with|508,512
her|513,516
<EOL>|517,518
daughter|518,526
when|527,531
she|532,535
began|536,541
to|542,544
feel|545,549
weak|550,554
,|554,555
lightheaded|556,567
,|567,568
and|569,572
nauseous|573,581
.|581,582
<EOL>|583,584
She|584,587
has|588,591
had|592,595
a|596,597
few|598,601
syncopal|602,610
episodes|611,619
in|620,622
the|623,626
past|627,631
,|631,632
which|633,638
she|639,642
<EOL>|643,644
reports|644,651
were|652,656
concurrent|657,667
with|668,672
other|673,678
health|679,685
problems|686,694
such|695,699
as|700,702
a|703,704
<EOL>|705,706
recent|706,712
PNA|713,716
in|717,719
_|720,721
_|721,722
_|722,723
with|724,728
hemoptysis|729,739
treated|740,747
at|748,750
_|751,752
_|752,753
_|753,754
(|755,756
CT|756,758
scan|759,763
<EOL>|764,765
showed|765,771
RML|772,775
brochiectasis|776,789
and|790,793
some|794,798
consolidation|799,812
;|812,813
bronch|814,820
showed|821,827
<EOL>|828,829
copious|829,836
mucoid|837,843
secretions|844,854
RML|855,858
>|858,859
lingula|859,866
>|866,867
RUL|867,870
with|871,875
some|876,880
blood|881,886
,|886,887
pt|888,890
<EOL>|891,892
was|892,895
scheduled|896,905
for|906,909
rpt|910,913
CT|914,916
scan|917,921
on|922,924
_|925,926
_|926,927
_|927,928
.|928,929
<EOL>|929,930
.|930,931
<EOL>|931,932
On|932,934
_|935,936
_|936,937
_|937,938
,|938,939
she|940,943
sat|944,947
down|948,952
in|953,955
her|956,959
chair|960,965
and|966,969
then|970,974
passed|975,981
out|982,985
,|985,986
and|987,990
was|991,994
<EOL>|995,996
unresponsive|996,1008
for|1009,1012
a|1013,1014
few|1015,1018
seconds|1019,1026
.|1026,1027
The|1028,1031
pt|1032,1034
denies|1035,1041
prodrome|1042,1050
or|1051,1053
<EOL>|1054,1055
palpitations|1055,1067
,|1067,1068
and|1069,1072
regained|1073,1081
consciousness|1082,1095
quickly|1096,1103
with|1104,1108
no|1109,1111
<EOL>|1112,1113
confusion|1113,1122
afterwards|1123,1133
.|1133,1134
No|1135,1137
seizure|1138,1145
like|1146,1150
activity|1151,1159
witnessed|1160,1169
,|1169,1170
no|1171,1173
<EOL>|1174,1175
lose|1175,1179
of|1180,1182
bowel|1183,1188
or|1189,1191
bladder|1192,1199
.|1199,1200
Denies|1201,1207
any|1208,1211
recent|1212,1218
exertion|1219,1227
or|1228,1230
<EOL>|1231,1232
miturition|1232,1242
prior|1243,1248
to|1249,1251
episode|1252,1259
.|1259,1260
Denies|1261,1267
CP|1268,1270
,|1270,1271
palpitations|1272,1284
,|1284,1285
SOB|1286,1289
prior|1290,1295
<EOL>|1296,1297
or|1297,1299
after|1300,1305
the|1306,1309
episode|1310,1317
.|1317,1318
She|1319,1322
remembers|1323,1332
the|1333,1336
episode|1337,1344
.|1344,1345
She|1346,1349
states|1350,1356
she|1357,1360
<EOL>|1361,1362
has|1362,1365
been|1366,1370
coughing|1371,1379
for|1380,1383
the|1384,1387
past|1388,1392
few|1393,1396
days|1397,1401
,|1401,1402
occasionally|1403,1415
productive|1416,1426
<EOL>|1427,1428
with|1428,1432
phlegm|1433,1439
,|1439,1440
nonbloody|1441,1450
,|1450,1451
but|1452,1455
has|1456,1459
otherwise|1460,1469
been|1470,1474
well|1475,1479
,|1479,1480
with|1481,1485
no|1486,1488
<EOL>|1489,1490
fevers|1490,1496
/|1496,1497
chills|1497,1503
.|1503,1504
Her|1505,1508
last|1509,1513
echo|1514,1518
for|1519,1522
AR|1523,1525
_|1526,1527
_|1527,1528
_|1528,1529
years|1530,1535
ago|1536,1539
.|1539,1540
<EOL>|1540,1541
.|1541,1542
<EOL>|1542,1543
In|1543,1545
the|1546,1549
ED|1550,1552
,|1552,1553
initial|1554,1561
vitals|1562,1568
were|1569,1573
98.5|1574,1578
96|1579,1581
145|1582,1585
/|1585,1586
86|1586,1588
20|1589,1591
97|1592,1594
%|1594,1595
.|1595,1596
Labs|1597,1601
were|1602,1606
<EOL>|1607,1608
notable|1608,1615
for|1616,1619
WBC|1620,1623
12.0|1624,1628
(|1629,1630
with|1630,1634
N|1635,1636
76|1637,1639
.|1639,1640
5|1640,1641
%|1641,1642
,|1642,1643
L|1644,1645
17.3|1646,1650
%|1650,1651
)|1651,1652
,|1652,1653
Hct|1654,1657
32.6|1658,1662
.|1662,1663
UA|1665,1667
<EOL>|1668,1669
showed|1669,1675
lg|1676,1678
leuk|1679,1683
and|1684,1687
18|1688,1690
WBC|1691,1694
.|1694,1695
Vitals|1696,1702
prior|1703,1708
to|1709,1711
transfer|1712,1720
were|1721,1725
<EOL>|1726,1727
98|1727,1729
-|1729,1730
85|1730,1732
-|1732,1733
146|1733,1736
/|1736,1737
75|1737,1739
-|1739,1740
25|1740,1742
-|1742,1743
98|1743,1745
.|1745,1746
<EOL>|1746,1747
.|1747,1748
<EOL>|1748,1749
Currently|1749,1758
on|1759,1761
the|1762,1765
medicine|1766,1774
floor|1775,1780
,|1780,1781
she|1782,1785
feels|1786,1791
"|1792,1793
fine|1793,1797
"|1797,1798
and|1799,1802
does|1803,1807
not|1808,1811
<EOL>|1812,1813
feel|1813,1817
dizzy|1818,1823
or|1824,1826
lightheaded|1827,1838
.|1838,1839
She|1840,1843
denies|1844,1850
fever|1851,1856
,|1856,1857
chills|1858,1864
,|1864,1865
vision|1866,1872
<EOL>|1873,1874
changes|1874,1881
,|1881,1882
shortness|1883,1892
of|1893,1895
breath|1896,1902
,|1902,1903
chest|1904,1909
pain|1910,1914
,|1914,1915
abdominal|1916,1925
pain|1926,1930
,|1930,1931
<EOL>|1932,1933
nausea|1933,1939
,|1939,1940
vomiting|1941,1949
,|1949,1950
diarrhea|1951,1959
,|1959,1960
constipation|1961,1973
,|1973,1974
BRBPR|1975,1980
,|1980,1981
melena|1982,1988
,|1988,1989
<EOL>|1990,1991
hematochezia|1991,2003
,|2003,2004
dysuria|2005,2012
,|2012,2013
hematuria|2014,2023
.|2023,2024
She|2025,2028
does|2029,2033
say|2034,2037
she|2038,2041
lost|2042,2046
a|2047,2048
few|2049,2052
<EOL>|2053,2054
pounds|2054,2060
in|2061,2063
the|2064,2067
last|2068,2072
few|2073,2076
weeks|2077,2082
and|2083,2086
has|2087,2090
not|2091,2094
had|2095,2098
a|2099,2100
great|2101,2106
appetite|2107,2115
<EOL>|2116,2117
for|2117,2120
about|2121,2126
a|2127,2128
month|2129,2134
.|2134,2135
<EOL>|2135,2136
<EOL>|2137,2138
Past|2138,2142
Medical|2143,2150
History|2151,2158
:|2158,2159
<EOL>|2159,2160
HTN|2160,2163
<EOL>|2163,2164
Hypothyroidism|2164,2178
<EOL>|2178,2179
Sjo|2179,2182
_|2182,2183
_|2183,2184
_|2184,2185
'|2185,2186
s|2186,2187
Syd|2188,2191
<EOL>|2191,2192
<EOL>|2192,2193
<EOL>|2194,2195
Social|2195,2201
History|2202,2209
:|2209,2210
<EOL>|2210,2211
_|2211,2212
_|2212,2213
_|2213,2214
<EOL>|2214,2215
Family|2215,2221
History|2222,2229
:|2229,2230
<EOL>|2230,2231
Long|2231,2235
history|2236,2243
of|2244,2246
hypertension|2247,2259
in|2260,2262
her|2263,2266
family|2267,2273
.|2273,2274
She|2276,2279
does|2280,2284
report|2285,2291
<EOL>|2292,2293
that|2293,2297
her|2298,2301
father|2302,2308
's|2308,2310
family|2311,2317
has|2318,2321
a|2322,2323
history|2324,2331
of|2332,2334
multiple|2335,2343
cancers|2344,2351
.|2351,2352
She|2354,2357
<EOL>|2358,2359
has|2359,2362
a|2363,2364
grandfather|2365,2376
with|2377,2381
a|2382,2383
history|2384,2391
of|2392,2394
stomach|2395,2402
cancer|2403,2409
and|2410,2413
an|2414,2416
uncle|2417,2422
<EOL>|2423,2424
with|2424,2428
a|2429,2430
history|2431,2438
of|2439,2441
throat|2442,2448
cancer|2449,2455
.|2455,2456
She|2458,2461
denies|2462,2468
any|2469,2472
history|2473,2480
of|2481,2483
<EOL>|2484,2485
colon|2485,2490
cancers|2491,2498
.|2498,2499
Father|2500,2506
had|2507,2510
stroke|2511,2517
.|2517,2518
No|2519,2521
family|2522,2528
h|2529,2530
/|2530,2531
o|2531,2532
MI|2533,2535
.|2535,2536
Mother|2537,2543
had|2544,2547
a|2548,2549
<EOL>|2550,2551
heart|2551,2556
valve|2557,2562
replaced|2563,2571
(|2572,2573
pt|2573,2575
not|2576,2579
sure|2580,2584
which|2585,2590
one|2591,2594
)|2594,2595
.|2595,2596
<EOL>|2596,2597
<EOL>|2597,2598
<EOL>|2599,2600
Physical|2600,2608
Exam|2609,2613
:|2613,2614
<EOL>|2614,2615
ADMISSION|2615,2624
EXAM|2625,2629
:|2629,2630
<EOL>|2630,2631
<EOL>|2631,2632
VS|2632,2634
-|2635,2636
Temp|2637,2641
98.1|2642,2646
F|2646,2647
,|2647,2648
BP|2649,2651
112|2652,2655
/|2655,2656
70|2656,2658
,|2658,2659
HR|2660,2662
96|2663,2665
,|2665,2666
R|2667,2668
18|2669,2671
,|2671,2672
O2|2673,2675
-|2675,2676
sat|2676,2679
96|2680,2682
%|2682,2683
RA|2684,2686
<EOL>|2686,2687
GENERAL|2687,2694
-|2695,2696
thin|2697,2701
-|2701,2702
appearing|2702,2711
woman|2712,2717
in|2718,2720
NAD|2721,2724
,|2724,2725
comfortable|2726,2737
,|2737,2738
appropriate|2739,2750
<EOL>|2750,2751
HEENT|2751,2756
-|2757,2758
NC|2759,2761
/|2761,2762
AT|2762,2764
,|2764,2765
PERRL|2766,2771
,|2771,2772
EOMI|2773,2777
,|2777,2778
sclerae|2779,2786
anicteric|2787,2796
,|2796,2797
MMM|2798,2801
,|2801,2802
OP|2803,2805
clear|2806,2811
<EOL>|2811,2812
NECK|2812,2816
-|2817,2818
supple|2819,2825
,|2825,2826
no|2827,2829
thyromegaly|2830,2841
,|2841,2842
no|2843,2845
JVD|2846,2849
,|2849,2850
carotid|2851,2858
bruits|2859,2865
(|2866,2867
likely|2867,2873
<EOL>|2874,2875
radiating|2875,2884
sounds|2885,2891
from|2892,2896
aortic|2897,2903
regurgitation|2904,2917
)|2917,2918
<EOL>|2918,2919
LUNGS|2919,2924
-|2925,2926
CTA|2927,2930
bilat|2931,2936
,|2936,2937
no|2938,2940
r|2941,2942
/|2942,2943
rh|2943,2945
/|2945,2946
wh|2946,2948
,|2948,2949
good|2950,2954
air|2955,2958
movement|2959,2967
,|2967,2968
resp|2969,2973
<EOL>|2974,2975
unlabored|2975,2984
,|2984,2985
no|2986,2988
accessory|2989,2998
muscle|2999,3005
use|3006,3009
<EOL>|3009,3010
HEART|3010,3015
-|3016,3017
RRR|3018,3021
,|3021,3022
3|3023,3024
+|3024,3025
mid-systolic|3026,3038
murmur|3039,3045
loudest|3046,3053
at|3054,3056
LLS|3057,3060
border|3061,3067
,|3067,3068
<EOL>|3069,3070
radiates|3070,3078
to|3079,3081
axilla|3082,3088
,|3088,3089
nl|3090,3092
S1|3093,3095
-|3095,3096
S2|3096,3098
<EOL>|3098,3099
ABDOMEN|3099,3106
-|3107,3108
NABS|3109,3113
,|3113,3114
soft|3115,3119
/|3119,3120
NT|3120,3122
/|3122,3123
ND|3123,3125
,|3125,3126
no|3127,3129
masses|3130,3136
or|3137,3139
HSM|3140,3143
,|3143,3144
no|3145,3147
<EOL>|3148,3149
rebound|3149,3156
/|3156,3157
guarding|3157,3165
<EOL>|3165,3166
EXTREMITIES|3166,3177
-|3178,3179
WWP|3180,3183
,|3183,3184
no|3185,3187
c|3188,3189
/|3189,3190
c|3190,3191
/|3191,3192
e|3192,3193
,|3193,3194
2|3195,3196
+|3196,3197
peripheral|3198,3208
pulses|3209,3215
(|3216,3217
radials|3217,3224
,|3224,3225
DPs|3226,3229
)|3229,3230
<EOL>|3230,3231
NEURO|3231,3236
-|3237,3238
awake|3239,3244
,|3244,3245
A|3246,3247
&|3247,3248
Ox3|3248,3251
,|3251,3252
muscle|3253,3259
strength|3260,3268
_|3269,3270
_|3270,3271
_|3271,3272
b|3273,3274
/|3274,3275
l|3275,3276
.|3276,3277
<EOL>|3277,3278
.|3278,3279
<EOL>|3279,3280
DISCHARGE|3280,3289
EXAM|3290,3294
:|3294,3295
Unchanged|3296,3305
with|3306,3310
previous|3311,3319
,|3319,3320
except|3321,3327
for|3328,3331
the|3332,3335
<EOL>|3336,3337
following|3337,3346
:|3346,3347
<EOL>|3347,3348
VS|3348,3350
-|3351,3352
Temp|3353,3357
97|3358,3360
.|3360,3361
8F|3361,3363
,|3363,3364
BP|3365,3367
123|3368,3371
/|3371,3372
74|3372,3374
,|3374,3375
HR|3376,3378
82|3379,3381
,|3381,3382
R|3383,3384
16|3385,3387
,|3387,3388
O2|3389,3391
-|3391,3392
sat|3392,3395
98|3396,3398
%|3398,3399
RA|3400,3402
<EOL>|3402,3403
LUNGS|3403,3408
-|3409,3410
CTA|3411,3414
bilat|3415,3420
,|3420,3421
no|3422,3424
r|3425,3426
/|3426,3427
rh|3427,3429
/|3429,3430
wh|3430,3432
,|3432,3433
good|3434,3438
air|3439,3442
movement|3443,3451
,|3451,3452
resp|3453,3457
<EOL>|3458,3459
unlabored|3459,3468
,|3468,3469
no|3470,3472
accessory|3473,3482
muscle|3483,3489
use|3490,3493
<EOL>|3493,3494
HEART|3494,3499
-|3500,3501
RRR|3502,3505
,|3505,3506
3|3507,3508
+|3508,3509
mid-systolic|3510,3522
murmur|3523,3529
loudest|3530,3537
at|3538,3540
_|3541,3542
_|3542,3543
_|3543,3544
border|3545,3551
,|3551,3552
<EOL>|3553,3554
radiates|3554,3562
to|3563,3565
_|3566,3567
_|3567,3568
_|3568,3569
,|3569,3570
_|3571,3572
_|3572,3573
_|3573,3574
S1|3575,3577
-|3577,3578
S2|3578,3580
<EOL>|3580,3581
<EOL>|3581,3582
<EOL>|3583,3584
Pertinent|3584,3593
Results|3594,3601
:|3601,3602
<EOL>|3602,3603
ADMISSION|3603,3612
LABS|3613,3617
:|3617,3618
<EOL>|3618,3619
_|3619,3620
_|3620,3621
_|3621,3622
05|3623,3625
:|3625,3626
50PM|3626,3630
BLOOD|3631,3636
WBC|3637,3640
-|3640,3641
12|3641,3643
.|3643,3644
0|3644,3645
*|3645,3646
#|3646,3647
RBC|3648,3651
-|3651,3652
3|3652,3653
.|3653,3654
48|3654,3656
*|3656,3657
Hgb|3658,3661
-|3661,3662
11|3662,3664
.|3664,3665
4|3665,3666
*|3666,3667
Hct|3668,3671
-|3671,3672
32|3672,3674
.|3674,3675
6|3675,3676
*|3676,3677
<EOL>|3678,3679
MCV|3679,3682
-|3682,3683
94|3683,3685
MCH|3686,3689
-|3689,3690
32|3690,3692
.|3692,3693
7|3693,3694
*|3694,3695
MCHC|3696,3700
-|3700,3701
34.9|3701,3705
RDW|3706,3709
-|3709,3710
13.4|3710,3714
Plt|3715,3718
_|3719,3720
_|3720,3721
_|3721,3722
<EOL>|3722,3723
_|3723,3724
_|3724,3725
_|3725,3726
05|3727,3729
:|3729,3730
50PM|3730,3734
BLOOD|3735,3740
Neuts|3741,3746
-|3746,3747
76|3747,3749
.|3749,3750
5|3750,3751
*|3751,3752
Lymphs|3753,3759
-|3759,3760
17|3760,3762
.|3762,3763
3|3763,3764
*|3764,3765
Monos|3766,3771
-|3771,3772
5.2|3772,3775
<EOL>|3776,3777
Eos|3777,3780
-|3780,3781
0.7|3781,3784
Baso|3785,3789
-|3789,3790
0.4|3790,3793
<EOL>|3793,3794
_|3794,3795
_|3795,3796
_|3796,3797
05|3798,3800
:|3800,3801
50PM|3801,3805
BLOOD|3806,3811
Plt|3812,3815
_|3816,3817
_|3817,3818
_|3818,3819
<EOL>|3819,3820
_|3820,3821
_|3821,3822
_|3822,3823
05|3824,3826
:|3826,3827
50PM|3827,3831
BLOOD|3832,3837
Glucose|3838,3845
-|3845,3846
101|3846,3849
*|3849,3850
UreaN|3851,3856
-|3856,3857
15|3857,3859
Creat|3860,3865
-|3865,3866
0.7|3866,3869
Na|3870,3872
-|3872,3873
135|3873,3876
<EOL>|3877,3878
K|3878,3879
-|3879,3880
4.4|3880,3883
Cl|3884,3886
-|3886,3887
101|3887,3890
HCO3|3891,3895
-|3895,3896
26|3896,3898
AnGap|3899,3904
-|3904,3905
12|3905,3907
<EOL>|3907,3908
_|3908,3909
_|3909,3910
_|3910,3911
05|3912,3914
:|3914,3915
50PM|3915,3919
BLOOD|3920,3925
cTropnT|3926,3933
-|3933,3934
<|3934,3935
0|3935,3936
.|3936,3937
01|3937,3939
<EOL>|3939,3940
_|3940,3941
_|3941,3942
_|3942,3943
08|3944,3946
:|3946,3947
05AM|3947,3951
BLOOD|3952,3957
cTropnT|3958,3965
-|3965,3966
<|3966,3967
0.01|3967,3971
<EOL>|3971,3972
.|3972,3973
<EOL>|3973,3974
DISCHARGE|3974,3983
LABS|3984,3988
:|3988,3989
<EOL>|3989,3990
_|3990,3991
_|3991,3992
_|3992,3993
08|3994,3996
:|3996,3997
05AM|3997,4001
BLOOD|4002,4007
WBC|4008,4011
-|4011,4012
6.0|4012,4015
RBC|4016,4019
-|4019,4020
3|4020,4021
.|4021,4022
62|4022,4024
*|4024,4025
Hgb|4026,4029
-|4029,4030
11|4030,4032
.|4032,4033
8|4033,4034
*|4034,4035
Hct|4036,4039
-|4039,4040
34|4040,4042
.|4042,4043
1|4043,4044
*|4044,4045
<EOL>|4046,4047
MCV|4047,4050
-|4050,4051
94|4051,4053
MCH|4054,4057
-|4057,4058
32|4058,4060
.|4060,4061
7|4061,4062
*|4062,4063
MCHC|4064,4068
-|4068,4069
34.7|4069,4073
RDW|4074,4077
-|4077,4078
13.3|4078,4082
Plt|4083,4086
_|4087,4088
_|4088,4089
_|4089,4090
<EOL>|4090,4091
_|4091,4092
_|4092,4093
_|4093,4094
08|4095,4097
:|4097,4098
05AM|4098,4102
BLOOD|4103,4108
Plt|4109,4112
_|4113,4114
_|4114,4115
_|4115,4116
<EOL>|4116,4117
_|4117,4118
_|4118,4119
_|4119,4120
08|4121,4123
:|4123,4124
05AM|4124,4128
BLOOD|4129,4134
Glucose|4135,4142
-|4142,4143
100|4143,4146
UreaN|4147,4152
-|4152,4153
12|4153,4155
Creat|4156,4161
-|4161,4162
0.8|4162,4165
Na|4166,4168
-|4168,4169
136|4169,4172
<EOL>|4173,4174
K|4174,4175
-|4175,4176
4.4|4176,4179
Cl|4180,4182
-|4182,4183
101|4183,4186
HCO3|4187,4191
-|4191,4192
28|4192,4194
AnGap|4195,4200
-|4200,4201
11|4201,4203
<EOL>|4203,4204
_|4204,4205
_|4205,4206
_|4206,4207
08|4208,4210
:|4210,4211
05AM|4211,4215
BLOOD|4216,4221
Calcium|4222,4229
-|4229,4230
9.3|4230,4233
Phos|4234,4238
-|4238,4239
3.3|4239,4242
Mg|4243,4245
-|4245,4246
1.9|4246,4249
<EOL>|4249,4250
_|4250,4251
_|4251,4252
_|4252,4253
11|4254,4256
:|4256,4257
00AM|4257,4261
BLOOD|4262,4267
Iron|4268,4272
-|4272,4273
98|4273,4275
<EOL>|4275,4276
_|4276,4277
_|4277,4278
_|4278,4279
11|4280,4282
:|4282,4283
00AM|4283,4287
BLOOD|4288,4293
calTIBC|4294,4301
-|4301,4302
354|4302,4305
VitB12|4306,4312
-|4312,4313
1270|4313,4317
*|4317,4318
Folate|4319,4325
-|4325,4326
GREATER|4326,4333
<EOL>|4334,4335
TH|4335,4337
Ferritn|4338,4345
-|4345,4346
80|4346,4348
TRF|4349,4352
-|4352,4353
272|4353,4356
<EOL>|4356,4357
.|4357,4358
<EOL>|4358,4359
MICROBIOLOGY|4359,4371
:|4371,4372
<EOL>|4372,4373
_|4373,4374
_|4374,4375
_|4375,4376
Blood|4377,4382
Cx|4383,4385
:|4385,4386
Pending|4387,4394
<EOL>|4394,4395
_|4395,4396
_|4396,4397
_|4397,4398
Urine|4399,4404
Cx|4405,4407
:|4407,4408
pending|4409,4416
<EOL>|4416,4417
.|4417,4418
<EOL>|4418,4419
IMAGING|4419,4426
:|4426,4427
<EOL>|4427,4428
_|4428,4429
_|4429,4430
_|4430,4431
Video|4432,4437
swallow|4438,4445
study|4446,4451
:|4451,4452
Not|4453,4456
likely|4457,4463
aspiration|4464,4474
.|4474,4475
<EOL>|4476,4477
RECOMMENDATIONS|4477,4492
:|4492,4493
1.|4494,4496
PO|4497,4499
diet|4500,4504
of|4505,4507
thin|4508,4512
liquids|4513,4520
and|4521,4524
soft|4525,4529
solids|4530,4536
2|4537,4538
.|4538,4539
<EOL>|4540,4541
Aspiration|4541,4551
precautions|4552,4563
including|4564,4573
:|4573,4574
<EOL>|4575,4576
a|4576,4577
)|4577,4578
keep|4579,4583
solids|4584,4590
soft|4591,4595
and|4596,4599
moist|4600,4605
b|4607,4608
)|4608,4609
use|4610,4613
liquid|4614,4620
wash|4621,4625
to|4626,4628
clear|4629,4634
<EOL>|4635,4636
solids|4636,4642
as|4643,4645
needed|4646,4652
<EOL>|4652,4653
c|4654,4655
)|4655,4656
alternate|4657,4666
bites|4667,4672
and|4673,4676
sips|4677,4681
3.|4682,4684
Meds|4685,4689
whole|4690,4695
with|4696,4700
water|4701,4706
4.|4707,4709
Regular|4710,4717
<EOL>|4718,4719
oral|4719,4723
care|4724,4728
<EOL>|4728,4729
5.|4729,4731
Suggest|4732,4739
nutritional|4740,4751
supplements|4752,4763
at|4764,4766
home|4767,4771
given|4772,4777
reports|4778,4785
of|4786,4788
<EOL>|4789,4790
recent|4790,4796
weight|4797,4803
loss|4804,4808
.|4808,4809
<EOL>|4809,4810
<EOL>|4811,4812
Brief|4812,4817
Hospital|4818,4826
Course|4827,4833
:|4833,4834
<EOL>|4834,4835
Ms.|4835,4838
_|4839,4840
_|4840,4841
_|4841,4842
is|4843,4845
a|4846,4847
pleasant|4848,4856
_|4857,4858
_|4858,4859
_|4859,4860
w|4861,4862
/|4862,4863
a|4864,4865
h|4866,4867
/|4867,4868
o|4868,4869
aortic|4870,4876
regurgitation|4877,4890
,|4890,4891
<EOL>|4892,4893
hypothyroidism|4893,4907
,|4907,4908
Sjogrens|4909,4917
,|4917,4918
and|4919,4922
HTN|4923,4926
who|4927,4930
presents|4931,4939
as|4940,4942
a|4943,4944
transfer|4945,4953
<EOL>|4954,4955
from|4955,4959
_|4960,4961
_|4961,4962
_|4962,4963
after|4964,4969
a|4970,4971
syncopal|4972,4980
episode|4981,4988
on|4989,4991
_|4992,4993
_|4993,4994
_|4994,4995
AM|4996,4998
.|4998,4999
Upon|5000,5004
admission|5005,5014
,|5014,5015
<EOL>|5016,5017
she|5017,5020
was|5021,5024
hemodynamically|5025,5040
stable|5041,5047
,|5047,5048
but|5049,5052
was|5053,5056
found|5057,5062
to|5063,5065
have|5066,5070
<EOL>|5071,5072
asymptomatic|5072,5084
pyuria|5085,5091
,|5091,5092
cough|5093,5098
,|5098,5099
and|5100,5103
a|5104,5105
WBC|5106,5109
of|5110,5112
12.0|5113,5117
.|5117,5118
<EOL>|5118,5119
.|5119,5120
<EOL>|5120,5121
ACTIVE|5121,5127
ISSUES|5128,5134
:|5134,5135
<EOL>|5135,5136
.|5136,5137
<EOL>|5137,5138
#|5138,5139
Syncope|5139,5146
:|5146,5147
Pt|5148,5150
's|5150,5152
syncopal|5153,5161
episode|5162,5169
appears|5170,5177
to|5178,5180
be|5181,5183
c|5184,5185
/|5185,5186
w|5186,5187
vasovagal|5188,5197
<EOL>|5198,5199
syncope|5199,5206
,|5206,5207
likely|5208,5214
in|5215,5217
the|5218,5221
setting|5222,5229
of|5230,5232
her|5233,5236
asymptomatic|5237,5249
pyuria|5250,5256
.|5256,5257
She|5258,5261
<EOL>|5262,5263
also|5263,5267
had|5268,5271
a|5272,5273
_|5274,5275
_|5275,5276
_|5276,5277
in|5278,5280
which|5281,5286
her|5287,5290
Tn|5291,5293
's|5293,5295
were|5296,5300
negative|5301,5309
X2|5310,5312
and|5313,5316
EKG|5317,5320
's|5320,5322
<EOL>|5323,5324
were|5324,5328
c|5329,5330
/|5330,5331
w|5331,5332
and|5333,5336
unchanged|5337,5346
from|5347,5351
previous|5352,5360
.|5360,5361
She|5362,5365
was|5366,5369
hemodynamically|5370,5385
<EOL>|5386,5387
stable|5387,5393
and|5394,5397
received|5398,5406
fluids|5407,5413
and|5414,5417
bactrim|5418,5425
(|5426,5427
see|5427,5430
below|5431,5436
)|5436,5437
.|5437,5438
Given|5439,5444
her|5445,5448
<EOL>|5449,5450
h|5450,5451
/|5451,5452
o|5452,5453
aortic|5454,5460
regurgitation|5461,5474
,|5474,5475
an|5476,5478
Echo|5479,5483
was|5484,5487
ordered|5488,5495
but|5496,5499
will|5500,5504
be|5505,5507
<EOL>|5508,5509
obtained|5509,5517
by|5518,5520
the|5521,5524
pt|5525,5527
on|5528,5530
an|5531,5533
outpatient|5534,5544
basis|5545,5550
.|5550,5551
<EOL>|5551,5552
.|5552,5553
<EOL>|5553,5554
#|5554,5555
Pyuria|5555,5561
:|5561,5562
She|5563,5566
had|5567,5570
18|5571,5573
WBC|5574,5577
and|5578,5581
Lg|5582,5584
leuk|5585,5589
esterase|5590,5598
on|5599,5601
UA|5602,5604
on|5605,5607
admission|5608,5617
,|5617,5618
<EOL>|5619,5620
although|5620,5628
she|5629,5632
had|5633,5636
no|5637,5639
bacteria|5640,5648
on|5649,5651
UA|5652,5654
or|5655,5657
Sx|5658,5660
of|5661,5663
burning|5664,5671
/|5671,5672
dysuria|5672,5679
.|5679,5680
<EOL>|5681,5682
Given|5682,5687
her|5688,5691
syncopal|5692,5700
episode|5701,5708
in|5709,5711
the|5712,5715
setting|5716,5723
of|5724,5726
a|5727,5728
UTI|5729,5732
,|5732,5733
treatment|5734,5743
<EOL>|5744,5745
with|5745,5749
bactrim|5750,5757
was|5758,5761
started|5762,5769
in|5770,5772
the|5773,5776
ED|5777,5779
and|5780,5783
continued|5784,5793
for|5794,5797
a|5798,5799
total|5800,5805
of|5806,5808
<EOL>|5809,5810
4|5810,5811
days|5812,5816
.|5816,5817
<EOL>|5817,5818
.|5818,5819
<EOL>|5819,5820
#|5820,5821
Leukocytosis|5821,5833
:|5833,5834
Her|5835,5838
WBC|5839,5842
of|5843,5845
12.0|5846,5850
is|5851,5853
likely|5854,5860
in|5861,5863
the|5864,5867
setting|5868,5875
of|5876,5878
her|5879,5882
<EOL>|5883,5884
UTI|5884,5887
.|5887,5888
She|5889,5892
was|5893,5896
treated|5897,5904
with|5905,5909
PO|5910,5912
bactrim|5913,5920
as|5921,5923
above|5924,5929
.|5929,5930
<EOL>|5931,5932
.|5932,5933
<EOL>|5933,5934
INACTIVE|5934,5942
ISSUES|5943,5949
:|5949,5950
<EOL>|5950,5951
.|5951,5952
<EOL>|5952,5953
#|5953,5954
Anemia|5954,5960
:|5960,5961
Hct|5962,5965
_|5966,5967
_|5967,5968
_|5968,5969
is|5970,5972
32.6|5973,5977
,|5977,5978
slightly|5979,5987
down|5988,5992
from|5993,5997
baseline|5998,6006
of|6007,6009
~|6010,6011
35|6011,6013
.|6013,6014
<EOL>|6015,6016
Her|6016,6019
Iron|6020,6024
studies|6025,6032
,|6032,6033
B12|6034,6037
,|6037,6038
and|6039,6042
Folate|6043,6049
were|6050,6054
within|6055,6061
normal|6062,6068
limits|6069,6075
.|6075,6076
<EOL>|6076,6077
.|6077,6078
<EOL>|6078,6079
#|6079,6080
HTN|6080,6083
:|6083,6084
Her|6085,6088
home|6089,6093
lisinopril|6094,6104
was|6105,6108
decreased|6109,6118
to|6119,6121
10mg|6122,6126
PO|6127,6129
qday|6130,6134
,|6134,6135
in|6136,6138
the|6139,6142
<EOL>|6143,6144
setting|6144,6151
of|6152,6154
her|6155,6158
syncope|6159,6166
in|6167,6169
order|6170,6175
to|6176,6178
ensure|6179,6185
her|6186,6189
BP|6190,6192
does|6193,6197
not|6198,6201
drop|6202,6206
<EOL>|6207,6208
too|6208,6211
low|6212,6215
.|6215,6216
<EOL>|6216,6217
.|6217,6218
<EOL>|6218,6219
#|6219,6220
Hypothyroidism|6220,6234
:|6234,6235
continued|6236,6245
home|6246,6250
levothyroxin|6251,6263
.|6263,6264
<EOL>|6264,6265
.|6265,6266
<EOL>|6266,6267
TRANSITIONS|6267,6278
OF|6279,6281
CARE|6282,6286
:|6286,6287
<EOL>|6287,6288
-|6288,6289
_|6290,6291
_|6291,6292
_|6292,6293
Iron|6294,6298
studies|6299,6306
wnl|6307,6310
,|6310,6311
B12|6312,6315
1270|6316,6320
,|6320,6321
and|6322,6325
Folate|6326,6332
>|6333,6334
20|6334,6336
.|6336,6337
<EOL>|6337,6338
-|6338,6339
Pt|6340,6342
will|6343,6347
obtain|6348,6354
Echo|6355,6359
as|6360,6362
outpt|6363,6368
.|6368,6369
<EOL>|6369,6370
<EOL>|6371,6372
Medications|6372,6383
on|6384,6386
Admission|6387,6396
:|6396,6397
<EOL>|6397,6398
Lisinopril|6398,6408
20mg|6409,6413
PO|6414,6416
qday|6417,6421
<EOL>|6421,6422
Levothyroxine|6422,6435
50mcg|6436,6441
PO|6442,6444
qday|6445,6449
<EOL>|6449,6450
<EOL>|6450,6451
<EOL>|6452,6453
Discharge|6453,6462
Medications|6463,6474
:|6474,6475
<EOL>|6475,6476
1.|6476,6478
levothyroxine|6479,6492
50|6493,6495
mcg|6496,6499
Tablet|6500,6506
Sig|6507,6510
:|6510,6511
One|6512,6515
(|6516,6517
1|6517,6518
)|6518,6519
Tablet|6520,6526
PO|6527,6529
DAILY|6530,6535
<EOL>|6536,6537
(|6537,6538
Daily|6538,6543
)|6543,6544
.|6544,6545
<EOL>|6547,6548
2.|6548,6550
lisinopril|6551,6561
10|6562,6564
mg|6565,6567
Tablet|6568,6574
Sig|6575,6578
:|6578,6579
One|6580,6583
(|6584,6585
1|6585,6586
)|6586,6587
Tablet|6588,6594
PO|6595,6597
DAILY|6598,6603
(|6604,6605
Daily|6605,6610
)|6610,6611
.|6611,6612
<EOL>|6612,6613
Disp|6613,6617
:|6617,6618
*|6618,6619
30|6619,6621
Tablet|6622,6628
(|6628,6629
s|6629,6630
)|6630,6631
*|6631,6632
Refills|6633,6640
:|6640,6641
*|6641,6642
2|6642,6643
*|6643,6644
<EOL>|6644,6645
3.|6645,6647
sulfamethoxazole|6648,6664
-|6664,6665
trimethoprim|6665,6677
800|6678,6681
-|6681,6682
160|6682,6685
mg|6686,6688
Tablet|6689,6695
Sig|6696,6699
:|6699,6700
One|6701,6704
(|6705,6706
1|6706,6707
)|6707,6708
<EOL>|6709,6710
Tablet|6710,6716
PO|6717,6719
BID|6720,6723
(|6724,6725
2|6725,6726
times|6727,6732
a|6733,6734
day|6735,6738
)|6738,6739
for|6740,6743
2|6744,6745
days|6746,6750
.|6750,6751
<EOL>|6751,6752
Disp|6752,6756
:|6756,6757
*|6757,6758
4|6758,6759
Tablet|6760,6766
(|6766,6767
s|6767,6768
)|6768,6769
*|6769,6770
Refills|6771,6778
:|6778,6779
*|6779,6780
0|6780,6781
*|6781,6782
<EOL>|6782,6783
4.|6783,6785
Fish|6786,6790
Oil|6791,6794
Oral|6796,6800
<EOL>|6800,6801
5.|6801,6803
calcium|6804,6811
Oral|6813,6817
<EOL>|6817,6818
<EOL>|6818,6819
<EOL>|6820,6821
Discharge|6821,6830
Disposition|6831,6842
:|6842,6843
<EOL>|6843,6844
Home|6844,6848
<EOL>|6848,6849
<EOL>|6850,6851
Discharge|6851,6860
Diagnosis|6861,6870
:|6870,6871
<EOL>|6871,6872
Primary|6872,6879
diagnosis|6880,6889
:|6889,6890
<EOL>|6890,6891
Syncope|6891,6898
<EOL>|6898,6899
<EOL>|6899,6900
Secondary|6900,6909
diagnoses|6910,6919
:|6919,6920
<EOL>|6920,6921
Hypothyroidism|6921,6935
<EOL>|6935,6936
Hypertension|6936,6948
<EOL>|6948,6949
<EOL>|6949,6950
<EOL>|6951,6952
Discharge|6952,6961
Condition|6962,6971
:|6971,6972
<EOL>|6972,6973
Mental|6973,6979
Status|6980,6986
:|6986,6987
Clear|6988,6993
and|6994,6997
coherent|6998,7006
.|7006,7007
<EOL>|7007,7008
Level|7008,7013
of|7014,7016
Consciousness|7017,7030
:|7030,7031
Alert|7032,7037
and|7038,7041
interactive|7042,7053
.|7053,7054
<EOL>|7054,7055
Activity|7055,7063
Status|7064,7070
:|7070,7071
Ambulatory|7072,7082
-|7083,7084
Independent|7085,7096
.|7096,7097
<EOL>|7097,7098
<EOL>|7098,7099
<EOL>|7100,7101
Discharge|7101,7110
Instructions|7111,7123
:|7123,7124
<EOL>|7124,7125
Dear|7125,7129
Ms.|7130,7133
_|7134,7135
_|7135,7136
_|7136,7137
,|7137,7138
<EOL>|7138,7139
<EOL>|7139,7140
It|7140,7142
was|7143,7146
a|7147,7148
pleasure|7149,7157
providing|7158,7167
care|7168,7172
for|7173,7176
you|7177,7180
here|7181,7185
at|7186,7188
the|7189,7192
_|7193,7194
_|7194,7195
_|7195,7196
<EOL>|7197,7198
_|7198,7199
_|7199,7200
_|7200,7201
.|7201,7202
You|7204,7207
were|7208,7212
admitted|7213,7221
after|7222,7227
having|7228,7234
a|7235,7236
syncopal|7237,7245
<EOL>|7246,7247
(|7247,7248
fainting|7248,7256
)|7256,7257
episode|7258,7265
on|7266,7268
_|7269,7270
_|7270,7271
_|7271,7272
.|7272,7273
You|7275,7278
were|7279,7283
found|7284,7289
to|7290,7292
have|7293,7297
some|7298,7302
<EOL>|7303,7304
evidence|7304,7312
of|7313,7315
a|7316,7317
urinary|7318,7325
tract|7326,7331
infection|7332,7341
and|7342,7345
were|7346,7350
treated|7351,7358
with|7359,7363
an|7364,7366
<EOL>|7367,7368
antibiotic|7368,7378
called|7379,7385
Bactrim|7386,7393
.|7393,7394
Your|7396,7400
chest|7401,7406
x-ray|7407,7412
at|7413,7415
the|7416,7419
other|7420,7425
<EOL>|7426,7427
hospital|7427,7435
did|7436,7439
not|7440,7443
show|7444,7448
evidence|7449,7457
of|7458,7460
a|7461,7462
pneumonia|7463,7472
.|7472,7473
We|7475,7477
monitored|7478,7487
<EOL>|7488,7489
your|7489,7493
heart|7494,7499
rhythm|7500,7506
overnight|7507,7516
and|7517,7520
did|7521,7524
not|7525,7528
note|7529,7533
any|7534,7537
abnormalities|7538,7551
.|7551,7552
<EOL>|7554,7555
Your|7555,7559
electrocardiogram|7560,7577
did|7578,7581
not|7582,7585
show|7586,7590
any|7591,7594
changes|7595,7602
.|7602,7603
Your|7605,7609
blood|7610,7615
<EOL>|7616,7617
pressure|7617,7625
remained|7626,7634
stable|7635,7641
.|7641,7642
You|7644,7647
will|7648,7652
need|7653,7657
an|7658,7660
ultrasound|7661,7671
of|7672,7674
the|7675,7678
<EOL>|7679,7680
heart|7680,7685
for|7686,7689
further|7690,7697
evaluation|7698,7708
(|7709,7710
echocardiogram|7710,7724
)|7724,7725
,|7725,7726
but|7727,7730
this|7731,7735
can|7736,7739
be|7740,7742
<EOL>|7743,7744
done|7744,7748
after|7749,7754
you|7755,7758
leave|7759,7764
the|7765,7768
_|7769,7770
_|7770,7771
_|7771,7772
.|7772,7773
<EOL>|7774,7775
<EOL>|7775,7776
Your|7776,7780
condition|7781,7790
has|7791,7794
improved|7795,7803
and|7804,7807
you|7808,7811
can|7812,7815
be|7816,7818
discharged|7819,7829
to|7830,7832
home|7833,7837
.|7837,7838
<EOL>|7838,7839
<EOL>|7839,7840
The|7840,7843
following|7844,7853
changes|7854,7861
were|7862,7866
made|7867,7871
to|7872,7874
your|7875,7879
medications|7880,7891
:|7891,7892
<EOL>|7892,7893
<EOL>|7893,7894
NEW|7894,7897
:|7897,7898
<EOL>|7899,7900
-|7900,7901
Bactrim|7901,7908
double|7909,7915
-|7915,7916
strength|7916,7924
tab|7925,7928
,|7928,7929
1|7930,7931
tab|7932,7935
by|7936,7938
mouth|7939,7944
twice|7945,7950
daily|7951,7956
for|7957,7960
2|7961,7962
<EOL>|7963,7964
more|7964,7968
days|7969,7973
(|7974,7975
to|7975,7977
treat|7978,7983
urinary|7984,7991
tract|7992,7997
infection|7998,8007
)|8007,8008
<EOL>|8008,8009
<EOL>|8009,8010
CHANGED|8010,8017
:|8017,8018
<EOL>|8018,8019
-|8019,8020
DECREASED|8021,8030
Lisinopril|8031,8041
to|8042,8044
10mg|8045,8049
by|8050,8052
mouth|8053,8058
daily|8059,8064
<EOL>|8064,8065
<EOL>|8065,8066
Please|8066,8072
keep|8073,8077
your|8078,8082
follow|8083,8089
-|8089,8090
up|8090,8092
appointments|8093,8105
as|8106,8108
scheduled|8109,8118
below|8119,8124
.|8124,8125
We|8127,8129
<EOL>|8130,8131
are|8131,8134
also|8135,8139
working|8140,8147
to|8148,8150
schedule|8151,8159
your|8160,8164
echocardiogram|8165,8179
.|8179,8180
<EOL>|8180,8181
<EOL>|8181,8182
Of|8182,8184
note|8185,8189
,|8189,8190
while|8191,8196
you|8197,8200
were|8201,8205
here|8206,8210
you|8211,8214
had|8215,8218
a|8219,8220
video|8221,8226
swallow|8227,8234
study|8235,8240
that|8241,8245
<EOL>|8246,8247
did|8247,8250
not|8251,8254
show|8255,8259
evidence|8260,8268
that|8269,8273
you|8274,8277
are|8278,8281
aspirating|8282,8292
when|8293,8297
you|8298,8301
swallow|8302,8309
.|8309,8310
<EOL>|8312,8313
You|8313,8316
can|8317,8320
continue|8321,8329
to|8330,8332
eat|8333,8336
a|8337,8338
regular|8339,8346
diet|8347,8351
.|8351,8352
<EOL>|8352,8353
<EOL>|8354,8355
Followup|8355,8363
Instructions|8364,8376
:|8376,8377
<EOL>|8377,8378
_|8378,8379
_|8379,8380
_|8380,8381
<EOL>|8381,8382

