 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|159,166|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|159,166|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|169,178|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|169,178|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|169,178|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Body Substance|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|189,197|true|false|false|||recorded
Attribute|Clinical Attribute|SIMPLE_SEGMENT|217,226|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|217,226|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|217,226|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|230,235|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|SIMPLE_SEGMENT|230,235|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|230,235|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|SIMPLE_SEGMENT|238,247|true|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|238,247|true|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|256,271|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|262,271|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|262,271|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|262,271|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|273,287|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|273,287|false|false|false|||diverticulitis
Finding|Classification|SIMPLE_SEGMENT|290,295|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|296,304|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|296,304|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|308,326|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|317,326|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|317,326|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|317,326|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|317,326|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|317,326|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|332,344|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|332,362|false|false|false|C0585462;C5890124|Laparoscopic sigmoid colectomy;Laparoscopic-assisted sigmoid colectomy|laparoscopic sigmoid colectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|345,352|false|false|false|C0227391|Sigmoid colon|sigmoid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|345,362|false|false|false|C0192866|Sigmoid colectomy|sigmoid colectomy
Event|Event|SIMPLE_SEGMENT|353,362|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|353,362|false|false|false|C0009274|Colectomy|colectomy
Event|Event|SIMPLE_SEGMENT|367,374|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|367,377|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|367,393|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|367,393|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|378,385|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|378,385|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|378,393|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|386,393|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|420,427|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|420,427|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|420,427|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|420,427|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|420,430|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|441,455|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|441,455|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|469,478|false|false|false|||diagnosed
Event|Event|SIMPLE_SEGMENT|491,498|false|false|false|||reports
Finding|Idea or Concept|SIMPLE_SEGMENT|505,510|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|505,510|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|SIMPLE_SEGMENT|511,518|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|511,518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|511,518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|511,518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|511,521|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|523,526|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Attribute|Clinical Attribute|SIMPLE_SEGMENT|527,531|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|527,531|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|527,531|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|527,531|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|562,572|false|false|false|||prescribed
Finding|Idea or Concept|SIMPLE_SEGMENT|578,581|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|578,581|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|582,588|false|false|false|||course
Drug|Organic Chemical|SIMPLE_SEGMENT|592,597|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|592,597|false|false|false|C0701042|Cipro|Cipro
Drug|Organic Chemical|SIMPLE_SEGMENT|598,604|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|598,604|false|false|false|C0699678|Flagyl|Flagyl
Event|Event|SIMPLE_SEGMENT|618,627|false|false|false|||completed
Finding|Finding|SIMPLE_SEGMENT|650,654|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|SIMPLE_SEGMENT|661,670|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|661,675|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|671,675|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|671,675|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|671,675|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|671,675|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|676,684|false|false|false|||returned
Finding|Intellectual Product|SIMPLE_SEGMENT|694,698|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|705,714|false|false|false|||finishing
Drug|Antibiotic|SIMPLE_SEGMENT|715,725|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|726,732|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|737,744|true|false|false|||reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|748,754|true|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|748,754|true|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|748,754|true|false|false|C0027497|Nausea|nausea
Finding|Finding|SIMPLE_SEGMENT|748,766|true|false|false|C3843946|Nausea or vomiting|nausea or vomiting
Event|Event|SIMPLE_SEGMENT|758,766|true|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|758,766|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|780,784|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|780,784|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|788,796|false|false|false|||maintain
Event|Event|SIMPLE_SEGMENT|797,806|false|false|false|||hydration
Finding|Finding|SIMPLE_SEGMENT|797,806|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|SIMPLE_SEGMENT|797,806|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Event|Event|SIMPLE_SEGMENT|823,829|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|823,829|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|823,829|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|839,847|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|839,847|false|false|false|C0003618|Desire for food|appetite
Finding|Finding|SIMPLE_SEGMENT|857,865|false|false|false|C2984079|Somewhat|somewhat
Event|Event|SIMPLE_SEGMENT|866,875|false|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|866,875|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|917,922|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|917,932|false|false|false|C0011135|Defecation|bowel movements
Event|Event|SIMPLE_SEGMENT|923,932|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|923,932|false|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|937,944|false|false|false|||reports
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|960,964|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|965,970|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Event|Event|SIMPLE_SEGMENT|965,970|false|false|false|||brown
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|971,976|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|971,986|false|false|false|C0011135|Defecation|bowel movements
Event|Event|SIMPLE_SEGMENT|977,986|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|977,986|false|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|997,1005|true|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|997,1005|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|997,1005|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|1010,1018|false|false|false|||presents
Finding|Intellectual Product|SIMPLE_SEGMENT|1038,1044|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|direct
Event|Event|SIMPLE_SEGMENT|1045,1054|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1045,1054|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Functional Concept|SIMPLE_SEGMENT|1059,1069|false|false|false|C0205269|Unresponsive to Treatment|refractory
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1070,1073|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Finding|Sign or Symptom|SIMPLE_SEGMENT|1070,1078|false|false|false|C0238551|Left lower quadrant pain|LLQ pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1074,1078|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1074,1078|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1074,1078|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1074,1078|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1083,1103|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1088,1095|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1088,1095|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1088,1095|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1088,1095|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1088,1095|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1088,1103|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1096,1103|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1096,1103|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1096,1103|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1105,1119|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|1105,1119|false|false|false|||diverticulitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1120,1129|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|1120,1129|false|false|false|||Migraines
Finding|Functional Concept|SIMPLE_SEGMENT|1130,1134|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1135,1141|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1142,1152|false|false|false|C0007642|Cellulitis|cellulitis
Event|Event|SIMPLE_SEGMENT|1142,1152|false|false|false|||cellulitis
Finding|Finding|SIMPLE_SEGMENT|1142,1152|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Finding|Functional Concept|SIMPLE_SEGMENT|1155,1161|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1155,1169|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1162,1169|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1162,1169|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1162,1169|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1162,1169|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1175,1181|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1175,1181|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1175,1181|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1175,1181|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1175,1189|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1182,1189|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1182,1189|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1182,1189|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1182,1189|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1191,1197|false|false|false|||father
Finding|Conceptual Entity|SIMPLE_SEGMENT|1191,1197|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|1191,1197|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1207,1214|false|true|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|1207,1214|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|1217,1225|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1217,1225|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1217,1225|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1217,1225|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1217,1230|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1217,1230|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1226,1230|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1226,1230|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1226,1230|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1240,1249|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1240,1249|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|1250,1254|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1250,1254|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1250,1254|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Classification|SIMPLE_SEGMENT|1293,1296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|1293,1296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Finding|SIMPLE_SEGMENT|1298,1302|false|false|false|C5575035|Well (answer to question)|well
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1304,1307|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1304,1307|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1304,1307|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1304,1307|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1304,1307|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1304,1307|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1304,1307|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|1309,1310|false|false|false|||A
Event|Event|SIMPLE_SEGMENT|1317,1320|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1325,1326|true|false|false|||R
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1331,1335|true|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1331,1335|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Event|Event|SIMPLE_SEGMENT|1331,1335|true|false|false|||RESP
Drug|Organic Chemical|SIMPLE_SEGMENT|1337,1341|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|1337,1341|false|false|false|||CTAB
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1342,1345|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1342,1345|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|1342,1345|false|false|false|||ABD
Event|Event|SIMPLE_SEGMENT|1353,1363|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|1353,1363|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1353,1363|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1364,1367|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Event|Event|SIMPLE_SEGMENT|1368,1381|false|false|false|||inferolateral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1385,1394|false|false|false|C0041638|Umbilical structure|umbilicus
Event|Event|SIMPLE_SEGMENT|1417,1425|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|1417,1425|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|SIMPLE_SEGMENT|1429,1436|true|false|false|||rebound
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1437,1440|true|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|SIMPLE_SEGMENT|1437,1440|true|false|false|||EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|1437,1440|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1445,1450|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1445,1450|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1445,1450|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1473,1482|false|false|false|||RADIOLOGY
Finding|Finding|SIMPLE_SEGMENT|1473,1482|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Idea or Concept|SIMPLE_SEGMENT|1473,1482|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|1473,1482|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1473,1482|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|RADIOLOGY
Finding|Idea or Concept|SIMPLE_SEGMENT|1484,1489|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Intellectual Product|SIMPLE_SEGMENT|1484,1496|false|false|false|C0460114|Final report|Final Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1490,1496|false|false|false|C4255046||Report
Event|Event|SIMPLE_SEGMENT|1490,1496|false|false|false|||Report
Finding|Intellectual Product|SIMPLE_SEGMENT|1490,1496|false|false|false|C0684224|Report (document)|Report
Procedure|Health Care Activity|SIMPLE_SEGMENT|1490,1496|false|false|false|C0700287|Reporting|Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1497,1506|false|false|false|C0882057||CT PELVIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1497,1506|false|false|false|C0412628|Computed tomography of pelvis|CT PELVIS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1500,1506|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1500,1506|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1500,1506|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|SIMPLE_SEGMENT|1500,1506|false|false|false|||PELVIS
Finding|Finding|SIMPLE_SEGMENT|1500,1506|false|false|false|C0812455|Pelvis problem|PELVIS
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1509,1517|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|1542,1549|false|false|false|||MEDICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1542,1549|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Idea or Concept|SIMPLE_SEGMENT|1542,1549|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Intellectual Product|SIMPLE_SEGMENT|1542,1549|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1542,1549|false|false|false|C0199168|Medical service|MEDICAL
Finding|Finding|SIMPLE_SEGMENT|1542,1559|false|false|false|C4745084|Medical Condition|MEDICAL CONDITION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1550,1559|false|false|false|C3864998||CONDITION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1550,1559|false|false|false|C0012634|Disease|CONDITION
Event|Event|SIMPLE_SEGMENT|1550,1559|false|false|false|||CONDITION
Finding|Conceptual Entity|SIMPLE_SEGMENT|1550,1559|false|false|false|C1705253|Logical Condition|CONDITION
Finding|Idea or Concept|SIMPLE_SEGMENT|1565,1569|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|1565,1569|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|1570,1573|false|false|false|||old
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1585,1599|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|1585,1599|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|1601,1611|false|false|false|||increasing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1612,1615|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Finding|Sign or Symptom|SIMPLE_SEGMENT|1612,1620|false|false|false|C0694551|Right lower quadrant pain|RLQ pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1616,1620|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1616,1620|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1616,1620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1616,1620|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1622,1632|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|1622,1632|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|1622,1632|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|SIMPLE_SEGMENT|1634,1642|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|1634,1642|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1657,1671|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|1657,1671|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|1680,1688|false|false|false|||junction
Finding|Functional Concept|SIMPLE_SEGMENT|1696,1706|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1696,1712|false|false|false|C0227389|Descending colon|descending colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1696,1712|false|false|false|C0153435;C0496863|Benign neoplasm of descending colon;Malignant neoplasm of descending colon|descending colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1696,1730|false|false|false|C0391910|Descending colon and sigmoid colon|descending colon and sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1707,1712|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1707,1712|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1707,1712|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|1707,1712|false|false|false|C0750873|COLON PROBLEM|colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1707,1730|false|false|false|C0545860|colon and sigmoid colon|colon and sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1717,1724|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1717,1730|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1717,1730|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1725,1730|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1725,1730|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1725,1730|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|1725,1730|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|1725,1730|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|SIMPLE_SEGMENT|1732,1738|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1732,1738|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Finding|SIMPLE_SEGMENT|1740,1755|false|false|false|C5425894|Mildly enlarged|mildly enlarged
Event|Event|SIMPLE_SEGMENT|1747,1755|false|false|false|||enlarged
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1747,1755|false|false|false|C1293134|Enlargement procedure|enlarged
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1756,1771|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Finding|Body Substance|SIMPLE_SEGMENT|1772,1777|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1772,1783|false|false|false|C0024204|lymph nodes|lymph nodes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1772,1783|false|false|false|C0154054|benign neoplasm of lymph nodes|lymph nodes
Event|Event|SIMPLE_SEGMENT|1791,1799|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1791,1799|false|true|false|C4722408|Reactive Therapy|reactive
Event|Event|SIMPLE_SEGMENT|1805,1811|false|false|false|||nature
Finding|Functional Concept|SIMPLE_SEGMENT|1805,1811|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|1805,1811|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|SIMPLE_SEGMENT|1816,1823|true|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|1816,1823|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|1816,1823|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|1816,1823|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1816,1823|true|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|1837,1849|true|false|false|||contemplated
Event|Event|SIMPLE_SEGMENT|1853,1861|true|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|1853,1861|true|false|false|C1522577|follow-up|followup
Event|Event|SIMPLE_SEGMENT|1866,1877|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|1896,1902|false|false|false|||assess
Drug|Organic Chemical|SIMPLE_SEGMENT|1907,1915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1907,1915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|1907,1915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|1907,1915|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|1907,1915|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|1907,1915|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Event|SIMPLE_SEGMENT|1916,1926|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|1916,1926|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|1916,1926|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1937,1945|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|1937,1945|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|1937,1945|false|false|false|C2607943|findings aspects|findings
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1961,1966|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|1961,1966|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1961,1966|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|1967,1970|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1975,1978|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1975,1978|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1975,1978|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1985,1988|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1985,1988|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1985,1988|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1985,1988|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1994,1997|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1994,1997|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2005,2008|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2005,2008|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2005,2008|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2005,2008|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2005,2008|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2012,2015|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2012,2015|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2012,2015|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2012,2015|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2012,2015|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2012,2015|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2021,2025|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2021,2025|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2040,2043|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2060,2065|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2060,2065|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2060,2065|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2066,2069|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2077,2080|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2077,2080|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2077,2080|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2087,2090|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2087,2090|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2087,2090|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2087,2090|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2097,2100|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2097,2100|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2108,2111|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2108,2111|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2108,2111|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2108,2111|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2108,2111|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2115,2118|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2115,2118|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2115,2118|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2115,2118|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2115,2118|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2115,2118|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2124,2128|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2124,2128|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2143,2146|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2163,2168|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2163,2168|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2163,2168|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2169,2172|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2178,2181|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2178,2181|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2178,2181|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2188,2191|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2188,2191|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2188,2191|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2188,2191|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2197,2200|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2197,2200|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2208,2211|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2208,2211|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2208,2211|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2208,2211|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2208,2211|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2215,2218|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2215,2218|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2215,2218|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2215,2218|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2215,2218|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2215,2218|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2224,2228|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2224,2228|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2244,2247|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2264,2269|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2264,2269|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2264,2269|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2270,2273|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2290,2295|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2290,2295|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2290,2295|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2300,2303|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|2300,2303|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2300,2303|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2325,2330|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2325,2330|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2325,2330|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2335,2338|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|2335,2338|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2335,2338|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2360,2365|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2360,2365|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2360,2365|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|2360,2373|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2360,2373|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2360,2373|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2366,2373|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2366,2373|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2366,2373|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2366,2373|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2366,2373|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2366,2373|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2420,2424|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2420,2424|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2420,2424|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2449,2454|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2449,2454|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2449,2454|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|2449,2462|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2449,2462|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2449,2462|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2455,2462|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2455,2462|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2455,2462|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2455,2462|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2455,2462|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2455,2462|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2508,2512|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2508,2512|false|false|false|C0005367|Bicarbonates|HCO3
Event|Event|SIMPLE_SEGMENT|2508,2512|false|false|false|||HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2508,2512|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2537,2542|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2537,2542|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2537,2542|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2543,2546|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2543,2546|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|2543,2546|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|2543,2546|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|2543,2546|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|2543,2546|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|2543,2546|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2543,2546|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2551,2554|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2551,2554|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2551,2554|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2551,2554|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|2551,2554|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|2551,2554|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|2551,2554|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2562,2565|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|2562,2565|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|2562,2565|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|2562,2565|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2562,2565|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2571,2578|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|2571,2578|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2609,2614|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2609,2614|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2609,2614|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2615,2618|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2615,2618|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|2615,2618|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|2615,2618|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|2615,2618|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|2615,2618|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|2615,2618|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2615,2618|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2622,2625|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2622,2625|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2622,2625|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2622,2625|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|2622,2625|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|2622,2625|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|2622,2625|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2632,2635|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|2632,2635|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|2632,2635|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|2632,2635|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2632,2635|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2641,2648|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|2641,2648|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Event|Event|SIMPLE_SEGMENT|2641,2648|false|false|false|||AlkPhos
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2653,2660|false|false|false|C0002712|amylase|Amylase
Drug|Enzyme|SIMPLE_SEGMENT|2653,2660|false|false|false|C0002712|amylase|Amylase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2653,2660|false|false|false|C0002712|amylase|Amylase
Event|Event|SIMPLE_SEGMENT|2653,2660|false|false|false|||Amylase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2653,2660|false|false|false|C0201883|Amylase measurement|Amylase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2689,2694|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2689,2694|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2689,2694|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2689,2702|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2695,2702|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2695,2702|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2695,2702|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|2695,2702|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|2695,2702|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|2695,2702|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2695,2702|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2708,2715|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2708,2715|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2708,2715|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2708,2715|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|2708,2715|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|2708,2715|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|2708,2715|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2708,2715|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2749,2754|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2749,2754|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2749,2754|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2749,2762|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2755,2762|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2755,2762|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2755,2762|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|2755,2762|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|2755,2762|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|2755,2762|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2755,2762|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2767,2774|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2767,2774|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2767,2774|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2767,2774|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|2767,2774|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|2767,2774|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|2767,2774|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2767,2774|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2807,2812|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2807,2812|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2807,2812|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2813,2818|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|2813,2818|false|false|false|C0042313|vancomycin|Vanco
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2840,2844|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|SWAB
Drug|Substance|SIMPLE_SEGMENT|2840,2844|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|SWAB
Event|Event|SIMPLE_SEGMENT|2840,2844|false|false|false|||SWAB
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2840,2844|false|false|false|C0563454|Taking of swab|SWAB
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2849,2853|false|false|false|C1515974|Anatomic Site|Site
Finding|Intellectual Product|SIMPLE_SEGMENT|2849,2853|false|false|false|C1546778||Site
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2855,2862|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2855,2862|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2855,2862|true|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2855,2862|true|false|false|C0941288|Abdomen problem|ABDOMEN
Drug|Substance|SIMPLE_SEGMENT|2869,2874|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|SIMPLE_SEGMENT|2869,2874|true|false|false|||Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2869,2874|true|false|false|C1546638|Fluid Specimen Code|Fluid
Event|Event|SIMPLE_SEGMENT|2889,2893|true|false|false|||sent
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2898,2902|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|2898,2902|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2898,2902|true|false|false|C0563454|Taking of swab|swab
Event|Event|SIMPLE_SEGMENT|2903,2912|true|false|false|||transport
Finding|Cell Function|SIMPLE_SEGMENT|2903,2912|true|false|false|C0005528;C1519628;C1705822|Biological Transport;Molecular Transport;Transfer Technique|transport
Finding|Functional Concept|SIMPLE_SEGMENT|2903,2912|true|false|false|C0005528;C1519628;C1705822|Biological Transport;Molecular Transport;Transfer Technique|transport
Finding|Molecular Function|SIMPLE_SEGMENT|2903,2912|true|false|false|C0005528;C1519628;C1705822|Biological Transport;Molecular Transport;Transfer Technique|transport
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2903,2918|true|false|false|C1548752|Transport Media,|transport media
Anatomy|Tissue|SIMPLE_SEGMENT|2913,2918|false|false|false|C0162867;C1254021|Media layer;Tunica Media|media
Finding|Intellectual Product|SIMPLE_SEGMENT|2913,2918|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|media
Drug|Substance|SIMPLE_SEGMENT|2929,2935|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|2929,2935|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|2929,2935|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2929,2935|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|2955,2962|true|false|false|||syringe
Finding|Intellectual Product|SIMPLE_SEGMENT|2967,2973|true|false|false|C1546717||needle
Finding|Finding|SIMPLE_SEGMENT|2976,2979|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|2976,2979|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Event|Event|SIMPLE_SEGMENT|2984,2988|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|2984,2988|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|2984,2988|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Finding|SIMPLE_SEGMENT|2993,3000|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Finding|Pathologic Function|SIMPLE_SEGMENT|2993,3000|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3001,3004|false|false|false|C0220647|Carcinoma of unknown primary|cup
Event|Event|SIMPLE_SEGMENT|3001,3004|false|false|false|||cup
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3010,3020|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|3010,3020|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3010,3020|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3015,3020|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|3015,3020|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3015,3020|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|3022,3027|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|3060,3065|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|3060,3065|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|3060,3065|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|3070,3087|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|SIMPLE_SEGMENT|3089,3099|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|3089,3099|false|false|false|||LEUKOCYTES
Finding|Body Substance|SIMPLE_SEGMENT|3089,3099|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|SIMPLE_SEGMENT|3089,3099|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Event|Event|SIMPLE_SEGMENT|3128,3133|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|3128,3133|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|3128,3133|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|3138,3142|false|false|false|||GRAM
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3143,3151|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Event|Event|SIMPLE_SEGMENT|3143,3151|false|false|false|||POSITIVE
Finding|Classification|SIMPLE_SEGMENT|3143,3151|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|SIMPLE_SEGMENT|3143,3151|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Event|Event|SIMPLE_SEGMENT|3217,3225|false|false|false|||CLUSTERS
Drug|Substance|SIMPLE_SEGMENT|3229,3234|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|SIMPLE_SEGMENT|3229,3234|false|false|false|||FLUID
Finding|Intellectual Product|SIMPLE_SEGMENT|3229,3234|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3235,3242|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3235,3242|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3235,3242|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3235,3242|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3235,3242|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|3244,3249|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|3244,3249|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3262,3267|false|false|false|C0038160|Staphylococcal Infections|STAPH
Event|Event|SIMPLE_SEGMENT|3262,3267|false|false|false|||STAPH
Event|Event|SIMPLE_SEGMENT|3275,3279|false|false|false|||COAG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3275,3279|false|false|false|C0005790|Blood coagulation tests|COAG
Finding|Finding|SIMPLE_SEGMENT|3286,3294|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Finding|Intellectual Product|SIMPLE_SEGMENT|3286,3294|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Event|Event|SIMPLE_SEGMENT|3295,3301|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|3295,3301|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3295,3301|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|3295,3301|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|3295,3301|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3295,3301|false|false|false|C2911660|Growth action|GROWTH
Drug|Antibiotic|SIMPLE_SEGMENT|3304,3315|false|false|false|C0008947|clindamycin|CLINDAMYCIN
Drug|Organic Chemical|SIMPLE_SEGMENT|3304,3315|false|false|false|C0008947|clindamycin|CLINDAMYCIN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3316,3319|false|false|false|C0449201|PER (body structure)|PER
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3316,3319|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|PER
Event|Event|SIMPLE_SEGMENT|3316,3319|false|false|false|||PER
Finding|Functional Concept|SIMPLE_SEGMENT|3316,3319|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|PER
Finding|Gene or Genome|SIMPLE_SEGMENT|3316,3319|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|PER
Finding|Intellectual Product|SIMPLE_SEGMENT|3316,3319|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|PER
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3341,3348|false|false|false|C1764827;C1875400|ISOLATE COMPOUND;Isolate - microorganism|isolate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3341,3348|false|false|false|C1764827;C1875400|ISOLATE COMPOUND;Isolate - microorganism|isolate
Event|Event|SIMPLE_SEGMENT|3341,3348|false|false|false|||isolate
Event|Event|SIMPLE_SEGMENT|3352,3360|false|false|false|||presumed
Event|Event|SIMPLE_SEGMENT|3367,3376|false|false|false|||resistant
Finding|Functional Concept|SIMPLE_SEGMENT|3367,3376|false|true|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Finding|Idea or Concept|SIMPLE_SEGMENT|3367,3376|false|true|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3367,3376|false|true|false|C2827757|Antimicrobial Resistance Result|resistant
Finding|Functional Concept|SIMPLE_SEGMENT|3367,3379|false|true|false|C0332325|Resistant (qualifier value)|resistant to
Drug|Antibiotic|SIMPLE_SEGMENT|3380,3391|false|false|false|C0008947|clindamycin|clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|3380,3391|false|false|false|C0008947|clindamycin|clindamycin
Event|Event|SIMPLE_SEGMENT|3380,3391|false|false|false|||clindamycin
Event|Event|SIMPLE_SEGMENT|3415,3424|false|false|false|||detection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3415,3424|false|false|false|C1511790|Detection|detection
Finding|Functional Concept|SIMPLE_SEGMENT|3428,3437|false|false|false|C0205263|Induce (action)|inducible
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3438,3448|false|false|false|C1442099|Resistance|resistance
Event|Event|SIMPLE_SEGMENT|3438,3448|false|false|false|||resistance
Finding|Mental Process|SIMPLE_SEGMENT|3438,3448|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Physiologic Function|SIMPLE_SEGMENT|3438,3448|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Social Behavior|SIMPLE_SEGMENT|3438,3448|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3454,3471|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3464,3471|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3464,3471|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3464,3471|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3464,3471|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3464,3471|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|3503,3511|true|false|false|||ISOLATED
Event|Event|SIMPLE_SEGMENT|3517,3521|false|false|false|||ACID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3517,3526|false|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|3522,3526|false|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|3522,3526|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|3522,3526|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|3522,3526|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Activity|SIMPLE_SEGMENT|3527,3532|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Event|Event|SIMPLE_SEGMENT|3527,3532|false|false|false|||SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|3527,3532|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3527,3532|false|false|false|C0444186|Smear test|SMEAR
Finding|Idea or Concept|SIMPLE_SEGMENT|3534,3539|false|false|false|C1546485|Diagnosis Type - Final|Final
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3555,3564|true|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|3560,3564|true|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|3560,3564|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|3560,3564|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|3560,3564|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Event|SIMPLE_SEGMENT|3565,3572|true|false|false|||BACILLI
Event|Event|SIMPLE_SEGMENT|3573,3577|true|false|false|||SEEN
Finding|Intellectual Product|SIMPLE_SEGMENT|3581,3587|true|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Event|Activity|SIMPLE_SEGMENT|3588,3593|true|false|false|C1947932|Smear - instruction imperative|SMEAR
Event|Event|SIMPLE_SEGMENT|3588,3593|true|false|false|||SMEAR
Finding|Functional Concept|SIMPLE_SEGMENT|3588,3593|true|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3588,3593|true|false|false|C0444186|Smear test|SMEAR
Event|Event|SIMPLE_SEGMENT|3599,3603|false|false|false|||ACID
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3599,3608|false|false|false|C1318720|Acid fast stain|ACID FAST
Event|Event|SIMPLE_SEGMENT|3604,3608|false|false|false|||FAST
Finding|Finding|SIMPLE_SEGMENT|3604,3608|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|SIMPLE_SEGMENT|3604,3608|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|SIMPLE_SEGMENT|3604,3608|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3609,3616|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3609,3616|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3609,3616|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3609,3616|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3609,3616|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3641,3645|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|3641,3645|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|3641,3645|true|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3641,3645|true|false|false|C0563454|Taking of swab|swab
Finding|Intellectual Product|SIMPLE_SEGMENT|3657,3664|true|false|false|C3260738|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|optimal
Drug|Substance|SIMPLE_SEGMENT|3665,3673|true|false|false|C0370003|Specimen|specimen
Event|Event|SIMPLE_SEGMENT|3665,3673|true|false|false|||specimen
Finding|Body Substance|SIMPLE_SEGMENT|3665,3673|true|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|specimen
Finding|Functional Concept|SIMPLE_SEGMENT|3665,3673|true|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|specimen
Event|Activity|SIMPLE_SEGMENT|3678,3686|true|false|false|C0237820||recovery
Event|Event|SIMPLE_SEGMENT|3678,3686|true|false|false|||recovery
Finding|Organism Function|SIMPLE_SEGMENT|3678,3686|true|false|false|C2004454|Recovery - healing process|recovery
Event|Event|SIMPLE_SEGMENT|3691,3703|false|false|false|||mycobacteria
Event|Event|SIMPLE_SEGMENT|3725,3730|false|false|false|||fungi
Finding|Functional Concept|SIMPLE_SEGMENT|3725,3730|false|false|false|C0521033|Fungal|fungi
Finding|Classification|SIMPLE_SEGMENT|3735,3743|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|3735,3743|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3735,3743|false|false|false|C5237010|Expression Negative|negative
Finding|Classification|SIMPLE_SEGMENT|3735,3750|false|false|false|C4704700|Negative Results|negative result
Event|Event|SIMPLE_SEGMENT|3744,3750|false|false|false|||result
Finding|Finding|SIMPLE_SEGMENT|3744,3750|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|3744,3750|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|3744,3750|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Event|Event|SIMPLE_SEGMENT|3762,3773|false|false|false|||interpreted
Event|Event|SIMPLE_SEGMENT|3785,3792|false|false|false|||caution
Finding|Finding|SIMPLE_SEGMENT|3804,3812|false|false|false|C0332149|Possible|possible
Anatomy|Tissue|SIMPLE_SEGMENT|3813,3819|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|3813,3819|false|true|false|C1547928|Tissue Specimen Code|tissue
Event|Event|SIMPLE_SEGMENT|3820,3826|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|3820,3826|false|true|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|3820,3826|false|true|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3820,3826|false|true|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|3820,3826|false|true|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3830,3839|false|false|false|C1720922|Respiratory Aspiration|aspirated
Event|Event|SIMPLE_SEGMENT|3830,3839|false|false|false|||aspirated
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3830,3839|false|false|false|C0700198|Pulmonary aspiration|aspirated
Drug|Substance|SIMPLE_SEGMENT|3841,3846|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3841,3846|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|3863,3872|false|false|false|||submitted
Finding|Functional Concept|SIMPLE_SEGMENT|3878,3884|false|false|false|C0521033|Fungal|FUNGAL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3878,3892|false|false|false|C0200954|Mycology culture|FUNGAL CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3885,3892|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3885,3892|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3885,3892|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3885,3892|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3885,3892|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3918,3924|true|false|false|C2939457|Fungus Present|FUNGUS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3918,3933|true|false|false|C0427953|Specimen fungus isolated|FUNGUS ISOLATED
Event|Event|SIMPLE_SEGMENT|3925,3933|true|false|false|||ISOLATED
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3944,3948|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|3944,3948|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|3944,3948|true|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3944,3948|true|false|false|C0563454|Taking of swab|swab
Finding|Intellectual Product|SIMPLE_SEGMENT|3960,3967|true|false|false|C3260738|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|optimal
Drug|Substance|SIMPLE_SEGMENT|3968,3976|true|false|false|C0370003|Specimen|specimen
Event|Event|SIMPLE_SEGMENT|3968,3976|true|false|false|||specimen
Finding|Body Substance|SIMPLE_SEGMENT|3968,3976|true|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|specimen
Finding|Functional Concept|SIMPLE_SEGMENT|3968,3976|true|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|specimen
Event|Activity|SIMPLE_SEGMENT|3981,3989|true|false|false|C0237820||recovery
Event|Event|SIMPLE_SEGMENT|3981,3989|true|false|false|||recovery
Finding|Organism Function|SIMPLE_SEGMENT|3981,3989|true|false|false|C2004454|Recovery - healing process|recovery
Event|Event|SIMPLE_SEGMENT|3994,4006|false|false|false|||mycobacteria
Event|Event|SIMPLE_SEGMENT|4028,4033|false|false|false|||fungi
Finding|Functional Concept|SIMPLE_SEGMENT|4028,4033|false|false|false|C0521033|Fungal|fungi
Finding|Classification|SIMPLE_SEGMENT|4038,4046|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|4038,4046|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4038,4046|false|false|false|C5237010|Expression Negative|negative
Finding|Classification|SIMPLE_SEGMENT|4038,4053|false|false|false|C4704700|Negative Results|negative result
Event|Event|SIMPLE_SEGMENT|4047,4053|false|false|false|||result
Finding|Finding|SIMPLE_SEGMENT|4047,4053|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|4047,4053|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|4047,4053|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Event|Event|SIMPLE_SEGMENT|4065,4076|false|false|false|||interpreted
Event|Event|SIMPLE_SEGMENT|4088,4095|false|false|false|||caution
Finding|Finding|SIMPLE_SEGMENT|4107,4115|false|false|false|C0332149|Possible|possible
Anatomy|Tissue|SIMPLE_SEGMENT|4116,4122|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|4116,4122|false|true|false|C1547928|Tissue Specimen Code|tissue
Event|Event|SIMPLE_SEGMENT|4123,4129|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|4123,4129|false|true|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|4123,4129|false|true|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4123,4129|false|true|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4123,4129|false|true|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4133,4142|false|false|false|C1720922|Respiratory Aspiration|aspirated
Event|Event|SIMPLE_SEGMENT|4133,4142|false|false|false|||aspirated
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4133,4142|false|false|false|C0700198|Pulmonary aspiration|aspirated
Drug|Substance|SIMPLE_SEGMENT|4144,4149|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4144,4149|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|4166,4175|false|false|false|||submitted
Event|Event|SIMPLE_SEGMENT|4180,4189|false|false|false|||Pathology
Finding|Functional Concept|SIMPLE_SEGMENT|4180,4189|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|Pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|4180,4189|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|Pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4180,4189|false|false|false|C0919386|Pathology procedure|Pathology
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4180,4201|false|false|false|C4086729|Pathologic Examination|Pathology Examination
Event|Activity|SIMPLE_SEGMENT|4190,4201|false|false|false|C4321457|Examination|Examination
Event|Event|SIMPLE_SEGMENT|4190,4201|false|false|false|||Examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|4190,4201|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|Examination
Drug|Substance|SIMPLE_SEGMENT|4203,4211|false|false|false|C0370003|Specimen|SPECIMEN
Event|Event|SIMPLE_SEGMENT|4203,4211|false|false|false|||SPECIMEN
Finding|Body Substance|SIMPLE_SEGMENT|4203,4211|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Finding|Functional Concept|SIMPLE_SEGMENT|4203,4211|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4223,4230|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4223,4236|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4223,4236|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4231,4236|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4231,4236|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4231,4236|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|4231,4236|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|4231,4236|false|false|false|C0750873|COLON PROBLEM|colon
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4238,4247|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|4238,4247|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|4238,4247|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|4238,4247|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4238,4247|false|false|false|C0184661|Interventional procedure|Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4262,4271|false|false|false|C0945731||DIAGNOSIS
Event|Event|SIMPLE_SEGMENT|4262,4271|false|false|false|||DIAGNOSIS
Finding|Classification|SIMPLE_SEGMENT|4262,4271|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|SIMPLE_SEGMENT|4262,4271|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4262,4271|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4275,4282|false|false|false|C0227391|Sigmoid colon|Sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4275,4288|false|false|false|C0227391|Sigmoid colon|Sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4275,4288|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|Sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4283,4288|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4283,4288|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4283,4288|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|4283,4288|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|4283,4288|false|false|false|C0750873|COLON PROBLEM|colon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4300,4309|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4312,4319|false|false|false|C0009368|Colon structure (body structure)|Colonic
Finding|Functional Concept|SIMPLE_SEGMENT|4333,4343|false|false|false|C1300196|Organized|organizing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4344,4361|false|false|false|C0341363|Paracolic abscess|pericolic abscess
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4354,4361|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|4354,4361|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|4354,4361|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|4363,4373|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4363,4373|false|false|false|C0332290|Consistent with|consistent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4380,4401|false|false|false|C0341257|Perforated diverticulum|ruptured diverticulum
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4389,4401|false|false|false|C0012817|Diverticulum|diverticulum
Event|Event|SIMPLE_SEGMENT|4389,4401|false|false|false|||diverticulum
Finding|Intellectual Product|SIMPLE_SEGMENT|4389,4401|false|false|false|C1546602||diverticulum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4417,4437|false|false|false|C1184738|Set of regional lymph nodes|regional lymph nodes
Finding|Body Substance|SIMPLE_SEGMENT|4426,4431|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4426,4437|false|false|false|C0024204|lymph nodes|lymph nodes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4426,4437|false|false|false|C0154054|benign neoplasm of lymph nodes|lymph nodes
Finding|Functional Concept|SIMPLE_SEGMENT|4443,4452|true|false|false|C0439674|Intrinsic origin|intrinsic
Anatomy|Tissue|SIMPLE_SEGMENT|4453,4460|true|false|false|C0026724|Mucous Membrane|mucosal
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4461,4474|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|4461,4474|true|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|4461,4474|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|4475,4479|true|false|false|||seen
Event|Event|SIMPLE_SEGMENT|4481,4489|false|false|false|||Clinical
Finding|Intellectual Product|SIMPLE_SEGMENT|4481,4489|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|Clinical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4491,4505|false|false|false|C0012813|Diverticulitis|Diverticulitis
Event|Event|SIMPLE_SEGMENT|4491,4505|false|false|false|||Diverticulitis
Event|Event|SIMPLE_SEGMENT|4509,4518|false|false|false|||RADIOLOGY
Finding|Finding|SIMPLE_SEGMENT|4509,4518|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Idea or Concept|SIMPLE_SEGMENT|4509,4518|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|4509,4518|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4509,4518|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|RADIOLOGY
Finding|Idea or Concept|SIMPLE_SEGMENT|4520,4525|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Intellectual Product|SIMPLE_SEGMENT|4520,4532|false|false|false|C0460114|Final report|Final Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4526,4532|false|false|false|C4255046||Report
Event|Event|SIMPLE_SEGMENT|4526,4532|false|false|false|||Report
Finding|Intellectual Product|SIMPLE_SEGMENT|4526,4532|false|false|false|C0684224|Report (document)|Report
Procedure|Health Care Activity|SIMPLE_SEGMENT|4526,4532|false|false|false|C0700287|Reporting|Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4533,4543|false|false|false|C1644645||CT ABDOMEN
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4533,4543|false|false|false|C0412620|CT of abdomen|CT ABDOMEN
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4533,4554|false|false|false|C0202840|CT of abdomen with contrast|CT ABDOMEN W/CONTRAST
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4536,4543|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4536,4543|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|4536,4543|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4536,4543|false|false|false|C0941288|Abdomen problem|ABDOMEN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4546,4554|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|4546,4554|false|false|false|||CONTRAST
Event|Event|SIMPLE_SEGMENT|4569,4575|false|false|false|||Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|4569,4575|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Event|Event|SIMPLE_SEGMENT|4577,4581|false|false|false|||Rule
Finding|Functional Concept|SIMPLE_SEGMENT|4586,4598|true|true|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Finding|SIMPLE_SEGMENT|4586,4602|true|true|false|C3842127|Subcutaneous air|subcutaneous air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4599,4602|true|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4599,4602|true|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4599,4602|true|true|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4599,4602|true|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4599,4602|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4599,4602|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4599,4602|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Substance|SIMPLE_SEGMENT|4606,4611|true|true|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4606,4611|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4606,4611|true|true|false|C1546638|Fluid Specimen Code|fluid
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4613,4624|false|false|false|C4072741|IV contrast|IV contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4616,4624|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|4616,4624|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|4632,4639|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|4632,4639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|4632,4639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|4632,4639|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4667,4681|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|4667,4681|false|false|false|||diverticulitis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4684,4690|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|4684,4690|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|4684,4690|false|false|false|C1546481|What subject filter - Status|status
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4696,4708|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4696,4726|false|false|false|C0585462;C5890124|Laparoscopic sigmoid colectomy;Laparoscopic-assisted sigmoid colectomy|laparoscopic sigmoid colectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4709,4716|false|false|false|C0227391|Sigmoid colon|sigmoid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4709,4726|false|false|false|C0192866|Sigmoid colectomy|sigmoid colectomy
Event|Event|SIMPLE_SEGMENT|4717,4726|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4717,4726|false|false|false|C0009274|Colectomy|colectomy
Event|Event|SIMPLE_SEGMENT|4737,4747|false|false|false|||incisional
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4737,4747|false|false|false|C0184898|Surgical incisions|incisional
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4749,4757|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|4749,4757|false|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|4759,4763|false|false|false|||Rule
Finding|Functional Concept|SIMPLE_SEGMENT|4768,4780|true|true|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Finding|SIMPLE_SEGMENT|4768,4784|true|true|false|C3842127|Subcutaneous air|subcutaneous air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4781,4784|true|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4781,4784|true|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4781,4784|true|true|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4781,4784|true|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4781,4784|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4781,4784|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4781,4784|true|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Substance|SIMPLE_SEGMENT|4788,4793|true|true|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4788,4793|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4788,4793|true|true|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|4795,4805|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4795,4805|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4795,4805|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4810,4816|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4810,4816|false|false|false|C1546481|What subject filter - Status|Status
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4822,4829|false|false|false|C0227391|Sigmoid colon|sigmoid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4822,4839|false|false|false|C0192866|Sigmoid colectomy|sigmoid colectomy
Event|Event|SIMPLE_SEGMENT|4830,4839|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4830,4839|false|false|false|C0009274|Colectomy|colectomy
Event|Event|SIMPLE_SEGMENT|4853,4859|false|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|4853,4859|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|SIMPLE_SEGMENT|4879,4883|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|4879,4883|false|false|false|C0332296|Free of (attribute)|free
Finding|Finding|SIMPLE_SEGMENT|4884,4899|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Finding|Functional Concept|SIMPLE_SEGMENT|4884,4899|false|false|false|C1522583;C4760449|Intraperitoneal (intended site);Intraperitoneal Route of Administration|intraperitoneal
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4900,4903|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4900,4903|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4900,4903|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4900,4903|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4900,4903|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4900,4903|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4900,4903|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Substance|SIMPLE_SEGMENT|4908,4913|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4908,4913|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4908,4913|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4926,4932|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4926,4932|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4926,4932|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|4926,4932|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|4926,4932|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|4943,4949|false|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|4943,4949|false|false|false|C1561574|Amount class - Amount|amount
Finding|Functional Concept|SIMPLE_SEGMENT|4963,4975|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Finding|SIMPLE_SEGMENT|4963,4979|false|false|false|C3842127|Subcutaneous air|subcutaneous air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4976,4979|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4976,4979|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4976,4979|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4976,4979|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4976,4979|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4976,4979|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4976,4979|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4997,5002|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4997,5002|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4997,5026|true|false|false|C2332167|Lower anterior abdominal wall|lower anterior abdominal wall
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5003,5011|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5003,5026|true|false|false|C0230193|Anterior abdominal wall|anterior abdominal wall
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5012,5021|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5012,5026|true|false|false|C0836916|Abdominal wall structure|abdominal wall
Event|Event|SIMPLE_SEGMENT|5027,5037|true|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5027,5037|true|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5027,5042|true|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|5057,5063|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|5057,5063|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5057,5063|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|5073,5081|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5073,5081|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5073,5084|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Drug|Substance|SIMPLE_SEGMENT|5094,5099|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5094,5099|true|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5094,5099|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5100,5110|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|5100,5110|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|5100,5110|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|5100,5110|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5100,5110|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|5115,5120|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5121,5129|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5121,5136|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5121,5136|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|5160,5168|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|5190,5196|false|false|false|||office
Finding|Idea or Concept|SIMPLE_SEGMENT|5190,5196|false|false|false|C1549636|Address type - Office|office
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5213,5222|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|5213,5227|false|true|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5223,5227|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5223,5227|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5223,5227|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5223,5227|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|5228,5234|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5228,5234|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|5235,5242|false|true|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|5235,5242|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|5235,5242|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|5235,5242|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5247,5261|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|5247,5261|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|5262,5267|false|false|false|||flare
Finding|Finding|SIMPLE_SEGMENT|5262,5267|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|SIMPLE_SEGMENT|5262,5267|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|SIMPLE_SEGMENT|5280,5285|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|5280,5285|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|5280,5285|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|5298,5306|true|false|false|||remained
Event|Event|SIMPLE_SEGMENT|5308,5314|true|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|5308,5314|true|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|5336,5345|true|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|5336,5356|true|false|false|C0744727|Hematocrit decreased|decreased hematocrit
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5346,5356|true|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|SIMPLE_SEGMENT|5346,5356|true|false|false|||hematocrit
Finding|Finding|SIMPLE_SEGMENT|5346,5356|true|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5346,5356|true|false|false|C0018935|Hematocrit Measurement|hematocrit
Event|Event|SIMPLE_SEGMENT|5367,5374|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|5375,5380|false|false|false|C3714655|On IV|on IV
Drug|Organic Chemical|SIMPLE_SEGMENT|5381,5386|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5381,5386|false|false|false|C0701042|Cipro|Cipro
Event|Event|SIMPLE_SEGMENT|5381,5386|false|false|false|||Cipro
Drug|Organic Chemical|SIMPLE_SEGMENT|5389,5395|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5389,5395|false|false|false|C0699678|Flagyl|Flagyl
Event|Event|SIMPLE_SEGMENT|5389,5395|false|false|false|||Flagyl
Event|Event|SIMPLE_SEGMENT|5402,5405|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5402,5405|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5411,5414|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5411,5414|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|5411,5414|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|5411,5414|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5411,5414|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|5415,5424|false|false|false|||hydration
Finding|Finding|SIMPLE_SEGMENT|5415,5424|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|SIMPLE_SEGMENT|5415,5424|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5426,5430|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5426,5430|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5426,5430|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5426,5430|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5432,5441|false|false|false|||managment
Finding|Intellectual Product|SIMPLE_SEGMENT|5447,5453|false|false|false|C0031082|Periodicals|serial
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5454,5463|false|false|false|C0000726|Abdomen|abdominal
Event|Event|SIMPLE_SEGMENT|5464,5469|false|false|false|||exams
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5474,5477|false|false|false|C2713652|HDAC2 protein, human|HD2
Drug|Enzyme|SIMPLE_SEGMENT|5474,5477|false|false|false|C2713652|HDAC2 protein, human|HD2
Finding|Gene or Genome|SIMPLE_SEGMENT|5474,5477|false|false|false|C1706172|HDAC2 wt Allele|HD2
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5478,5481|false|false|false|C1438777;C1873129|HDAC7 protein, human;HDAC9 protein, human|HD7
Drug|Enzyme|SIMPLE_SEGMENT|5478,5481|false|false|false|C1438777;C1873129|HDAC7 protein, human;HDAC9 protein, human|HD7
Finding|Gene or Genome|SIMPLE_SEGMENT|5478,5481|false|false|false|C1422386;C3539637|HDAC9 gene;HDAC9 wt Allele|HD7
Event|Event|SIMPLE_SEGMENT|5486,5495|false|false|false|||underwent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5498,5501|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|5498,5501|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5502,5509|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|5505,5509|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5505,5509|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|5516,5524|false|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|5525,5538|false|false|false|||uncomplicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5540,5554|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|5540,5554|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|5560,5569|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|5579,5584|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|5595,5604|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|5595,5604|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|5595,5604|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5595,5604|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5595,5604|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|5606,5613|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|5606,5613|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5606,5613|false|false|false|C0040808|Treatment Protocols|regimen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5619,5628|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|5619,5633|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5629,5633|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5629,5633|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5629,5633|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5629,5633|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5634,5643|false|false|false|||responded
Finding|Finding|SIMPLE_SEGMENT|5644,5648|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|5655,5663|false|false|false|C0728755|Dilaudid|Dilaudid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5655,5663|false|false|false|C0728755|Dilaudid|Dilaudid
Event|Event|SIMPLE_SEGMENT|5655,5663|false|false|false|||Dilaudid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5694,5700|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|5694,5700|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|5694,5700|false|false|false|C0015733|Feces|stools
Event|Event|SIMPLE_SEGMENT|5706,5715|true|false|false|||continued
Event|Event|SIMPLE_SEGMENT|5719,5727|true|false|false|||ambulate
Finding|Finding|SIMPLE_SEGMENT|5719,5727|true|false|false|C4036205|Ambulate|ambulate
Event|Event|SIMPLE_SEGMENT|5737,5747|true|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|5737,5747|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Activity|SIMPLE_SEGMENT|5753,5760|true|false|false|C1705116|Refused|refused
Finding|Idea or Concept|SIMPLE_SEGMENT|5753,5760|true|false|false|C1548564|Refused - Completion Status for valid values|refused
Event|Event|SIMPLE_SEGMENT|5773,5783|true|false|false|||injections
Finding|Functional Concept|SIMPLE_SEGMENT|5773,5783|true|false|false|C1828121|Injection Route of Administration|injections
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5773,5783|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injections
Procedure|Health Care Activity|SIMPLE_SEGMENT|5785,5793|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5785,5793|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Event|Event|SIMPLE_SEGMENT|5795,5802|false|false|false|||options
Finding|Finding|SIMPLE_SEGMENT|5795,5802|false|false|true|C0683525;C1518601|Options;treatment options|options
Finding|Functional Concept|SIMPLE_SEGMENT|5795,5802|false|false|true|C0683525;C1518601|Options;treatment options|options
Event|Event|SIMPLE_SEGMENT|5808,5817|false|false|false|||discussed
Finding|Body Substance|SIMPLE_SEGMENT|5822,5829|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5822,5829|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5822,5829|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|5843,5850|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|SIMPLE_SEGMENT|5843,5850|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|5843,5850|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5843,5850|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Event|SIMPLE_SEGMENT|5852,5859|false|false|false|||planned
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5869,5872|true|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5869,5872|true|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5869,5872|true|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Event|Event|SIMPLE_SEGMENT|5869,5872|true|false|false|||TPN
Finding|Gene or Genome|SIMPLE_SEGMENT|5869,5872|true|false|false|C1420583;C3813711|TAPBP gene;TAPBP wt Allele|TPN
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5869,5872|true|false|false|C0030548|Parenteral Nutrition, Total|TPN
Event|Event|SIMPLE_SEGMENT|5875,5879|true|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5875,5879|true|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Event|Event|SIMPLE_SEGMENT|5888,5897|true|false|false|||indicated
Event|Event|SIMPLE_SEGMENT|5908,5915|false|false|false|||started
Drug|Food|SIMPLE_SEGMENT|5919,5925|false|false|false|C0218063|Ensure (product)|Ensure
Event|Event|SIMPLE_SEGMENT|5926,5937|false|false|false|||supplements
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5939,5956|false|false|false|C2972960||Operative consent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5949,5956|false|false|false|C2923685||consent
Event|Event|SIMPLE_SEGMENT|5949,5956|false|false|false|||consent
Finding|Idea or Concept|SIMPLE_SEGMENT|5949,5956|false|false|false|C1511481;C1554192;C5702721|ActClass - consent;Consent;Consent (record artifact)|consent
Finding|Intellectual Product|SIMPLE_SEGMENT|5949,5956|false|false|false|C1511481;C1554192;C5702721|ActClass - consent;Consent;Consent (record artifact)|consent
Event|Event|SIMPLE_SEGMENT|5958,5965|false|false|false|||labwork
Event|Event|SIMPLE_SEGMENT|5967,5970|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5967,5970|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|5975,5978|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|5975,5978|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5975,5978|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|5984,5993|false|false|false|||collected
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5997,6000|false|false|false|C1438985|HDAC8 protein, human|HD8
Drug|Enzyme|SIMPLE_SEGMENT|5997,6000|false|false|false|C1438985|HDAC8 protein, human|HD8
Finding|Gene or Genome|SIMPLE_SEGMENT|5997,6000|false|false|false|C3810557|HDAC8 wt Allele|HD8
Event|Event|SIMPLE_SEGMENT|6014,6017|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6014,6017|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Event|Event|SIMPLE_SEGMENT|6032,6039|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|6032,6039|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|6032,6039|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|6032,6039|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6032,6039|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|6041,6049|false|false|false|||Continue
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6055,6058|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6055,6058|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|6055,6058|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|6055,6058|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6055,6058|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|6061,6068|false|false|false|||Surgery
Finding|Finding|SIMPLE_SEGMENT|6061,6068|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|SIMPLE_SEGMENT|6061,6068|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|6061,6068|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6061,6068|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Event|SIMPLE_SEGMENT|6105,6111|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|6117,6130|false|false|false|||uncomplicated
Event|Event|SIMPLE_SEGMENT|6142,6150|false|false|false|||observed
Event|Event|SIMPLE_SEGMENT|6155,6159|false|false|false|||PACU
Event|Event|SIMPLE_SEGMENT|6165,6176|false|false|false|||transferred
Finding|Gene or Genome|SIMPLE_SEGMENT|6189,6193|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Event|Event|SIMPLE_SEGMENT|6194,6203|false|false|false|||Continued
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6209,6212|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6209,6212|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|6209,6212|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|6209,6212|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6209,6212|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|6214,6217|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6214,6217|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Event|Event|SIMPLE_SEGMENT|6223,6228|false|false|false|||foley
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6230,6233|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6230,6233|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Event|Event|SIMPLE_SEGMENT|6230,6233|false|false|false|||PCA
Finding|Finding|SIMPLE_SEGMENT|6230,6233|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|SIMPLE_SEGMENT|6230,6233|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|SIMPLE_SEGMENT|6230,6233|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6230,6233|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6238,6242|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6238,6242|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6238,6242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6238,6242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6238,6253|false|false|false|C0002766|Pain management (procedure)|pain management
Event|Event|SIMPLE_SEGMENT|6243,6253|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|6243,6253|false|true|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|6243,6253|false|true|false|C0376636|Disease Management|management
Drug|Organic Chemical|SIMPLE_SEGMENT|6269,6275|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6269,6275|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|SIMPLE_SEGMENT|6269,6275|false|false|false|||relief
Finding|Finding|SIMPLE_SEGMENT|6269,6275|false|false|false|C0564405|Feeling relief|relief
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6287,6295|false|false|false|C3870119;C3870120;C3870121;C3870126;C5886131||Reported
Event|Event|SIMPLE_SEGMENT|6287,6295|false|false|false|||Reported
Finding|Functional Concept|SIMPLE_SEGMENT|6287,6295|false|false|false|C0684224;C4319718;C5703234|Report (document);Reported;Reported Information|Reported
Finding|Idea or Concept|SIMPLE_SEGMENT|6287,6295|false|false|false|C0684224;C4319718;C5703234|Report (document);Reported;Reported Information|Reported
Finding|Intellectual Product|SIMPLE_SEGMENT|6287,6295|false|false|false|C0684224;C4319718;C5703234|Report (document);Reported;Reported Information|Reported
Procedure|Health Care Activity|SIMPLE_SEGMENT|6287,6295|false|false|false|C0700287|Reporting|Reported
Event|Event|SIMPLE_SEGMENT|6296,6302|false|false|false|||flatus
Finding|Sign or Symptom|SIMPLE_SEGMENT|6296,6302|false|false|false|C0016204|Flatulence|flatus
Event|Event|SIMPLE_SEGMENT|6319,6321|false|false|false|||BM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6323,6330|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6323,6330|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|6323,6330|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6346,6349|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6346,6349|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6346,6349|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|6346,6349|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|6346,6349|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|6346,6349|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|6346,6349|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6365,6370|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|6365,6377|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|6371,6377|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6371,6377|false|false|false|C0037709||sounds
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6391,6399|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6391,6399|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|6391,6399|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6391,6399|false|false|false|C0184898|Surgical incisions|incision
Event|Event|SIMPLE_SEGMENT|6406,6415|false|false|false|||increased
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6416,6424|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|6416,6424|false|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|6425,6434|false|false|false|||extending
Event|Event|SIMPLE_SEGMENT|6438,6443|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|6438,6443|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6448,6458|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|6448,6458|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|6448,6458|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6448,6458|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Event|Event|SIMPLE_SEGMENT|6459,6466|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|6472,6483|true|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|6472,6483|true|false|false|C2986411|Improvement|improvement
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6488,6493|true|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|6488,6493|true|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|6488,6493|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|6488,6493|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|6488,6493|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6499,6502|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6499,6502|false|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6499,6502|false|false|false|C1568891|HGS protein, human|hrs
Event|Event|SIMPLE_SEGMENT|6499,6502|false|false|false|||hrs
Finding|Gene or Genome|SIMPLE_SEGMENT|6499,6502|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Drug|Antibiotic|SIMPLE_SEGMENT|6504,6509|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|6504,6509|false|false|false|C0250482|Zosyn|Zosyn
Event|Event|SIMPLE_SEGMENT|6510,6515|false|false|false|||added
Event|Event|SIMPLE_SEGMENT|6519,6526|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|6519,6526|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6519,6526|false|false|false|C0040808|Treatment Protocols|regimen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6528,6532|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6528,6532|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6528,6532|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6534,6544|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|6534,6544|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6534,6544|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|6545,6553|false|false|false|||switched
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6560,6570|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|6560,6570|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6560,6570|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|6576,6580|false|false|false|||pump
Finding|Molecular Function|SIMPLE_SEGMENT|6576,6580|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Event|Event|SIMPLE_SEGMENT|6581,6588|false|false|false|||removed
Finding|Gene or Genome|SIMPLE_SEGMENT|6599,6603|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6599,6603|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|SIMPLE_SEGMENT|6604,6609|false|false|false|||spike
Drug|Antibiotic|SIMPLE_SEGMENT|6623,6634|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|6623,6634|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|6635,6642|false|false|false|||started
Anatomy|Cell|SIMPLE_SEGMENT|6644,6647|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|6684,6691|false|false|false|||Reports
Finding|Intellectual Product|SIMPLE_SEGMENT|6684,6691|false|false|false|C0684224|Report (document)|Reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|6684,6691|false|false|false|C0700287|Reporting|Reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6706,6712|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|6706,6712|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|6706,6712|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|SIMPLE_SEGMENT|6713,6719|false|false|false|C0206046|Zofran|zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6713,6719|false|false|false|C0206046|Zofran|zofran
Event|Event|SIMPLE_SEGMENT|6713,6719|false|false|false|||zofran
Event|Event|SIMPLE_SEGMENT|6728,6737|false|false|false|||effective
Drug|Organic Chemical|SIMPLE_SEGMENT|6739,6748|false|false|false|C0701017|Compazine|Compazine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6739,6748|false|false|false|C0701017|Compazine|Compazine
Event|Event|SIMPLE_SEGMENT|6739,6748|false|false|false|||Compazine
Event|Event|SIMPLE_SEGMENT|6749,6754|false|false|false|||added
Event|Event|SIMPLE_SEGMENT|6758,6765|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|6758,6765|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6758,6765|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|6771,6779|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|6771,6779|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|6771,6779|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|SIMPLE_SEGMENT|6781,6788|false|false|false|||effects
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6790,6793|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6790,6793|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|6790,6793|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|6790,6793|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6790,6793|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|6794,6803|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|6813,6822|false|false|false|||consulted
Drug|Antibiotic|SIMPLE_SEGMENT|6833,6843|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|6833,6843|false|false|false|||antibiotic
Event|Event|SIMPLE_SEGMENT|6845,6852|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|6845,6852|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6845,6852|false|false|false|C0040808|Treatment Protocols|regimen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6864,6871|true|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|6867,6871|true|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6867,6871|true|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6875,6878|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6875,6878|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Event|Event|SIMPLE_SEGMENT|6899,6908|true|false|false|||intra-abd
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6910,6918|true|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|6910,6918|true|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|6910,6918|true|false|false|C2607943|findings aspects|findings
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6920,6925|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|SIMPLE_SEGMENT|6920,6925|false|false|false|||Wound
Finding|Body Substance|SIMPLE_SEGMENT|6920,6925|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|6920,6925|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|6920,6925|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Event|Event|SIMPLE_SEGMENT|6926,6932|false|false|false|||opened
Event|Event|SIMPLE_SEGMENT|6952,6960|false|false|false|||Cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|6952,6960|false|true|false|C0010453|Culture (Anthropological)|Cultures
Drug|Substance|SIMPLE_SEGMENT|6972,6977|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6972,6977|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6972,6977|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|6978,6982|false|false|false|||sent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6991,6995|false|false|false|C1515974|Anatomic Site|Site
Finding|Intellectual Product|SIMPLE_SEGMENT|6991,6995|false|false|false|C1546778||Site
Event|Event|SIMPLE_SEGMENT|6996,7002|false|false|false|||packed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7012,7020|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|SIMPLE_SEGMENT|7012,7020|false|false|false|||dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7012,7020|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|7012,7020|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|7012,7020|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7012,7020|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7022,7032|false|false|false|C0009450|Communicable Diseases|Infectious
Event|Event|SIMPLE_SEGMENT|7022,7032|false|false|false|||Infectious
Event|Event|SIMPLE_SEGMENT|7034,7042|false|false|false|||reaction
Finding|Functional Concept|SIMPLE_SEGMENT|7034,7042|false|false|false|C0443286|Reaction|reaction
Finding|Finding|SIMPLE_SEGMENT|7043,7049|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7043,7049|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7054,7057|false|true|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|GAS
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|7054,7057|false|true|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|GAS
Drug|Substance|SIMPLE_SEGMENT|7054,7057|false|true|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|GAS
Event|Event|SIMPLE_SEGMENT|7054,7057|false|false|false|||GAS
Finding|Gene or Genome|SIMPLE_SEGMENT|7054,7057|false|true|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|GAS
Finding|Intellectual Product|SIMPLE_SEGMENT|7054,7057|false|true|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|GAS
Finding|Molecular Function|SIMPLE_SEGMENT|7054,7057|false|true|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|GAS
Finding|Sign or Symptom|SIMPLE_SEGMENT|7054,7057|false|true|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|GAS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7061,7075|false|false|false|C0374989|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|staphylococcus
Event|Event|SIMPLE_SEGMENT|7061,7075|false|false|false|||staphylococcus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7061,7082|false|false|false|C1318973|Staphylococcus aureus infection|staphylococcus aureus
Event|Event|SIMPLE_SEGMENT|7076,7082|false|false|false|||aureus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7084,7089|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7084,7089|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|7084,7089|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7084,7089|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|7084,7089|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|7084,7089|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Body Substance|SIMPLE_SEGMENT|7084,7094|false|false|false|C3669207|Nasal swab (specimen)|Nasal swab
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7084,7094|false|false|false|C4318939|Nasal Swab Test|Nasal swab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7090,7094|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|7090,7094|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|7090,7094|false|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7090,7094|false|false|false|C0563454|Taking of swab|swab
Event|Event|SIMPLE_SEGMENT|7107,7116|false|false|false|||collected
Event|Event|SIMPLE_SEGMENT|7119,7123|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|7127,7132|false|false|false|||Micro
Finding|Conceptual Entity|SIMPLE_SEGMENT|7127,7132|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|SIMPLE_SEGMENT|7127,7132|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7127,7132|false|false|false|C0085672|Microbiology procedure|Micro
Drug|Antibiotic|SIMPLE_SEGMENT|7134,7145|false|false|false|C0008947|clindamycin|Clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|7134,7145|false|false|false|C0008947|clindamycin|Clindamycin
Event|Event|SIMPLE_SEGMENT|7149,7154|false|false|false|||added
Event|Event|SIMPLE_SEGMENT|7159,7166|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|7159,7166|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7159,7166|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|7168,7176|false|false|false|||Cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|7168,7176|false|false|false|C0010453|Culture (Anthropological)|Cultures
Event|Event|SIMPLE_SEGMENT|7182,7190|false|false|false|||followed
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7196,7201|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|7196,7201|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|7196,7201|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|7196,7201|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|7196,7201|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|7202,7209|false|false|false|||checked
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7223,7226|false|false|false|C1506708|MAX protein, human|max
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7223,7226|false|false|false|C1506708|MAX protein, human|max
Event|Event|SIMPLE_SEGMENT|7223,7226|false|false|false|||max
Finding|Finding|SIMPLE_SEGMENT|7223,7226|false|false|false|C0919516;C0919551;C4760036|MAX gene;Max (cigarettes);Oncogene MAX|max
Finding|Gene or Genome|SIMPLE_SEGMENT|7223,7226|false|false|false|C0919516;C0919551;C4760036|MAX gene;Max (cigarettes);Oncogene MAX|max
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7243,7253|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7243,7253|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7243,7253|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7243,7253|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7243,7253|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|7254,7259|false|false|false|||noted
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7279,7284|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|7279,7284|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|7279,7284|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|7279,7284|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7279,7292|false|false|false|C0855657|Wound Culture|wound culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7285,7292|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7285,7292|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7285,7292|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7285,7292|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7285,7292|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Finding|SIMPLE_SEGMENT|7285,7301|false|false|false|C0159125|Culture positive|culture positive
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7293,7301|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|7293,7301|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|7293,7301|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|7293,7301|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|7293,7305|false|false|false|C1446409|Positive|positive for
Event|Event|SIMPLE_SEGMENT|7306,7310|false|false|false|||MSSA
Finding|Finding|SIMPLE_SEGMENT|7306,7310|false|false|false|C2355591|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|MSSA
Drug|Antibiotic|SIMPLE_SEGMENT|7315,7324|false|false|false|C0027324|nafcillin|Nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|7315,7324|false|false|false|C0027324|nafcillin|Nafcillin
Event|Event|SIMPLE_SEGMENT|7315,7324|false|false|false|||Nafcillin
Event|Event|SIMPLE_SEGMENT|7325,7330|false|false|false|||added
Event|Event|SIMPLE_SEGMENT|7337,7346|false|false|false|||continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7358,7363|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|7358,7363|false|false|false|C0042313|vancomycin|Vanco
Event|Event|SIMPLE_SEGMENT|7358,7363|false|false|false|||Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|7366,7371|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|7366,7371|false|false|false|C0250482|Zosyn|Zosyn
Event|Event|SIMPLE_SEGMENT|7372,7384|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|7392,7400|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|7392,7400|false|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|7402,7410|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|7402,7410|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|7402,7410|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7402,7410|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7416,7421|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7416,7421|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|7416,7421|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7416,7421|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|7416,7421|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|7416,7421|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Body Substance|SIMPLE_SEGMENT|7416,7426|false|false|false|C3669207|Nasal swab (specimen)|Nasal swab
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7416,7426|false|false|false|C4318939|Nasal Swab Test|Nasal swab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7422,7426|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|7422,7426|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|7422,7426|false|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7422,7426|false|false|false|C0563454|Taking of swab|swab
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7431,7436|false|false|false|C0038160|Staphylococcal Infections|Staph
Event|Event|SIMPLE_SEGMENT|7431,7436|false|false|false|||Staph
Event|Event|SIMPLE_SEGMENT|7437,7445|false|false|false|||cultured
Event|Event|SIMPLE_SEGMENT|7446,7455|false|false|false|||collected
Finding|Body Substance|SIMPLE_SEGMENT|7457,7464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7457,7464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7457,7464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7466,7473|false|false|false|||reports
Finding|Intellectual Product|SIMPLE_SEGMENT|7466,7473|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|7466,7473|false|false|false|C0700287|Reporting|reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7474,7480|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|7474,7480|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7474,7480|false|false|false|C0027497|Nausea|nausea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7481,7486|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|7487,7494|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|7487,7494|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|7487,7494|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|7500,7506|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|7500,7506|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|7517,7523|false|false|false|||eating
Event|Event|SIMPLE_SEGMENT|7531,7537|false|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|7531,7537|false|false|false|C1561574|Amount class - Amount|amount
Drug|Food|SIMPLE_SEGMENT|7549,7553|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|7549,7553|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7549,7553|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|SIMPLE_SEGMENT|7549,7553|false|false|false|||food
Event|Event|SIMPLE_SEGMENT|7559,7568|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7559,7568|false|false|false|C0549178|Continuous|continued
Event|Event|SIMPLE_SEGMENT|7569,7575|false|false|false|||flatus
Finding|Sign or Symptom|SIMPLE_SEGMENT|7569,7575|false|false|false|C0016204|Flatulence|flatus
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7580,7586|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|SIMPLE_SEGMENT|7580,7586|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Event|Event|SIMPLE_SEGMENT|7580,7586|false|false|false|||liquid
Finding|Finding|SIMPLE_SEGMENT|7580,7586|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7580,7586|false|false|false|C0301571|Liquid diet|liquid
Finding|Body Substance|SIMPLE_SEGMENT|7580,7592|false|false|false|C1550307;C2129214|Liquid Stool substance;Loose stool|liquid stool
Finding|Sign or Symptom|SIMPLE_SEGMENT|7580,7592|false|false|false|C1550307;C2129214|Liquid Stool substance;Loose stool|liquid stool
Event|Event|SIMPLE_SEGMENT|7587,7592|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|7587,7592|false|false|false|C0015733|Feces|stool
Event|Event|SIMPLE_SEGMENT|7594,7604|false|false|false|||production
Event|Occupational Activity|SIMPLE_SEGMENT|7594,7604|false|false|false|C0033268|production|production
Finding|Intellectual Product|SIMPLE_SEGMENT|7594,7604|false|false|false|C1548180|Production Processing ID|production
Event|Event|SIMPLE_SEGMENT|7606,7615|false|false|false|||Continues
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7621,7624|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7621,7624|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|7621,7624|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|7621,7624|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7621,7624|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7641,7651|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7641,7651|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|7641,7651|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7641,7651|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7641,7651|false|false|false|C0201975|Creatinine measurement|Creatinine
Finding|Body Substance|SIMPLE_SEGMENT|7670,7675|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|7670,7675|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|7670,7675|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7670,7682|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7670,7682|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|SIMPLE_SEGMENT|7676,7682|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|7676,7682|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|7676,7682|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|7684,7694|false|false|false|||Ambulating
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7710,7713|false|false|false|C5816720|Isolated lipoma of filum terminale|LFT
Event|Event|SIMPLE_SEGMENT|7710,7713|false|false|false|||LFT
Finding|Gene or Genome|SIMPLE_SEGMENT|7710,7713|false|false|false|C1537580|LIX1 gene|LFT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7710,7713|false|false|false|C0023901|Liver Function Tests|LFT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7710,7715|false|false|false|C0023901|Liver Function Tests|LFT's
Event|Event|SIMPLE_SEGMENT|7726,7734|false|false|false|||elevated
Finding|Finding|SIMPLE_SEGMENT|7738,7742|false|false|false|C5575035|Well (answer to question)|well
Drug|Antibiotic|SIMPLE_SEGMENT|7754,7765|false|false|false|C0008947|clindamycin|Clindamycin
Drug|Organic Chemical|SIMPLE_SEGMENT|7754,7765|false|false|false|C0008947|clindamycin|Clindamycin
Event|Event|SIMPLE_SEGMENT|7754,7765|false|false|false|||Clindamycin
Event|Event|SIMPLE_SEGMENT|7766,7778|false|false|false|||discontinued
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7786,7793|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7786,7793|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7786,7793|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7786,7793|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7786,7793|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7794,7804|false|false|false|C1442099|Resistance|resistance
Event|Event|SIMPLE_SEGMENT|7794,7804|false|false|false|||resistance
Finding|Mental Process|SIMPLE_SEGMENT|7794,7804|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Physiologic Function|SIMPLE_SEGMENT|7794,7804|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Social Behavior|SIMPLE_SEGMENT|7794,7804|false|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Drug|Antibiotic|SIMPLE_SEGMENT|7807,7816|false|false|false|C0027324|nafcillin|Nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|7807,7816|false|false|false|C0027324|nafcillin|Nafcillin
Event|Event|SIMPLE_SEGMENT|7807,7816|false|false|false|||Nafcillin
Event|Event|SIMPLE_SEGMENT|7817,7826|false|false|false|||continued
Finding|Body Substance|SIMPLE_SEGMENT|7828,7835|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7828,7835|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7828,7835|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7838,7844|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|7838,7844|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|7838,7844|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|7845,7853|false|false|false|||contiues
Event|Event|SIMPLE_SEGMENT|7857,7864|false|false|false|||improve
Event|Event|SIMPLE_SEGMENT|7875,7883|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|7875,7883|false|false|false|C0277797|Apyrexial|afebrile
Finding|Finding|SIMPLE_SEGMENT|7885,7898|false|false|false|C0750394|White blood cell count decreased|decreased WBC
Anatomy|Cell|SIMPLE_SEGMENT|7895,7898|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|7895,7898|false|false|false|||WBC
Finding|Finding|SIMPLE_SEGMENT|7904,7912|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|7904,7912|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7913,7923|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|7913,7923|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|7913,7923|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7928,7933|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|7928,7933|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|7928,7933|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|7928,7933|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|7928,7933|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7944,7952|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|7944,7952|false|false|false|||erythema
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7954,7957|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7954,7957|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|7954,7957|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|7954,7957|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7954,7957|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|7958,7966|false|false|false|||switched
Event|Activity|SIMPLE_SEGMENT|7970,7981|false|false|false|C0024501|Maintenance|maintenance
Event|Event|SIMPLE_SEGMENT|7970,7981|false|false|false|||maintenance
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7990,7995|true|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7990,7995|true|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|7990,7995|true|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7990,7995|true|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|7990,7995|true|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|7990,7995|true|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Body Substance|SIMPLE_SEGMENT|7990,8000|true|false|false|C3669207|Nasal swab (specimen)|Nasal swab
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7990,8000|true|false|false|C4318939|Nasal Swab Test|Nasal swab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7996,8000|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|SIMPLE_SEGMENT|7996,8000|true|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|SIMPLE_SEGMENT|7996,8000|true|false|false|||swab
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7996,8000|true|false|false|C0563454|Taking of swab|swab
Event|Event|SIMPLE_SEGMENT|8004,8010|true|false|false|||growth
Finding|Finding|SIMPLE_SEGMENT|8004,8010|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8004,8010|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|SIMPLE_SEGMENT|8004,8010|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|SIMPLE_SEGMENT|8004,8010|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8004,8010|true|false|false|C2911660|Growth action|growth
Event|Event|SIMPLE_SEGMENT|8012,8021|false|false|false|||Continues
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8022,8025|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8022,8025|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|8022,8025|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|8022,8025|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8022,8025|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Drug|Antibiotic|SIMPLE_SEGMENT|8028,8037|false|false|false|C0027324|nafcillin|Nafcillin
Drug|Organic Chemical|SIMPLE_SEGMENT|8028,8037|false|false|false|C0027324|nafcillin|Nafcillin
Event|Event|SIMPLE_SEGMENT|8039,8047|false|false|false|||Improved
Event|Event|SIMPLE_SEGMENT|8052,8058|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|8052,8058|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|8052,8058|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|8060,8069|false|false|false|||Continues
Event|Event|SIMPLE_SEGMENT|8075,8085|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|8075,8085|false|false|false|C5441521|Complaint (finding)|complaints
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8102,8108|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|8102,8108|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8102,8108|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|8111,8120|false|false|false|||improving
Event|Event|SIMPLE_SEGMENT|8131,8141|false|false|false|||responsive
Finding|Functional Concept|SIMPLE_SEGMENT|8131,8141|false|false|false|C0205342|Responsive|responsive
Drug|Organic Chemical|SIMPLE_SEGMENT|8145,8154|false|false|false|C0701017|Compazine|Compazine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8145,8154|false|false|false|C0701017|Compazine|Compazine
Event|Event|SIMPLE_SEGMENT|8145,8154|false|false|false|||Compazine
Event|Event|SIMPLE_SEGMENT|8191,8199|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|8191,8199|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|SIMPLE_SEGMENT|8207,8216|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8207,8216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8207,8216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8207,8216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8207,8216|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|8217,8220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8217,8220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8222,8232|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|8222,8232|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|8222,8232|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|8222,8232|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8222,8232|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|SIMPLE_SEGMENT|8233,8242|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|8246,8254|false|false|false|||decrease
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8272,8282|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|8272,8282|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|8272,8282|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|8272,8282|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8272,8282|false|false|false|C0201975|Creatinine measurement|Creatinine
Finding|Finding|SIMPLE_SEGMENT|8272,8288|false|false|false|C0428279|Finding of creatinine level|Creatinine level
Event|Event|SIMPLE_SEGMENT|8297,8306|false|false|false|||collected
Event|Event|SIMPLE_SEGMENT|8311,8315|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8311,8315|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8311,8315|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8311,8315|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|8330,8331|false|false|false|||_
Event|Event|SIMPLE_SEGMENT|8337,8343|false|false|false|||called
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8349,8352|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8349,8352|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8349,8352|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8349,8352|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8349,8352|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8349,8352|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8349,8352|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8349,8352|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|8349,8352|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8349,8352|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8349,8352|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|8362,8371|false|false|false|||Continued
Drug|Food|SIMPLE_SEGMENT|8385,8389|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|8385,8389|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8385,8389|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|SIMPLE_SEGMENT|8385,8389|false|false|false|||food
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8408,8414|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|8408,8414|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8408,8414|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|8416,8424|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|8430,8436|false|false|false|||eating
Finding|Organism Function|SIMPLE_SEGMENT|8430,8436|false|false|false|C0013470|Eating|eating
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8446,8455|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8446,8455|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|8446,8455|false|false|false|||narcotics
Event|Event|SIMPLE_SEGMENT|8456,8468|false|false|false|||discontinued
Drug|Antibiotic|SIMPLE_SEGMENT|8474,8480|false|false|false|C0700517|Keflex|Keflex
Drug|Organic Chemical|SIMPLE_SEGMENT|8474,8480|false|false|false|C0700517|Keflex|Keflex
Event|Event|SIMPLE_SEGMENT|8474,8480|false|false|false|||Keflex
Event|Event|SIMPLE_SEGMENT|8481,8489|false|false|false|||switched
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8493,8503|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Drug|Substance|SIMPLE_SEGMENT|8493,8503|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Event|Event|SIMPLE_SEGMENT|8493,8503|false|false|false|||suspension
Finding|Functional Concept|SIMPLE_SEGMENT|8493,8503|false|false|false|C1705537|Suspension (action)|suspension
Finding|Body Substance|SIMPLE_SEGMENT|8511,8518|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8511,8518|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8511,8518|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8523,8529|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|8523,8529|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|8530,8534|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|8530,8534|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|8538,8546|false|false|false|||tolerate
Event|Event|SIMPLE_SEGMENT|8556,8559|false|false|false|||set
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8568,8573|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|8568,8573|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|8568,8573|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|8568,8573|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|8568,8573|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8568,8578|false|false|false|C0886052;C1272654|Wound care management;wound care|wound care
Event|Activity|SIMPLE_SEGMENT|8574,8578|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8574,8578|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8574,8578|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8574,8578|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8583,8594|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8583,8594|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8583,8594|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8583,8594|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8583,8607|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8598,8607|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8598,8607|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|8609,8616|false|false|false|C1170371|Lexapro|Lexapro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8609,8616|false|false|false|C1170371|Lexapro|Lexapro
Drug|Organic Chemical|SIMPLE_SEGMENT|8621,8628|false|false|false|C0594492|Nasonex|nasonex
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8621,8628|false|false|false|C0594492|Nasonex|nasonex
Event|Event|SIMPLE_SEGMENT|8621,8628|false|false|false|||nasonex
Event|Event|SIMPLE_SEGMENT|8632,8641|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8632,8641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8632,8641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8632,8641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8632,8641|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8632,8653|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8642,8653|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8642,8653|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8642,8653|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8642,8653|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8658,8670|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8658,8670|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8677,8683|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8697,8703|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8697,8703|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|8728,8739|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8728,8739|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|8728,8739|false|false|false|||Fluticasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8757,8762|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|8757,8762|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|8757,8762|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|8757,8762|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8757,8774|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8764,8774|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|SIMPLE_SEGMENT|8764,8774|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|SIMPLE_SEGMENT|8764,8774|false|false|false|||Suspension
Finding|Functional Concept|SIMPLE_SEGMENT|8764,8774|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8789,8794|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|8789,8794|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|8789,8794|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|8789,8794|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8795,8800|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8795,8800|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|8795,8800|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8795,8800|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|8795,8800|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|8795,8800|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|SIMPLE_SEGMENT|8801,8806|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|8821,8827|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8821,8827|false|false|false|C0282139|Colace|Colace
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8835,8842|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|8835,8842|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8835,8842|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8856,8863|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|8856,8863|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8856,8863|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|SIMPLE_SEGMENT|8875,8878|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8875,8878|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|8883,8889|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|8894,8906|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|8894,8906|false|false|false|C0009806|Constipation|constipation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8930,8937|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|8930,8937|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8930,8937|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|SIMPLE_SEGMENT|8942,8949|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8957,8966|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8957,8966|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8974,8980|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8974,8980|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8994,9000|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8994,9000|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|9028,9034|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9039,9046|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|9039,9046|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9039,9046|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Hormone|SIMPLE_SEGMENT|9053,9067|false|false|false|C0020268|hydrocortisone|Hydrocortisone
Drug|Organic Chemical|SIMPLE_SEGMENT|9053,9067|false|false|false|C0020268|hydrocortisone|Hydrocortisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9053,9067|false|false|false|C0020268|hydrocortisone|Hydrocortisone
Event|Event|SIMPLE_SEGMENT|9053,9067|false|false|false|||Hydrocortisone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9053,9067|false|false|false|C0201968|Cortisol Measurement|Hydrocortisone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9074,9079|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|Cream
Drug|Food|SIMPLE_SEGMENT|9074,9079|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|Cream
Event|Event|SIMPLE_SEGMENT|9080,9083|false|false|false|||Sig
Finding|Gene or Genome|SIMPLE_SEGMENT|9093,9097|false|false|false|C1858559|APPL1 gene|Appl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9098,9104|false|false|false|C1272938|Rectal Dosage Form|Rectal
Finding|Finding|SIMPLE_SEGMENT|9098,9104|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Finding|Functional Concept|SIMPLE_SEGMENT|9098,9104|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Event|Event|SIMPLE_SEGMENT|9105,9108|false|false|false|||TID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9113,9118|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|9121,9124|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9121,9124|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|9129,9135|false|false|false|||needed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9140,9151|false|false|false|C0019112|Hemorrhoids|hemorrhoids
Event|Event|SIMPLE_SEGMENT|9140,9151|false|false|false|||hemorrhoids
Drug|Antibiotic|SIMPLE_SEGMENT|9158,9168|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Organic Chemical|SIMPLE_SEGMENT|9158,9168|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9181,9191|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|SIMPLE_SEGMENT|9181,9191|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|SIMPLE_SEGMENT|9181,9191|false|false|false|||Suspension
Finding|Functional Concept|SIMPLE_SEGMENT|9181,9191|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9181,9210|false|false|false|C2348620|Suspension for Reconstitution Dosage Form|Suspension for Reconstitution
Event|Event|SIMPLE_SEGMENT|9196,9210|false|false|false|||Reconstitution
Finding|Idea or Concept|SIMPLE_SEGMENT|9262,9269|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9277,9284|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9277,9284|false|false|false|C0699142|Tylenol|Tylenol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9292,9298|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9312,9318|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9342,9348|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|9353,9358|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|9353,9358|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9353,9358|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9362,9366|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9362,9366|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9362,9366|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9362,9366|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|9373,9383|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9373,9383|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|SIMPLE_SEGMENT|9384,9387|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|SIMPLE_SEGMENT|9384,9387|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|SIMPLE_SEGMENT|9388,9392|false|false|false|||Work
Event|Occupational Activity|SIMPLE_SEGMENT|9388,9392|false|false|false|C0043227|Work|Work
Event|Event|SIMPLE_SEGMENT|9400,9405|false|false|false|||check
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9406,9411|false|false|false|C5575602|Cell Culture Serum|serum
Finding|Body Substance|SIMPLE_SEGMENT|9406,9411|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|SIMPLE_SEGMENT|9406,9411|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Finding|SIMPLE_SEGMENT|9406,9422|false|false|false|C0600061|Serum creatinine level|serum Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9406,9422|false|false|false|C0201976|Creatinine measurement, serum (procedure)|serum Creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9412,9422|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|9412,9422|false|false|false|C0010294|creatinine|Creatinine
Event|Event|SIMPLE_SEGMENT|9412,9422|false|false|false|||Creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|9412,9422|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9412,9422|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|SIMPLE_SEGMENT|9439,9445|false|false|false|||result
Finding|Finding|SIMPLE_SEGMENT|9439,9445|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|9439,9445|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|9439,9445|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9449,9452|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9449,9452|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9449,9452|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9449,9452|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|9449,9452|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9449,9452|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|9449,9452|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9449,9452|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|9449,9452|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|9449,9452|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|9449,9452|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9472,9483|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|9472,9483|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|9472,9483|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|9485,9489|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9485,9489|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9485,9489|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9485,9489|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|9495,9502|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|9495,9502|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|9505,9513|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9505,9513|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|9521,9530|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9521,9530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9521,9530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9521,9530|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9521,9530|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9521,9540|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9531,9540|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9531,9540|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9531,9540|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9531,9540|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9531,9540|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9561,9575|false|false|false|C0012813|Diverticulitis|Diverticulitis
Event|Event|SIMPLE_SEGMENT|9561,9575|false|false|false|||Diverticulitis
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9584,9589|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|9584,9589|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|9584,9589|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|9584,9589|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|9584,9589|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9584,9600|false|false|false|C0406832|Wound cellulitis|wound cellulitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9590,9600|false|false|false|C0007642|Cellulitis|cellulitis
Event|Event|SIMPLE_SEGMENT|9590,9600|false|false|false|||cellulitis
Finding|Finding|SIMPLE_SEGMENT|9590,9600|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Event|Event|SIMPLE_SEGMENT|9609,9620|false|false|false|||hypovolemia
Finding|Finding|SIMPLE_SEGMENT|9609,9620|false|false|false|C0546884|Hypovolemia|hypovolemia
Event|Event|SIMPLE_SEGMENT|9629,9634|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|9629,9634|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9629,9634|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9637,9646|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|9637,9646|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|9637,9646|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9648,9655|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|SIMPLE_SEGMENT|9648,9655|false|false|false|||Anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9648,9655|false|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9656,9670|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|SIMPLE_SEGMENT|9656,9670|false|false|false|||diverticulosis
Event|Event|SIMPLE_SEGMENT|9674,9683|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9674,9683|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9674,9683|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9674,9683|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9674,9683|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9684,9693|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9684,9693|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9684,9693|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9684,9693|false|false|false|C1705253|Logical Condition|Condition
Event|Event|SIMPLE_SEGMENT|9695,9701|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|9695,9701|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Finding|SIMPLE_SEGMENT|9724,9727|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|9724,9727|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Conceptual Entity|SIMPLE_SEGMENT|9728,9735|false|false|false|C1709915|Residue|residue
Drug|Food|SIMPLE_SEGMENT|9736,9740|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|9736,9740|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|9736,9740|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|9736,9740|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9750,9754|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9750,9754|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9750,9754|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9750,9754|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9750,9762|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9750,9762|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|SIMPLE_SEGMENT|9755,9762|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9755,9762|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|9755,9762|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|9755,9762|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|9755,9762|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|9755,9762|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|9755,9762|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9768,9772|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9768,9772|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9768,9772|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9768,9772|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9768,9783|false|false|false|C5848556|Oral medication (substance)|oral medication
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9768,9783|false|false|false|C0175795|Oral Medication|oral medication
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9773,9783|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9773,9783|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9773,9783|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9787,9796|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9787,9796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9787,9796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9787,9796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9787,9796|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9787,9809|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9787,9809|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9787,9809|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9797,9809|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9797,9809|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9797,9809|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|9818,9822|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|9828,9834|true|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|9828,9834|true|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|9838,9844|true|false|false|||return
Event|Event|SIMPLE_SEGMENT|9888,9898|false|false|false|||experience
Finding|Finding|SIMPLE_SEGMENT|9899,9902|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|9899,9902|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9903,9908|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9903,9908|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9903,9913|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9903,9913|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9909,9913|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9909,9913|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9909,9913|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9909,9913|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9915,9923|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|9915,9923|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|9915,9923|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9915,9923|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9915,9923|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|9925,9934|false|false|false|||squeezing
Event|Event|SIMPLE_SEGMENT|9939,9948|false|false|false|||tightness
Finding|Finding|SIMPLE_SEGMENT|9952,9955|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|9952,9955|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|9959,9968|false|true|false|C1546960|Patient Outcome - Worsening|worsening
Drug|Organic Chemical|SIMPLE_SEGMENT|9969,9974|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9969,9974|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|9969,9974|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|9969,9974|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|9978,9986|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|9978,9986|false|true|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|10001,10009|true|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|10001,10009|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|10021,10025|true|false|false|||keep
Drug|Substance|SIMPLE_SEGMENT|10030,10036|true|false|true|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|10030,10036|true|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|10030,10036|true|false|true|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10030,10036|true|false|true|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10046,10057|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10046,10057|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10046,10057|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10046,10057|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10077,10087|false|false|false|C0011175|Dehydration|dehydrated
Event|Event|SIMPLE_SEGMENT|10077,10087|false|false|false|||dehydrated
Event|Event|SIMPLE_SEGMENT|10095,10104|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|10105,10113|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|10105,10113|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|10116,10124|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|10116,10124|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10116,10124|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|10134,10141|false|false|false|||reasons
Finding|Idea or Concept|SIMPLE_SEGMENT|10134,10141|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Event|Event|SIMPLE_SEGMENT|10143,10148|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|10143,10148|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|10143,10148|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Finding|SIMPLE_SEGMENT|10143,10163|false|false|false|C5924540|Signs of dehydration|Signs of dehydration
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10152,10163|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10152,10163|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|SIMPLE_SEGMENT|10152,10163|false|false|false|||dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10152,10163|false|false|false|C4284399|Dehydration procedure|dehydration
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10177,10182|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10177,10182|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|SIMPLE_SEGMENT|10184,10199|false|false|false|C0039231|Tachycardia|rapid heartbeat
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10190,10199|false|false|false|C0232117|Pulse Rate|heartbeat
Event|Event|SIMPLE_SEGMENT|10190,10199|false|false|false|||heartbeat
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10190,10199|false|false|false|C0425583|Heart beat|heartbeat
Event|Event|SIMPLE_SEGMENT|10203,10210|false|false|false|||feeling
Finding|Mental Process|SIMPLE_SEGMENT|10203,10210|false|false|false|C1527305|Feelings|feeling
Finding|Sign or Symptom|SIMPLE_SEGMENT|10203,10216|false|false|false|C0849959|feeling dizzy|feeling dizzy
Finding|Sign or Symptom|SIMPLE_SEGMENT|10211,10216|false|false|false|C0012833|Dizziness|dizzy
Event|Event|SIMPLE_SEGMENT|10220,10225|false|false|false|||faint
Finding|Finding|SIMPLE_SEGMENT|10220,10225|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|SIMPLE_SEGMENT|10220,10225|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Event|Event|SIMPLE_SEGMENT|10247,10250|false|false|false|||see
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10251,10256|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10251,10256|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10251,10256|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Substance|SIMPLE_SEGMENT|10271,10279|false|false|false|C0520510|Materials|material
Event|Event|SIMPLE_SEGMENT|10271,10279|false|false|false|||material
Event|Event|SIMPLE_SEGMENT|10289,10294|false|false|false|||vomit
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10306,10311|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|10306,10320|false|false|false|C0011135|Defecation|bowel movement
Event|Event|SIMPLE_SEGMENT|10312,10320|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|10312,10320|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10329,10333|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10329,10333|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10329,10333|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10329,10333|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10341,10350|true|false|false|||improving
Event|Event|SIMPLE_SEGMENT|10375,10379|true|false|false|||gone
Event|Event|SIMPLE_SEGMENT|10398,10402|false|false|false|||Call
Finding|Functional Concept|SIMPLE_SEGMENT|10398,10402|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|SIMPLE_SEGMENT|10398,10402|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|SIMPLE_SEGMENT|10398,10402|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|SIMPLE_SEGMENT|10398,10402|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Event|Event|SIMPLE_SEGMENT|10406,10412|false|false|false|||return
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10433,10437|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10433,10437|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10433,10437|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10433,10437|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10450,10455|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|10450,10455|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|10450,10455|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Functional Concept|SIMPLE_SEGMENT|10462,10470|false|false|false|C0392747|Changing|changing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10471,10479|false|false|false|C1515974|Anatomic Site|location
Event|Event|SIMPLE_SEGMENT|10471,10479|false|false|false|||location
Finding|Intellectual Product|SIMPLE_SEGMENT|10471,10479|false|false|false|C1555588|Transaction counts and value totals - location|location
Event|Event|SIMPLE_SEGMENT|10483,10489|false|false|false|||moving
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10498,10503|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|10498,10503|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|10509,10513|false|false|false|||back
Event|Event|SIMPLE_SEGMENT|10522,10529|false|false|false|||driving
Event|Event|SIMPLE_SEGMENT|10533,10542|false|false|false|||operating
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10549,10558|false|false|false|C0337246|Contact with machinery|machinery
Event|Event|SIMPLE_SEGMENT|10549,10558|false|false|false|||machinery
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10572,10576|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10572,10576|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10572,10576|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10572,10576|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10578,10589|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10578,10589|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10578,10589|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10578,10589|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|10610,10616|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|10610,10616|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|10623,10628|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|10623,10628|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|10623,10628|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|10653,10660|false|false|false|||degrees
Finding|Intellectual Product|SIMPLE_SEGMENT|10653,10660|false|false|false|C0542560|Academic degree|degrees
Event|Event|SIMPLE_SEGMENT|10670,10677|false|false|false|||degrees
Finding|Intellectual Product|SIMPLE_SEGMENT|10670,10677|false|false|false|C0542560|Academic degree|degrees
Finding|Finding|SIMPLE_SEGMENT|10685,10692|true|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Finding|Idea or Concept|SIMPLE_SEGMENT|10685,10692|true|false|false|C1551395;C1552745;C1561576|Alert level - Serious;Device Alert Level - Serious;Equipment Alert Level - Serious|serious
Event|Event|SIMPLE_SEGMENT|10693,10699|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|10693,10699|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10693,10699|true|false|false|C4319952|Change - procedure|change
Event|Event|SIMPLE_SEGMENT|10709,10717|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|10709,10717|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10709,10717|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|SIMPLE_SEGMENT|10726,10729|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|10726,10729|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|10730,10738|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|10730,10738|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10730,10738|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|10745,10752|true|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|10745,10752|true|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|10768,10774|true|false|false|||resume
Finding|Idea or Concept|SIMPLE_SEGMENT|10787,10791|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10787,10791|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10787,10791|true|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10792,10803|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10792,10803|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10792,10803|true|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10792,10803|true|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|10808,10812|true|false|false|||take
Event|Event|SIMPLE_SEGMENT|10817,10820|true|false|false|||new
Finding|Finding|SIMPLE_SEGMENT|10817,10820|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|10817,10820|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10822,10826|true|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|SIMPLE_SEGMENT|10822,10826|true|false|false|||meds
Finding|Intellectual Product|SIMPLE_SEGMENT|10822,10826|true|false|false|C4284232|Medications|meds
Event|Event|SIMPLE_SEGMENT|10831,10838|true|false|false|||ordered
Event|Event|SIMPLE_SEGMENT|10843,10851|false|false|false|||Continue
Event|Event|SIMPLE_SEGMENT|10855,10863|false|false|false|||ambulate
Finding|Finding|SIMPLE_SEGMENT|10864,10885|false|false|false|C4489371|Several times per day|several times per day
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10872,10877|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|10882,10885|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10882,10885|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10889,10894|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|SIMPLE_SEGMENT|10889,10894|false|false|false|||WOUND
Finding|Body Substance|SIMPLE_SEGMENT|10889,10894|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|SIMPLE_SEGMENT|10889,10894|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|SIMPLE_SEGMENT|10889,10894|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10889,10899|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|SIMPLE_SEGMENT|10895,10899|false|false|false|C1947933|care activity|CARE
Event|Event|SIMPLE_SEGMENT|10895,10899|false|false|false|||CARE
Finding|Finding|SIMPLE_SEGMENT|10895,10899|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|10895,10899|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Procedure|Health Care Activity|SIMPLE_SEGMENT|10909,10917|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10909,10917|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10909,10923|false|false|false|C0332803|Surgical wound|surgical wound
Finding|Finding|SIMPLE_SEGMENT|10909,10923|false|false|false|C1628502|Surgical wound finding|surgical wound
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10918,10923|false|true|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|10918,10923|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|10918,10923|false|true|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|10918,10923|false|true|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|10918,10923|false|true|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10924,10928|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|10924,10928|false|false|false|C1546778||site
Finding|Functional Concept|SIMPLE_SEGMENT|10937,10943|false|false|false|C0392747|Changing|Change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10937,10943|false|false|false|C4319952|Change - procedure|Change
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10944,10951|false|false|false|C1706363|Packing Dosage Form|packing
Event|Activity|SIMPLE_SEGMENT|10944,10951|false|false|false|C2828395|Packing (action)|packing
Event|Event|SIMPLE_SEGMENT|10944,10951|false|false|false|||packing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10944,10951|false|false|false|C0184967|Insertion of pack (procedure)|packing
Finding|Intellectual Product|SIMPLE_SEGMENT|10961,10965|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|SIMPLE_SEGMENT|10970,10973|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10970,10973|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|10982,10988|false|false|false|||needed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10991,10995|false|false|false|C1999262|Pack|Pack
Event|Activity|SIMPLE_SEGMENT|10991,10995|false|false|false|C2828395|Packing (action)|Pack
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11025,11031|false|false|false|C0036082|Saline Solution|Saline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11025,11031|false|false|false|C0036082|Saline Solution|Saline
Event|Event|SIMPLE_SEGMENT|11025,11031|false|false|false|||Saline
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11025,11031|false|false|false|C0450082|Saline method|Saline
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11038,11048|false|false|false|C0184898|Surgical incisions|incisional
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11050,11056|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|11050,11056|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11050,11056|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|11050,11056|false|false|false|||cavity
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11086,11092|false|false|false|C3714578|Fix|adhere
Finding|Idea or Concept|SIMPLE_SEGMENT|11098,11103|false|false|false|C1547566|Paper Authorization|paper
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11104,11108|false|false|false|C1704747|Tape Dosage Form|tape
Event|Event|SIMPLE_SEGMENT|11104,11108|false|false|false|||tape
Finding|Gene or Genome|SIMPLE_SEGMENT|11104,11108|false|false|false|C1824539|CC2D1A gene|tape
Finding|Functional Concept|SIMPLE_SEGMENT|11112,11119|false|false|false|C0392747|Changing|Changed
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11139,11148|false|false|false|C0522534|Saturated|saturated
Event|Event|SIMPLE_SEGMENT|11152,11159|false|false|false|||prevent
Event|Event|SIMPLE_SEGMENT|11160,11170|false|false|false|||irritation
Finding|Intellectual Product|SIMPLE_SEGMENT|11160,11170|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|SIMPLE_SEGMENT|11160,11170|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|SIMPLE_SEGMENT|11160,11170|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11160,11170|false|false|false|C0441723|Irritation|irritation
Anatomy|Body System|SIMPLE_SEGMENT|11187,11191|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11187,11191|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11187,11191|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|11187,11191|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|11187,11191|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|11187,11191|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11198,11203|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|11198,11203|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|11198,11203|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|11198,11203|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|11198,11203|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|SIMPLE_SEGMENT|11204,11213|false|false|false|||continues
Event|Event|SIMPLE_SEGMENT|11217,11221|false|false|false|||weep
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11223,11227|false|false|false|C1999262|Pack|pack
Event|Activity|SIMPLE_SEGMENT|11223,11227|false|false|false|C2828395|Packing (action)|pack
Event|Event|SIMPLE_SEGMENT|11223,11227|false|false|false|||pack
Drug|Organic Chemical|SIMPLE_SEGMENT|11234,11241|false|false|false|C0967370|Aquacel|Aquacel
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|11245,11248|false|false|false|C0036875;C1842691|Diaphanospondylodysostosis;Disorders of Sex Development|DSD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11245,11248|false|false|false|C0036875;C1842691|Diaphanospondylodysostosis;Disorders of Sex Development|DSD
Event|Event|SIMPLE_SEGMENT|11245,11248|false|false|false|||DSD
Event|Event|SIMPLE_SEGMENT|11259,11265|false|false|false|||shower
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11279,11283|false|false|false|C1883550|Wash Dosage Form|wash
Event|Activity|SIMPLE_SEGMENT|11279,11283|false|false|false|C0441648|Wash (cleansing action)|wash
Event|Event|SIMPLE_SEGMENT|11279,11283|false|false|false|||wash
Finding|Functional Concept|SIMPLE_SEGMENT|11279,11283|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Finding|Gene or Genome|SIMPLE_SEGMENT|11279,11283|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Finding|Intellectual Product|SIMPLE_SEGMENT|11279,11283|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11279,11283|false|false|false|C2699154|Cell Wash|wash
Procedure|Health Care Activity|SIMPLE_SEGMENT|11291,11299|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11291,11299|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11291,11309|false|false|false|C0332803|Surgical wound|surgical incisions
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11291,11309|false|false|false|C0184898|Surgical incisions|surgical incisions
Event|Event|SIMPLE_SEGMENT|11300,11309|false|false|false|||incisions
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11300,11309|false|false|false|C0184898|Surgical incisions|incisions
Event|Event|SIMPLE_SEGMENT|11318,11326|false|false|false|||swimming
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11318,11326|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|SIMPLE_SEGMENT|11318,11326|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Gene or Genome|SIMPLE_SEGMENT|11331,11334|false|false|false|C1421225|TUB gene|tub
Event|Event|SIMPLE_SEGMENT|11335,11340|false|false|false|||baths
Procedure|Health Care Activity|SIMPLE_SEGMENT|11335,11340|false|false|false|C0150141|Bathing|baths
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11347,11352|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|11347,11352|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|11347,11352|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|11347,11352|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|11347,11352|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|11353,11363|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|11364,11370|false|false|false|||healed
Event|Event|SIMPLE_SEGMENT|11379,11383|false|false|false|||call
Event|Event|SIMPLE_SEGMENT|11388,11394|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|11388,11394|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11417,11421|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11417,11421|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11417,11421|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11417,11421|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|11423,11431|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|11423,11431|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|11423,11431|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11434,11441|false|false|false|C0041834|Erythema|redness
Event|Event|SIMPLE_SEGMENT|11434,11441|false|false|false|||redness
Finding|Finding|SIMPLE_SEGMENT|11434,11441|false|false|false|C0332575|Redness|redness
Event|Event|SIMPLE_SEGMENT|11446,11454|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|11446,11454|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|11446,11454|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11446,11454|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11464,11472|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11464,11472|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11464,11472|false|false|false|C0184898|Surgical incisions|incision
Event|Event|SIMPLE_SEGMENT|11473,11478|false|false|false|||sites
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11482,11492|false|false|false|C0010294|creatinine|CREATININE
Drug|Organic Chemical|SIMPLE_SEGMENT|11482,11492|false|false|false|C0010294|creatinine|CREATININE
Event|Event|SIMPLE_SEGMENT|11482,11492|false|false|false|||CREATININE
Finding|Physiologic Function|SIMPLE_SEGMENT|11482,11492|false|false|false|C4551889|Creatinine metabolic function|CREATININE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11482,11492|false|false|false|C0201975|Creatinine measurement|CREATININE
Event|Event|SIMPLE_SEGMENT|11515,11520|false|false|false|||check
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11526,11536|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|11526,11536|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|11526,11536|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|11526,11536|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11526,11536|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|11553,11557|false|false|false|||call
Finding|Functional Concept|SIMPLE_SEGMENT|11553,11557|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|11553,11557|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|11553,11557|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|11553,11557|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11578,11581|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11578,11581|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11578,11581|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11578,11581|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|11578,11581|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11578,11581|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|11578,11581|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11578,11581|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|11578,11581|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|11578,11581|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|11578,11581|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|11584,11590|false|false|false|||office
Finding|Idea or Concept|SIMPLE_SEGMENT|11584,11590|false|false|false|C1549636|Address type - Office|office
Event|Event|SIMPLE_SEGMENT|11601,11607|false|false|false|||result
Finding|Finding|SIMPLE_SEGMENT|11601,11607|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|11601,11607|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|11601,11607|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Procedure|Health Care Activity|SIMPLE_SEGMENT|11612,11620|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11621,11633|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11621,11633|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11621,11633|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

