 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|44,53|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|44,53|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|44,58|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|78,87|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|78,87|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|78,92|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|134,137|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|145,152|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|145,152|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|154,166|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|154,166|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|169,178|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|169,178|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|169,178|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Body Substance|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|189,197|true|false|false|||recorded
Attribute|Clinical Attribute|SIMPLE_SEGMENT|217,226|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|217,226|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|217,226|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|230,235|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|SIMPLE_SEGMENT|230,235|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|230,235|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|SIMPLE_SEGMENT|238,247|true|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|238,247|true|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|256,271|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|262,271|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|262,271|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|262,271|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Finding|SIMPLE_SEGMENT|273,277|false|false|false|C0016928|Gait|Gait
Finding|Finding|SIMPLE_SEGMENT|273,289|false|false|false|C0231686|Gait, Unsteady|Gait instability
Event|Event|SIMPLE_SEGMENT|278,289|false|false|false|||instability
Finding|Finding|SIMPLE_SEGMENT|278,289|false|false|false|C1444783|Instability|instability
Finding|Finding|SIMPLE_SEGMENT|291,305|false|false|false|C0743800|multiple falls|multiple falls
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|300,305|false|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|300,305|false|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|300,305|false|false|false|C0085639|Falls|falls
Finding|Classification|SIMPLE_SEGMENT|308,313|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|314,322|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|314,322|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|326,344|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|335,344|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|335,344|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|335,344|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|335,344|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|335,344|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|354,361|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|354,361|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,361|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|354,361|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|354,364|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|354,380|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|354,380|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|365,372|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|365,372|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|365,380|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|373,380|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|394,402|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|394,402|false|false|false|C2987187|Pleasant|pleasant
Finding|Functional Concept|SIMPLE_SEGMENT|403,408|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|403,415|false|false|false|C0230370|Structure of right hand|right handed
Finding|Idea or Concept|SIMPLE_SEGMENT|420,424|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|420,424|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|429,433|false|false|false|||male
Finding|Finding|SIMPLE_SEGMENT|429,433|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|439,443|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|439,443|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Drug|Organic Chemical|SIMPLE_SEGMENT|449,457|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|449,457|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|449,457|false|false|false|||coumadin
Event|Event|SIMPLE_SEGMENT|472,483|false|false|false|||independent
Finding|Finding|SIMPLE_SEGMENT|472,483|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|independent
Finding|Idea or Concept|SIMPLE_SEGMENT|472,483|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|independent
Event|Event|SIMPLE_SEGMENT|485,491|false|false|false|||living
Finding|Idea or Concept|SIMPLE_SEGMENT|520,524|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|525,530|false|false|false|||state
Finding|Functional Concept|SIMPLE_SEGMENT|525,530|false|false|false|C1442792|State|state
Finding|Finding|SIMPLE_SEGMENT|525,540|false|false|false|C0683314|personal health|state of health
Event|Event|SIMPLE_SEGMENT|534,540|false|false|false|||health
Finding|Idea or Concept|SIMPLE_SEGMENT|534,540|false|false|false|C0018684|Health|health
Finding|Idea or Concept|SIMPLE_SEGMENT|556,560|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|556,560|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|SIMPLE_SEGMENT|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|585,592|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|601,606|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|614,621|false|false|false|||periods
Finding|Organism Function|SIMPLE_SEGMENT|614,621|false|false|false|C0025344|Menstruation|periods
Event|Event|SIMPLE_SEGMENT|625,637|false|false|false|||disorganized
Event|Event|SIMPLE_SEGMENT|639,645|false|false|false|||speech
Finding|Organism Function|SIMPLE_SEGMENT|639,645|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|639,645|false|false|false|C0846595|Speech assessment|speech
Finding|Finding|SIMPLE_SEGMENT|650,654|false|false|false|C0016928|Gait|gait
Finding|Finding|SIMPLE_SEGMENT|650,666|false|false|false|C0231686|Gait, Unsteady|gait instability
Event|Event|SIMPLE_SEGMENT|655,666|false|false|false|||instability
Finding|Finding|SIMPLE_SEGMENT|655,666|false|false|false|C1444783|Instability|instability
Finding|Finding|SIMPLE_SEGMENT|684,690|true|false|false|C1561668|History of fall|a fall
Event|Event|SIMPLE_SEGMENT|686,690|true|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|686,690|true|true|false|C0085639|Falls|fall
Finding|Gene or Genome|SIMPLE_SEGMENT|707,710|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|719,724|false|false|false|||broke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|733,737|false|false|false|C0035561|Bone structure of rib|ribs
Drug|Food|SIMPLE_SEGMENT|745,751|false|false|false|C0009237|Coffee|coffee
Event|Event|SIMPLE_SEGMENT|752,757|false|false|false|||table
Finding|Intellectual Product|SIMPLE_SEGMENT|752,757|false|false|false|C1706074|Data Table|table
Anatomy|Body Location or Region|SIMPLE_SEGMENT|780,784|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|780,784|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|780,784|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|780,784|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|780,791|true|false|false|C0018674|Craniocerebral Trauma|head trauma
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|785,791|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|785,791|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|785,791|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|804,811|true|false|false|||scanned
Event|Event|SIMPLE_SEGMENT|818,821|true|false|false|||OSH
Event|Event|SIMPLE_SEGMENT|836,842|false|false|false|||speech
Finding|Organism Function|SIMPLE_SEGMENT|836,842|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|836,842|false|false|false|C0846595|Speech assessment|speech
Event|Event|SIMPLE_SEGMENT|847,859|false|false|false|||unsteadiness
Finding|Finding|SIMPLE_SEGMENT|847,859|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|SIMPLE_SEGMENT|865,870|false|false|false|||waxed
Event|Event|SIMPLE_SEGMENT|875,880|false|false|false|||waned
Event|Event|SIMPLE_SEGMENT|918,925|false|false|false|||reports
Finding|Finding|SIMPLE_SEGMENT|940,944|false|false|false|C4281574|Much|much
Event|Event|SIMPLE_SEGMENT|945,953|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|963,968|false|false|false|||takes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|973,982|false|false|false|C0012798|Diuretics|diuretics
Event|Event|SIMPLE_SEGMENT|973,982|false|false|false|||diuretics
Event|Event|SIMPLE_SEGMENT|994,1000|false|false|false|||period
Finding|Organism Function|SIMPLE_SEGMENT|994,1000|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|SIMPLE_SEGMENT|994,1000|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|SIMPLE_SEGMENT|1008,1012|false|false|false|||lost
Event|Event|SIMPLE_SEGMENT|1018,1021|false|false|false|||lbs
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1018,1021|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|SIMPLE_SEGMENT|1042,1049|false|false|false|||sorting
Event|Event|SIMPLE_SEGMENT|1050,1056|false|false|false|||papers
Finding|Intellectual Product|SIMPLE_SEGMENT|1076,1081|false|false|false|C1706074|Data Table|table
Event|Event|SIMPLE_SEGMENT|1091,1095|false|false|false|||fell
Event|Event|SIMPLE_SEGMENT|1101,1109|false|false|false|||standing
Event|Event|SIMPLE_SEGMENT|1125,1134|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1125,1134|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|1139,1146|true|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1151,1154|true|false|false|||LOC
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1159,1163|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1159,1163|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1159,1163|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1159,1163|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1159,1170|true|false|false|C0018674|Craniocerebral Trauma|head trauma
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1164,1170|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|1164,1170|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|1164,1170|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|1179,1183|true|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1179,1183|true|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|1187,1192|true|false|false|||stand
Event|Event|SIMPLE_SEGMENT|1198,1200|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|1205,1213|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|1205,1213|false|false|false|C0549178|Continuous|continue
Event|Event|SIMPLE_SEGMENT|1219,1223|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|1219,1223|false|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|1234,1240|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|1266,1269|false|false|false|||got
Event|Event|SIMPLE_SEGMENT|1283,1287|false|false|false|||fell
Event|Event|SIMPLE_SEGMENT|1315,1321|true|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1326,1329|true|false|false|||LOC
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1333,1337|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1333,1337|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1333,1337|true|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|1333,1337|true|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1333,1337|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1339,1345|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|1339,1345|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|1339,1345|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|1347,1354|true|false|false|||blaming
Event|Event|SIMPLE_SEGMENT|1359,1370|false|false|false|||instability
Finding|Finding|SIMPLE_SEGMENT|1359,1370|false|false|false|C1444783|Instability|instability
Event|Event|SIMPLE_SEGMENT|1379,1387|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1379,1387|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1400,1406|true|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1400,1406|true|false|false|C0153933|Benign neoplasm of tongue|tongue
Event|Event|SIMPLE_SEGMENT|1400,1406|true|false|false|||tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|1400,1406|true|false|false|C0872394|Procedure on tongue|tongue
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1400,1413|true|false|false|C0241424|Tongue biting|tongue biting
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1407,1413|true|false|false|C0005658|bite injury|biting
Event|Event|SIMPLE_SEGMENT|1407,1413|true|false|false|||biting
Finding|Physiologic Function|SIMPLE_SEGMENT|1407,1413|true|false|false|C2584293|Biting|biting
Event|Event|SIMPLE_SEGMENT|1417,1421|true|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1417,1421|true|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1425,1430|true|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1431,1438|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1431,1438|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1431,1438|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Finding|SIMPLE_SEGMENT|1431,1449|false|false|false|C0876938;C4319531|Bladder Continence Question;Urinary bladder control|bladder continence
Finding|Intellectual Product|SIMPLE_SEGMENT|1431,1449|false|false|false|C0876938;C4319531|Bladder Continence Question;Urinary bladder control|bladder continence
Event|Event|SIMPLE_SEGMENT|1439,1449|false|false|false|||continence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1463,1466|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|1463,1466|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|1463,1466|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|1498,1510|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|1498,1510|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|1525,1534|false|false|false|||concerned
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1545,1550|false|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|1545,1550|false|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|1545,1550|false|false|false|C0085639|Falls|falls
Event|Event|SIMPLE_SEGMENT|1555,1562|false|false|false|||brought
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1594,1603|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|1594,1603|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|1594,1603|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|1594,1603|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1594,1603|false|false|false|C0011900|Diagnosis|diagnosis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1607,1612|false|false|false|C0378717|elongation factor DmS-II|DM II
Finding|Idea or Concept|SIMPLE_SEGMENT|1630,1635|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|1630,1635|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|SIMPLE_SEGMENT|1636,1639|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|1649,1656|false|false|false|||started
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1657,1661|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1657,1661|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|1657,1661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|1657,1661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1657,1675|false|false|false|C0359086|Oral hypoglycemic|oral hypoglycemics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1662,1675|false|false|false|C0020616|Hypoglycemic Agents|hypoglycemics
Event|Event|SIMPLE_SEGMENT|1662,1675|false|false|false|||hypoglycemics
Event|Event|SIMPLE_SEGMENT|1689,1696|false|false|false|||reports
Finding|Finding|SIMPLE_SEGMENT|1704,1707|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|1704,1707|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|1716,1720|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|1716,1720|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1716,1720|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1716,1720|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|1729,1733|false|false|false|||seen
Finding|Intellectual Product|SIMPLE_SEGMENT|1764,1768|false|false|false|C1561540|Transaction counts and value totals - week|week
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1794,1801|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1794,1801|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1797,1801|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1797,1801|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1797,1801|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|1797,1801|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1797,1801|false|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|1808,1817|false|false|false|||completed
Finding|Intellectual Product|SIMPLE_SEGMENT|1832,1836|false|false|false|C1561540|Transaction counts and value totals - week|week
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1853,1857|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1853,1857|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1853,1857|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|1853,1857|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1853,1857|false|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|1862,1869|false|false|false|||scanned
Event|Event|SIMPLE_SEGMENT|1876,1884|true|false|false|||revealed
Event|Event|SIMPLE_SEGMENT|1888,1893|true|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|1888,1893|true|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1907,1919|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1907,1919|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1915,1919|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|1915,1919|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|1932,1936|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Cell Component|SIMPLE_SEGMENT|1968,1975|true|false|false|C1660780|midline cell component|midline
Finding|Finding|SIMPLE_SEGMENT|1968,1981|true|false|false|C4086580|Midline Shift|midline shift
Event|Event|SIMPLE_SEGMENT|1976,1981|true|false|false|||shift
Finding|Functional Concept|SIMPLE_SEGMENT|1976,1981|true|false|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1976,1981|true|false|false|C2347509|Physical Shift|shift
Event|Event|SIMPLE_SEGMENT|1983,1995|false|false|false|||Neurosurgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1983,1995|false|false|false|C0524850|Neurosurgical Procedures|Neurosurgery
Event|Event|SIMPLE_SEGMENT|2000,2009|false|false|false|||contacted
Event|Event|SIMPLE_SEGMENT|2014,2024|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|2014,2024|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2014,2024|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|2033,2037|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|2046,2054|false|false|false|C0332149|Possible|possible
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2055,2059|false|false|false|C5890809||role
Event|Event|SIMPLE_SEGMENT|2055,2059|false|false|false|||role
Finding|Conceptual Entity|SIMPLE_SEGMENT|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Intellectual Product|SIMPLE_SEGMENT|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Social Behavior|SIMPLE_SEGMENT|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Body Substance|SIMPLE_SEGMENT|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2084,2092|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|2084,2092|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|2084,2092|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|SIMPLE_SEGMENT|2098,2118|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2103,2110|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2103,2110|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2103,2110|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2103,2110|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2103,2110|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2103,2118|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2111,2118|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2111,2118|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2111,2118|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2120,2125|false|false|false|C0378717|elongation factor DmS-II|DM II
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2127,2130|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2127,2130|false|false|false|||HTN
Drug|Organic Chemical|SIMPLE_SEGMENT|2156,2164|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2156,2164|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|2156,2164|false|false|false|||coumadin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2166,2174|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2166,2174|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2166,2174|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2166,2177|false|false|false|C0376358|Malignant neoplasm of prostate|prostate CA
Event|Event|SIMPLE_SEGMENT|2175,2177|false|false|false|||CA
Event|Event|SIMPLE_SEGMENT|2179,2186|false|false|false|||treated
Finding|Functional Concept|SIMPLE_SEGMENT|2206,2212|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2206,2220|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2213,2220|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2213,2220|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2213,2220|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2213,2220|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2226,2232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2226,2232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2226,2232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2226,2232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2226,2240|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2233,2240|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2233,2240|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2233,2240|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2233,2240|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2262,2270|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2262,2270|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2262,2270|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2262,2270|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2262,2275|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2262,2275|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2271,2275|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2271,2275|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2271,2275|false|false|false|C0582103|Medical Examination|Exam
Finding|Finding|SIMPLE_SEGMENT|2277,2289|false|false|false|C4533677|at admission|At Admission
Event|Event|SIMPLE_SEGMENT|2280,2289|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2280,2289|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|2293,2296|false|false|false|||Gen
Finding|Classification|SIMPLE_SEGMENT|2293,2296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|2293,2296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|2305,2316|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|2305,2316|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2318,2321|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2318,2321|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2318,2321|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2318,2321|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2323,2328|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2330,2336|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|2346,2350|false|false|false|||EOMs
Finding|Functional Concept|SIMPLE_SEGMENT|2346,2350|false|false|false|C0241886|Extraocular|EOMs
Event|Event|SIMPLE_SEGMENT|2351,2357|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2351,2357|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2362,2367|false|false|false|C0024109|Lung|Lungs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2369,2372|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|2369,2372|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2369,2372|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2369,2372|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2386,2393|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2386,2393|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|SIMPLE_SEGMENT|2416,2435|false|false|false|C0232258|Pansystolic murmur|holosystolic murmur
Event|Event|SIMPLE_SEGMENT|2429,2435|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|2429,2435|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2437,2440|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2437,2440|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2442,2446|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2442,2446|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2448,2450|false|false|false|||NT
Event|Event|SIMPLE_SEGMENT|2464,2468|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|2464,2468|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2464,2468|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|2473,2477|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2478,2486|false|false|false|||perfused
Finding|Mental Process|SIMPLE_SEGMENT|2495,2501|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2495,2508|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|SIMPLE_SEGMENT|2495,2508|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2502,2508|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|2502,2508|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|2502,2508|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|2510,2515|false|false|false|||Awake
Finding|Finding|SIMPLE_SEGMENT|2510,2515|false|false|false|C0234422|Awake (finding)|Awake
Event|Event|SIMPLE_SEGMENT|2520,2531|false|false|false|||cooperative
Event|Event|SIMPLE_SEGMENT|2537,2541|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2537,2541|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2537,2541|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|2550,2556|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|2550,2556|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|2550,2556|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|2558,2569|false|false|false|||Orientation
Finding|Mental Process|SIMPLE_SEGMENT|2558,2569|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|SIMPLE_SEGMENT|2571,2579|false|false|false|||Oriented
Finding|Finding|SIMPLE_SEGMENT|2571,2579|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|SIMPLE_SEGMENT|2571,2589|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2583,2589|false|false|false|C5890614||person
Event|Event|SIMPLE_SEGMENT|2583,2589|false|false|false|||person
Finding|Intellectual Product|SIMPLE_SEGMENT|2583,2589|false|false|false|C1522390|Person Info|person
Event|Activity|SIMPLE_SEGMENT|2591,2596|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|2591,2596|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|2591,2596|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|2591,2596|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|2608,2614|false|false|false|||Recall
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|2608,2614|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|SIMPLE_SEGMENT|2608,2614|false|false|false|C0034770|Mental Recall|Recall
Event|Event|SIMPLE_SEGMENT|2620,2627|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2631,2640|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|SIMPLE_SEGMENT|2633,2640|false|false|false|||minutes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2642,2650|false|false|false|C2706915||Language
Event|Event|SIMPLE_SEGMENT|2642,2650|false|false|false|||Language
Finding|Intellectual Product|SIMPLE_SEGMENT|2642,2650|false|false|false|C0033348|Programming Languages|Language
Event|Event|SIMPLE_SEGMENT|2652,2658|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|2652,2658|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2652,2658|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|2662,2668|false|false|false|||fluent
Finding|Idea or Concept|SIMPLE_SEGMENT|2670,2674|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|2675,2688|false|false|false|||comprehension
Finding|Mental Process|SIMPLE_SEGMENT|2675,2688|false|false|false|C0162340|Comprehension|comprehension
Event|Event|SIMPLE_SEGMENT|2690,2700|false|false|false|||Difficulty
Finding|Finding|SIMPLE_SEGMENT|2690,2700|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Finding|Finding|SIMPLE_SEGMENT|2690,2705|false|false|false|C0332218|Difficult (qualifier value)|Difficulty with
Event|Event|SIMPLE_SEGMENT|2706,2716|false|false|false|||repitition
Event|Event|SIMPLE_SEGMENT|2718,2724|false|false|false|||Naming
Finding|Mental Process|SIMPLE_SEGMENT|2718,2724|false|false|false|C0233735|Naming (function)|Naming
Event|Event|SIMPLE_SEGMENT|2725,2731|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2725,2731|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2736,2746|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|SIMPLE_SEGMENT|2736,2746|true|false|false|||dysarthria
Event|Event|SIMPLE_SEGMENT|2761,2767|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2770,2777|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2770,2784|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2770,2784|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2778,2784|false|false|false|C0027740|Nerve|Nerves
Event|Event|SIMPLE_SEGMENT|2793,2799|true|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2804,2810|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|2819,2824|false|false|false|||round
Event|Event|SIMPLE_SEGMENT|2829,2837|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2829,2837|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|SIMPLE_SEGMENT|2829,2846|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2841,2846|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2841,2846|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|2841,2846|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2841,2846|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2841,2846|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|SIMPLE_SEGMENT|2867,2873|false|false|false|C0234621|Visual|Visual
Event|Event|SIMPLE_SEGMENT|2874,2880|false|false|false|||fields
Event|Event|SIMPLE_SEGMENT|2885,2889|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|2893,2906|false|false|false|||confrontation
Finding|Finding|SIMPLE_SEGMENT|2893,2906|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2893,2906|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2893,2906|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|SIMPLE_SEGMENT|2921,2932|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2921,2942|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|SIMPLE_SEGMENT|2933,2942|true|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2933,2942|true|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2943,2949|true|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2943,2949|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2970,2979|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|SIMPLE_SEGMENT|2970,2979|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2984,2987|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|2984,2987|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2989,2995|false|false|false|C0015450|Face|Facial
Event|Event|SIMPLE_SEGMENT|2996,3004|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|2996,3004|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3009,3018|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|3009,3018|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3009,3018|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3009,3018|false|false|false|C2229507|sensory exam|sensation
Event|Event|SIMPLE_SEGMENT|3019,3025|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3019,3025|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3030,3039|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3030,3039|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3030,3039|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3041,3045|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|SIMPLE_SEGMENT|3041,3045|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|SIMPLE_SEGMENT|3041,3045|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|SIMPLE_SEGMENT|3047,3054|false|false|false|||Hearing
Finding|Finding|SIMPLE_SEGMENT|3047,3054|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|3047,3054|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|SIMPLE_SEGMENT|3055,3061|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3055,3061|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3065,3070|false|false|false|||voice
Finding|Idea or Concept|SIMPLE_SEGMENT|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|SIMPLE_SEGMENT|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|SIMPLE_SEGMENT|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3079,3086|false|false|false|C0700374|Palate|Palatal
Event|Event|SIMPLE_SEGMENT|3087,3096|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3087,3096|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|SIMPLE_SEGMENT|3097,3108|false|false|false|||symmetrical
Finding|Finding|SIMPLE_SEGMENT|3097,3108|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3114,3133|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3138,3147|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|SIMPLE_SEGMENT|3148,3154|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3173,3179|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3173,3179|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|3173,3179|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|SIMPLE_SEGMENT|3173,3187|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|SIMPLE_SEGMENT|3180,3187|true|false|false|C1660780|midline cell component|midline
Event|Event|SIMPLE_SEGMENT|3196,3210|true|false|false|||fasciculations
Finding|Sign or Symptom|SIMPLE_SEGMENT|3196,3210|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|SIMPLE_SEGMENT|3213,3218|false|false|false|||Motor
Finding|Functional Concept|SIMPLE_SEGMENT|3213,3218|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3227,3231|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|3227,3231|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|SIMPLE_SEGMENT|3227,3231|false|false|false|||bulk
Event|Event|SIMPLE_SEGMENT|3236,3240|false|false|false|||tone
Finding|Finding|SIMPLE_SEGMENT|3257,3265|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|3257,3265|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3257,3275|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|SIMPLE_SEGMENT|3257,3275|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|SIMPLE_SEGMENT|3266,3275|true|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|3266,3275|true|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|3277,3284|true|false|false|||tremors
Finding|Sign or Symptom|SIMPLE_SEGMENT|3277,3284|true|false|false|C0040822|Tremor|tremors
Finding|Idea or Concept|SIMPLE_SEGMENT|3286,3294|false|false|false|C0808080|Strength (attribute)|Strength
Finding|Social Behavior|SIMPLE_SEGMENT|3300,3305|false|false|false|C0032863|Power (Psychology)|power
Finding|Intellectual Product|SIMPLE_SEGMENT|3322,3326|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Pathologic Function|SIMPLE_SEGMENT|3335,3349|false|false|false|C1504476|Pronator drift|pronator drift
Event|Event|SIMPLE_SEGMENT|3344,3349|false|false|false|||drift
Finding|Finding|SIMPLE_SEGMENT|3351,3355|false|false|false|C0016928|Gait|Gait
Finding|Finding|SIMPLE_SEGMENT|3351,3364|false|false|false|C0231686|Gait, Unsteady|Gait unsteady
Event|Event|SIMPLE_SEGMENT|3356,3364|false|false|false|||unsteady
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3366,3379|false|false|false|C1656968|rhomberg test|rhomberg test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3375,3379|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|3375,3379|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|3375,3379|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|3375,3379|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3375,3379|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3375,3379|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|3385,3397|false|false|false|||unsteadiness
Finding|Finding|SIMPLE_SEGMENT|3385,3397|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|SIMPLE_SEGMENT|3400,3409|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|3400,3409|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3400,3409|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3400,3409|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|3411,3417|false|false|false|||Intact
Finding|Finding|SIMPLE_SEGMENT|3411,3417|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3421,3426|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3421,3426|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3421,3426|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3421,3426|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|3421,3432|false|false|false|C0423553|Light touch|light touch
Event|Event|SIMPLE_SEGMENT|3427,3432|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|3427,3432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3427,3432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3427,3432|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|3434,3447|false|false|false|||propioception
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3462,3471|false|false|false|C0677519|Exposed to vibration|vibration
Event|Event|SIMPLE_SEGMENT|3462,3471|false|false|false|||vibration
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3462,3471|false|false|false|C0459800||vibration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3462,3471|false|false|false|C0455941|Vibration - treatment|vibration
Event|Event|SIMPLE_SEGMENT|3486,3494|false|false|false|||Reflexes
Finding|Finding|SIMPLE_SEGMENT|3486,3494|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3486,3494|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3486,3494|false|false|false|C0436145|Examination of reflexes|Reflexes
Finding|Functional Concept|SIMPLE_SEGMENT|3509,3514|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|SIMPLE_SEGMENT|3528,3532|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3548,3552|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|SIMPLE_SEGMENT|3553,3562|false|false|false|||downgoing
Event|Event|SIMPLE_SEGMENT|3576,3588|false|false|false|||Coordination
Finding|Functional Concept|SIMPLE_SEGMENT|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3590,3594|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3598,3602|false|false|false|C0230444|Shin|shin
Event|Event|SIMPLE_SEGMENT|3603,3609|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3603,3609|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3611,3617|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3623,3629|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Event|Event|SIMPLE_SEGMENT|3630,3636|false|false|false|||slowed
Event|Event|SIMPLE_SEGMENT|3641,3653|false|false|false|||overshooting
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3659,3665|false|false|false|C0230370|Structure of right hand|R hand
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3661,3665|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|SIMPLE_SEGMENT|3661,3665|false|false|false|C0741992|Hand problem|hand
Event|Event|SIMPLE_SEGMENT|3667,3677|false|false|false|||Difficulty
Finding|Finding|SIMPLE_SEGMENT|3667,3677|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Finding|Finding|SIMPLE_SEGMENT|3667,3682|false|false|false|C0332218|Difficult (qualifier value)|Difficulty with
Event|Event|SIMPLE_SEGMENT|3689,3700|false|false|false|||alternating
Finding|Functional Concept|SIMPLE_SEGMENT|3689,3700|false|false|false|C0332270|Alternating|alternating
Event|Event|SIMPLE_SEGMENT|3701,3710|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|3701,3710|false|false|false|C0026649|Movement|movements
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3716,3722|false|false|false|C0230370|Structure of right hand|R hand
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3718,3722|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|SIMPLE_SEGMENT|3718,3722|false|false|false|C0741992|Hand problem|hand
Event|Event|SIMPLE_SEGMENT|3728,3737|false|false|false|||DISCHARGE
Finding|Body Substance|SIMPLE_SEGMENT|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3728,3737|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3746,3749|false|false|false|||VSS
Event|Event|SIMPLE_SEGMENT|3750,3753|false|false|false|||Gen
Finding|Classification|SIMPLE_SEGMENT|3750,3753|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|3750,3753|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3755,3758|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3755,3758|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3755,3758|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3755,3758|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3760,3765|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3767,3773|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|3781,3785|false|false|false|||EOMs
Finding|Functional Concept|SIMPLE_SEGMENT|3781,3785|false|false|false|C0241886|Extraocular|EOMs
Finding|Finding|SIMPLE_SEGMENT|3786,3792|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3797,3802|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|SIMPLE_SEGMENT|3804,3809|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3814,3821|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|3814,3821|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|SIMPLE_SEGMENT|3844,3863|false|false|false|C0232258|Pansystolic murmur|holosystolic murmur
Event|Event|SIMPLE_SEGMENT|3857,3863|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3857,3863|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3865,3868|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3865,3868|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3906,3911|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3906,3911|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3906,3911|true|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3915,3923|true|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|3915,3923|true|false|false|||erythema
Finding|Finding|SIMPLE_SEGMENT|3925,3929|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3925,3929|true|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3930,3934|true|false|false|C5575035|Well (answer to question)|well
Finding|Mental Process|SIMPLE_SEGMENT|3953,3959|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3953,3966|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|SIMPLE_SEGMENT|3953,3966|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3960,3966|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|3960,3966|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|3960,3966|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|3968,3973|false|false|false|||Awake
Finding|Finding|SIMPLE_SEGMENT|3968,3973|false|false|false|C0234422|Awake (finding)|Awake
Event|Event|SIMPLE_SEGMENT|3978,3989|false|false|false|||cooperative
Event|Event|SIMPLE_SEGMENT|3995,3999|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|3995,3999|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3995,3999|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|4008,4014|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|4008,4014|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|4008,4014|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|4016,4027|false|false|false|||Orientation
Finding|Mental Process|SIMPLE_SEGMENT|4016,4027|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|SIMPLE_SEGMENT|4029,4037|false|false|false|||Oriented
Finding|Finding|SIMPLE_SEGMENT|4029,4037|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|SIMPLE_SEGMENT|4029,4047|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4041,4047|false|false|false|C5890614||person
Event|Event|SIMPLE_SEGMENT|4041,4047|false|false|false|||person
Finding|Intellectual Product|SIMPLE_SEGMENT|4041,4047|false|false|false|C1522390|Person Info|person
Event|Activity|SIMPLE_SEGMENT|4049,4054|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|4049,4054|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|4049,4054|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4049,4054|false|false|false|C1533810||place
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4066,4074|false|false|false|C2706915||Language
Event|Event|SIMPLE_SEGMENT|4066,4074|false|false|false|||Language
Finding|Intellectual Product|SIMPLE_SEGMENT|4066,4074|false|false|false|C0033348|Programming Languages|Language
Event|Event|SIMPLE_SEGMENT|4076,4082|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|4076,4082|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4076,4082|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|4086,4092|false|false|false|||fluent
Finding|Idea or Concept|SIMPLE_SEGMENT|4094,4098|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|4099,4112|false|false|false|||comprehension
Finding|Mental Process|SIMPLE_SEGMENT|4099,4112|false|false|false|C0162340|Comprehension|comprehension
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4115,4122|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4115,4129|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4115,4129|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4123,4129|false|false|false|C0027740|Nerve|Nerves
Finding|Functional Concept|SIMPLE_SEGMENT|4138,4144|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|tested
Finding|Intellectual Product|SIMPLE_SEGMENT|4138,4144|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|tested
Event|Event|SIMPLE_SEGMENT|4149,4155|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|4149,4155|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|4161,4166|false|false|false|||Motor
Finding|Functional Concept|SIMPLE_SEGMENT|4161,4166|false|false|false|C1513492|motor movement|Motor
Event|Event|SIMPLE_SEGMENT|4172,4180|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|4172,4180|false|false|false|C0808080|Strength (attribute)|strength
Finding|Pathologic Function|SIMPLE_SEGMENT|4203,4217|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|SIMPLE_SEGMENT|4212,4217|true|false|false|||drift
Finding|Finding|SIMPLE_SEGMENT|4219,4223|true|false|false|C0016928|Gait|Gait
Event|Event|SIMPLE_SEGMENT|4233,4240|true|false|false|||walking
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|SIMPLE_SEGMENT|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|SIMPLE_SEGMENT|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Event|SIMPLE_SEGMENT|4249,4259|true|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|4249,4259|true|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|4262,4271|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|4262,4271|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4262,4271|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4262,4271|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|4281,4287|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|4281,4287|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|4294,4302|false|false|false|||Reflexes
Finding|Finding|SIMPLE_SEGMENT|4294,4302|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4294,4302|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4294,4302|false|false|false|C0436145|Examination of reflexes|Reflexes
Finding|Functional Concept|SIMPLE_SEGMENT|4317,4322|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|SIMPLE_SEGMENT|4336,4340|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4356,4360|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|SIMPLE_SEGMENT|4361,4370|false|false|false|||downgoing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4416,4421|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4416,4421|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4416,4421|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4422,4425|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4431,4434|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4431,4434|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4431,4434|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4441,4444|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4441,4444|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4441,4444|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4441,4444|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4451,4454|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4451,4454|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4461,4464|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4461,4464|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4461,4464|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4461,4464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4461,4464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4468,4471|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4468,4471|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4468,4471|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4468,4471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4468,4471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4468,4471|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4477,4481|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4477,4481|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4496,4499|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4516,4521|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4516,4521|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4516,4521|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4538,4543|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4538,4543|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4538,4543|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4538,4551|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4538,4551|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4538,4551|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4544,4551|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4544,4551|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4544,4551|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4544,4551|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4544,4551|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4544,4551|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4598,4602|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4598,4602|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4598,4602|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4627,4632|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4627,4632|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4627,4632|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4627,4640|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|4633,4640|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|4633,4640|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|4633,4640|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4633,4640|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4658,4663|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4658,4663|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4658,4663|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4665,4670|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4665,4670|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|SIMPLE_SEGMENT|4665,4670|false|false|false|||HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4665,4670|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|SIMPLE_SEGMENT|4676,4679|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4697,4702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4697,4702|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4697,4702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4717,4724|false|false|false|C0881943||CT Head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4717,4724|false|false|false|C0202691|CAT scan of head|CT Head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4720,4724|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4720,4724|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4720,4724|false|false|false|C0362076|Problems with head|Head
Event|Event|SIMPLE_SEGMENT|4720,4724|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4720,4724|false|false|false|C0876917|Procedure on head|Head
Event|Event|SIMPLE_SEGMENT|4731,4741|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4731,4741|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4731,4741|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|4759,4765|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|4759,4765|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|4759,4765|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|4778,4782|false|false|false|||foci
Finding|Finding|SIMPLE_SEGMENT|4778,4782|false|false|false|C4321394|Foci|foci
Event|Event|SIMPLE_SEGMENT|4786,4800|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|4786,4800|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4786,4800|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Event|Event|SIMPLE_SEGMENT|4802,4811|false|false|false|||measuring
Finding|Finding|SIMPLE_SEGMENT|4830,4836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4830,4836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|4837,4845|false|false|false|||reflects
Event|Event|SIMPLE_SEGMENT|4861,4865|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4877,4887|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|SIMPLE_SEGMENT|4877,4887|false|false|false|||meningioma
Event|Event|SIMPLE_SEGMENT|4905,4913|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|4905,4913|false|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|4930,4938|false|false|false|||subacute
Event|Event|SIMPLE_SEGMENT|4942,4949|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|4942,4949|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|4942,4949|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|SIMPLE_SEGMENT|4955,4965|false|false|false|||considered
Event|Event|SIMPLE_SEGMENT|4971,4977|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|4971,4977|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4971,4977|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|4983,4987|false|false|false|||Loss
Finding|Finding|SIMPLE_SEGMENT|4983,4987|false|false|false|C5890125|Loss (adaptation)|Loss
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5002,5017|false|false|false|C1511938|Cellular Differentiation Qualifier|differentiation
Event|Event|SIMPLE_SEGMENT|5002,5017|false|false|false|||differentiation
Finding|Cell Function|SIMPLE_SEGMENT|5002,5017|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Finding|Functional Concept|SIMPLE_SEGMENT|5002,5017|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Finding|Finding|SIMPLE_SEGMENT|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Functional Concept|SIMPLE_SEGMENT|5030,5034|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5051,5055|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|5051,5055|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|5063,5070|false|false|false|||reflect
Finding|Intellectual Product|SIMPLE_SEGMENT|5074,5079|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|SIMPLE_SEGMENT|5074,5087|false|false|false|C0333548|Acute infarct|acute infarct
Event|Event|SIMPLE_SEGMENT|5080,5087|false|false|false|||infarct
Finding|Pathologic Function|SIMPLE_SEGMENT|5080,5087|false|false|false|C0021308|Infarction|infarct
Event|Event|SIMPLE_SEGMENT|5091,5094|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|5091,5094|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5091,5094|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|5091,5094|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5091,5099|false|false|false|C0412674|MRI of head|MRI Head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5095,5099|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5095,5099|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5095,5099|false|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5095,5099|false|false|false|C0876917|Procedure on head|Head
Event|Event|SIMPLE_SEGMENT|5105,5110|false|false|false|||Acute
Finding|Intellectual Product|SIMPLE_SEGMENT|5105,5110|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Event|Event|SIMPLE_SEGMENT|5133,5144|false|false|false|||infarctions
Finding|Pathologic Function|SIMPLE_SEGMENT|5133,5144|false|false|false|C0021308|Infarction|infarctions
Event|Event|SIMPLE_SEGMENT|5162,5167|false|false|false|||focus
Finding|Functional Concept|SIMPLE_SEGMENT|5162,5167|false|false|false|C1285542|Has focus|focus
Finding|Functional Concept|SIMPLE_SEGMENT|5176,5180|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5201,5211|false|false|false|C0550215||Appearance
Event|Event|SIMPLE_SEGMENT|5201,5211|false|false|false|||Appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|5201,5211|false|false|false|C2051406|patient appearance regarding mental status exam|Appearance
Event|Event|SIMPLE_SEGMENT|5231,5237|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|5231,5237|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|5231,5237|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|5241,5249|false|false|false|||somewhat
Finding|Finding|SIMPLE_SEGMENT|5241,5249|false|false|false|C2984079|Somewhat|somewhat
Event|Event|SIMPLE_SEGMENT|5277,5286|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|5287,5296|false|false|false|||attention
Finding|Intellectual Product|SIMPLE_SEGMENT|5287,5296|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|SIMPLE_SEGMENT|5287,5296|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Event|Event|SIMPLE_SEGMENT|5300,5308|true|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|5300,5308|true|false|false|C1522577|follow-up|followup
Event|Event|SIMPLE_SEGMENT|5310,5317|true|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|5310,5317|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5310,5317|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|5330,5340|true|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|5330,5340|true|true|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5330,5340|true|true|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|5344,5351|false|false|false|||exclude
Event|Event|SIMPLE_SEGMENT|5356,5364|true|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5356,5364|true|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|SIMPLE_SEGMENT|5356,5367|true|false|false|C0150312|Present|presence of
Event|Event|SIMPLE_SEGMENT|5383,5387|true|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5393,5404|true|false|false|C0025286|Meningioma|meningiomas
Event|Event|SIMPLE_SEGMENT|5393,5404|true|false|false|||meningiomas
Finding|Functional Concept|SIMPLE_SEGMENT|5412,5416|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5417,5431|true|false|false|C0016733;C0162783;C0549224|Frontal region;Prefrontal Cortex;frontal lobe|frontal region
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5417,5431|true|false|false|C0016733;C0162783;C0549224|Frontal region;Prefrontal Cortex;frontal lobe|frontal region
Drug|Amino Acid Sequence|SIMPLE_SEGMENT|5425,5431|true|false|false|C1514562|Protein Domain|region
Finding|Idea or Concept|SIMPLE_SEGMENT|5441,5452|true|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|5453,5457|true|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|5453,5464|true|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|5458,5464|true|false|false|||effect
Event|Event|SIMPLE_SEGMENT|5467,5471|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|5467,5471|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5467,5471|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Conceptual Entity|SIMPLE_SEGMENT|5484,5493|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|5484,5493|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Functional Concept|SIMPLE_SEGMENT|5494,5498|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5494,5522|false|false|false|C3484363||left ventricular hypertrophy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5494,5522|false|false|false|C0149721|Left Ventricular Hypertrophy|left ventricular hypertrophy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5499,5510|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5499,5522|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|SIMPLE_SEGMENT|5511,5522|false|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|5511,5522|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5535,5541|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5535,5541|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5535,5541|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5568,5576|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5577,5585|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5587,5591|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5592,5598|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5592,5604|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5599,5604|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5606,5614|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5606,5614|false|false|false|C1261287|Stenosis|stenosis
Finding|Intellectual Product|SIMPLE_SEGMENT|5616,5620|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5621,5627|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5621,5641|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|SIMPLE_SEGMENT|5628,5641|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5628,5641|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5628,5641|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5628,5641|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Functional Concept|SIMPLE_SEGMENT|5643,5648|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5643,5670|false|false|false|C4288280|Right Ventricular Free Wall|Right ventricular free wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5649,5660|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|5661,5665|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5661,5665|false|false|false|C0332296|Free of (attribute)|free
Event|Event|SIMPLE_SEGMENT|5672,5683|false|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|5672,5683|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5685,5694|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5685,5694|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|5685,5694|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5685,5701|false|false|false|C0034052|Pulmonary artery structure|Pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5695,5701|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5695,5701|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5702,5710|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5702,5723|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5711,5723|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5711,5723|false|false|false|||hypertension
Finding|Finding|SIMPLE_SEGMENT|5725,5732|false|false|false|C0700124|Dilated|Dilated
Finding|Functional Concept|SIMPLE_SEGMENT|5734,5743|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5734,5749|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5744,5749|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|5744,5749|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Intellectual Product|SIMPLE_SEGMENT|5752,5760|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|CLINICAL
Finding|Body Substance|SIMPLE_SEGMENT|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|5780,5791|false|false|false|C0332310|Has patient|patient has
Finding|Intellectual Product|SIMPLE_SEGMENT|5792,5796|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5797,5803|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|SIMPLE_SEGMENT|5797,5812|false|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|SIMPLE_SEGMENT|5804,5812|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5804,5812|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5827,5830|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Anatomy|Tissue|SIMPLE_SEGMENT|5827,5830|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5827,5830|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5827,5830|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Enzyme|SIMPLE_SEGMENT|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Event|Event|SIMPLE_SEGMENT|5827,5830|false|false|false|||ACC
Finding|Gene or Genome|SIMPLE_SEGMENT|5827,5830|false|false|false|C1412104;C3541413|ACACA gene;ACACA wt Allele|ACC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5831,5834|false|false|false|C0002880;C0272325|Autoimmune hemolytic anemia;Factor 8 deficiency, acquired|AHA
Drug|Organic Chemical|SIMPLE_SEGMENT|5831,5834|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5831,5834|false|false|false|C0050451|acetohydroxamic acid|AHA
Event|Event|SIMPLE_SEGMENT|5831,5834|false|false|false|||AHA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5836,5858|false|false|false|C0018824|Heart valve disease|Valvular Heart Disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5845,5850|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5845,5850|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5845,5850|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5845,5858|false|false|false|C0018799|Heart Diseases|Heart Disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5851,5858|false|false|false|C0012634|Disease|Disease
Event|Event|SIMPLE_SEGMENT|5859,5869|false|false|false|||Guidelines
Finding|Intellectual Product|SIMPLE_SEGMENT|5859,5869|false|false|false|C0162791;C0220845;C0282423|Guideline (Publication Type);Guidelines;guiding characteristics|Guidelines
Event|Event|SIMPLE_SEGMENT|5873,5879|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|5873,5879|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5873,5879|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5873,5882|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5873,5882|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|5883,5897|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5883,5897|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|5902,5911|false|false|false|||suggested
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5944,5956|false|false|false|C0014118|Endocarditis|endocarditis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5944,5968|false|false|false|C1396567|Endocarditis prophylaxis|endocarditis prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5957,5968|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|5969,5984|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|5969,5984|false|false|false|C0034866|Recommendation|recommendations
Procedure|Health Care Activity|SIMPLE_SEGMENT|5991,5995|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5991,5995|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5996,6004|true|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|5996,6004|true|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|5996,6004|true|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|6014,6025|true|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6014,6025|true|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|6033,6044|true|false|false|||recommended
Finding|Intellectual Product|SIMPLE_SEGMENT|6046,6054|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|Clinical
Event|Event|SIMPLE_SEGMENT|6056,6065|false|false|false|||decisions
Finding|Mental Process|SIMPLE_SEGMENT|6056,6065|false|false|false|C0679006|Decision|decisions
Event|Event|SIMPLE_SEGMENT|6080,6084|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|6080,6084|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|6080,6088|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|SIMPLE_SEGMENT|6089,6100|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6089,6100|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|6111,6116|false|false|false|||based
Event|Event|SIMPLE_SEGMENT|6121,6129|false|false|false|||clinical
Finding|Intellectual Product|SIMPLE_SEGMENT|6121,6129|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|SIMPLE_SEGMENT|6152,6156|false|false|false|||data
Finding|Idea or Concept|SIMPLE_SEGMENT|6152,6156|false|false|false|C1511726|Data|data
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Event|Event|SIMPLE_SEGMENT|6160,6163|false|false|false|||MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6160,6163|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6160,6163|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6160,6168|false|false|false|C1636167|Magnetic resonance angiography of vascular structure of head|MRA Head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6164,6168|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6164,6168|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6164,6168|false|false|false|C0362076|Problems with head|Head
Event|Event|SIMPLE_SEGMENT|6164,6168|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6164,6168|false|false|false|C0876917|Procedure on head|Head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6169,6173|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|6169,6173|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|6169,6173|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Intellectual Product|SIMPLE_SEGMENT|6179,6183|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Functional Concept|SIMPLE_SEGMENT|6184,6199|false|false|false|C0333482|atherosclerotic|atherosclerotic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6200,6207|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6200,6207|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6215,6229|false|false|false|C0004811|Structure of basilar artery|basilar artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6223,6229|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6223,6229|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|6244,6252|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|6244,6252|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6244,6255|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|SIMPLE_SEGMENT|6256,6261|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6262,6270|true|false|false|C0005847|Blood Vessel|vascular
Finding|Finding|SIMPLE_SEGMENT|6262,6284|true|false|false|C0241657|Abnormality of the vasculature|vascular abnormalities
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6271,6284|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|6271,6284|true|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|6271,6284|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|6285,6294|true|false|false|||involving
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6300,6312|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|6300,6312|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6313,6321|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|6313,6321|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|6313,6321|false|false|false|C0397581|Procedure on artery|arteries
Finding|Intellectual Product|SIMPLE_SEGMENT|6329,6334|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6335,6343|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6335,6350|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6335,6350|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|6364,6372|false|false|false|||admitted
Event|Occupational Activity|SIMPLE_SEGMENT|6394,6401|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|6394,6401|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|SIMPLE_SEGMENT|6419,6428|false|false|false|||emergency
Finding|Finding|SIMPLE_SEGMENT|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6419,6428|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|6419,6428|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|6419,6433|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Event|Event|SIMPLE_SEGMENT|6449,6455|false|false|false|||series
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6459,6464|false|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|6459,6464|false|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|6459,6464|false|false|false|C0085639|Falls|falls
Event|Event|SIMPLE_SEGMENT|6476,6478|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6486,6490|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6486,6490|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6486,6490|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6486,6490|false|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|6491,6503|false|false|false|||demonstrated
Finding|Functional Concept|SIMPLE_SEGMENT|6506,6510|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|6532,6536|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|6540,6544|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|SIMPLE_SEGMENT|6555,6560|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|6561,6567|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|6561,6567|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|6561,6567|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6585,6589|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6585,6589|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Functional Concept|SIMPLE_SEGMENT|6597,6601|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6625,6630|false|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|6625,6630|false|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|6625,6630|false|false|false|C0085639|Falls|falls
Drug|Organic Chemical|SIMPLE_SEGMENT|6636,6644|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6636,6644|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|6636,6644|false|false|false|||coumadin
Event|Event|SIMPLE_SEGMENT|6650,6654|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|6666,6672|false|false|false|||placed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|6679,6686|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|6679,6686|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6679,6686|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|6687,6694|false|false|false|||sliding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6695,6700|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|6695,6700|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|6695,6700|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|6695,6700|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|SIMPLE_SEGMENT|6720,6727|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|6720,6727|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6732,6744|false|true|false|C0020615|Hypoglycemia|hypoglycemia
Event|Event|SIMPLE_SEGMENT|6732,6744|false|false|false|||hypoglycemia
Finding|Finding|SIMPLE_SEGMENT|6732,6744|false|true|false|C5767385|Blood glucose below reference range (finding)|hypoglycemia
Event|Event|SIMPLE_SEGMENT|6745,6757|false|false|false|||contributing
Event|Event|SIMPLE_SEGMENT|6765,6777|false|false|false|||unsteadiness
Finding|Finding|SIMPLE_SEGMENT|6765,6777|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|SIMPLE_SEGMENT|6784,6787|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|6784,6787|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6784,6787|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|6784,6787|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6796,6800|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6796,6800|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6796,6800|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6796,6800|false|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|6805,6813|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|6820,6829|false|false|false|||confirmed
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6832,6842|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|SIMPLE_SEGMENT|6832,6842|false|false|false|||meningioma
Event|Event|SIMPLE_SEGMENT|6844,6853|false|false|false|||overlying
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6860,6872|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6860,6872|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6868,6872|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6868,6872|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|6889,6896|false|false|false|||infarct
Finding|Pathologic Function|SIMPLE_SEGMENT|6889,6896|false|false|false|C0021308|Infarction|infarct
Event|Event|SIMPLE_SEGMENT|6918,6923|false|false|false|||gyrus
Finding|Functional Concept|SIMPLE_SEGMENT|6931,6935|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|6964,6969|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|6977,6985|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6977,6985|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6993,7002|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|6993,7002|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|6993,7007|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Finding|Idea or Concept|SIMPLE_SEGMENT|7012,7020|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|7021,7024|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7021,7024|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|7034,7042|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7034,7042|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Intellectual Product|SIMPLE_SEGMENT|7054,7064|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|7065,7073|false|false|false|||resolved
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7082,7091|false|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|7082,7091|false|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|7082,7091|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|7102,7108|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|7102,7108|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|7122,7129|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|7122,7129|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|7134,7142|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|7155,7163|false|false|false|||appeared
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7182,7188|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|7182,7188|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|7182,7188|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|SIMPLE_SEGMENT|7196,7199|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|7196,7199|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7196,7199|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|7196,7199|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|7207,7218|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|7220,7230|false|false|false|||restarting
Drug|Organic Chemical|SIMPLE_SEGMENT|7240,7248|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7240,7248|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|7240,7248|false|false|false|||coumadin
Event|Event|SIMPLE_SEGMENT|7250,7257|false|false|false|||holding
Drug|Organic Chemical|SIMPLE_SEGMENT|7262,7270|false|false|false|C0699512|Dilantin|dilantin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7262,7270|false|false|false|C0699512|Dilantin|dilantin
Event|Event|SIMPLE_SEGMENT|7262,7270|false|false|false|||dilantin
Event|Activity|SIMPLE_SEGMENT|7275,7283|false|false|false|C1283174||checking
Event|Event|SIMPLE_SEGMENT|7275,7283|false|false|false|||checking
Event|Event|SIMPLE_SEGMENT|7288,7291|false|false|false|||EEG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7288,7291|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|SIMPLE_SEGMENT|7325,7334|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7325,7334|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|7325,7334|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|7365,7369|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|7365,7369|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7365,7369|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Event|Event|SIMPLE_SEGMENT|7377,7380|false|false|false|||MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7377,7380|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7377,7380|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7388,7393|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7388,7393|false|false|false|C0006111|Brain Diseases|brain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7398,7402|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|7398,7402|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|7398,7402|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|SIMPLE_SEGMENT|7414,7420|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7414,7420|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Pathologic Function|SIMPLE_SEGMENT|7421,7428|false|true|false|C0013922|Embolism|embolic
Event|Event|SIMPLE_SEGMENT|7429,7435|false|false|false|||nature
Finding|Functional Concept|SIMPLE_SEGMENT|7429,7435|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|7429,7435|false|false|false|C0349590;C1262865|Nature;Natures|nature
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7443,7450|false|false|false|C0038454|Cerebrovascular accident|strokes
Event|Event|SIMPLE_SEGMENT|7443,7450|false|false|false|||strokes
Event|Event|SIMPLE_SEGMENT|7469,7472|false|false|false|||see
Finding|Functional Concept|SIMPLE_SEGMENT|7496,7502|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7503,7507|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7503,7507|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7503,7507|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7503,7507|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7503,7511|false|false|false|C0412674|MRI of head|head MRI
Event|Event|SIMPLE_SEGMENT|7508,7511|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|7508,7511|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7508,7511|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|7508,7511|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|7523,7526|false|false|false|||saw
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7539,7547|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|7548,7557|false|false|false|||managment
Event|Event|SIMPLE_SEGMENT|7563,7574|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|7575,7583|false|false|false|||changing
Drug|Organic Chemical|SIMPLE_SEGMENT|7588,7597|true|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7588,7597|true|false|false|C0017642|glipizide|glipizide
Event|Event|SIMPLE_SEGMENT|7588,7597|true|false|false|||glipizide
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7604,7607|true|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7604,7607|true|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7604,7607|true|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7604,7607|true|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7604,7607|true|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|7618,7626|true|false|false|||starting
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|7627,7634|true|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7627,7634|true|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7627,7634|true|false|false|C0202098|Insulin measurement|insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|7640,7646|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7640,7646|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|7640,7646|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7640,7646|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|7652,7656|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|7657,7667|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|7708,7716|true|false|false|||episodes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7720,7732|true|false|false|C0020615|Hypoglycemia|hypoglycemia
Event|Event|SIMPLE_SEGMENT|7720,7732|true|false|false|||hypoglycemia
Finding|Finding|SIMPLE_SEGMENT|7720,7732|true|false|false|C5767385|Blood glucose below reference range (finding)|hypoglycemia
Event|Event|SIMPLE_SEGMENT|7753,7763|false|false|false|||standpoing
Finding|Idea or Concept|SIMPLE_SEGMENT|7765,7773|false|false|false|C4288901|In-House|in-house
Event|Event|SIMPLE_SEGMENT|7787,7791|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|7787,7791|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|7797,7806|false|false|false|||resultion
Finding|Functional Concept|SIMPLE_SEGMENT|7815,7820|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|SIMPLE_SEGMENT|7815,7835|false|false|false|C0457435|Right hemiparesis|right sided weakness
Event|Event|SIMPLE_SEGMENT|7827,7835|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7827,7835|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|7849,7861|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|SIMPLE_SEGMENT|7862,7871|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7862,7871|false|false|false|C0549178|Continuous|continued
Event|Event|SIMPLE_SEGMENT|7880,7886|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7887,7894|false|false|false|C1317973|Support - dental|support
Drug|Organic Chemical|SIMPLE_SEGMENT|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Vitamin|SIMPLE_SEGMENT|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Event|Event|SIMPLE_SEGMENT|7887,7894|false|false|false|||support
Finding|Conceptual Entity|SIMPLE_SEGMENT|7887,7894|false|false|false|C1521721|Supportive assistance|support
Procedure|Health Care Activity|SIMPLE_SEGMENT|7887,7894|false|false|false|C0344211|Supportive care|support
Event|Event|SIMPLE_SEGMENT|7901,7911|false|false|false|||ambulating
Event|Event|SIMPLE_SEGMENT|7919,7930|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|7934,7936|false|false|false|||go
Finding|Idea or Concept|SIMPLE_SEGMENT|7948,7952|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|7948,7952|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Event|Event|SIMPLE_SEGMENT|7953,7958|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7953,7958|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|7972,7978|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|7972,7978|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|7980,7984|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|7980,7984|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|7988,7995|false|false|false|||compete
Event|Event|SIMPLE_SEGMENT|7996,8005|false|false|false|||transfers
Finding|Finding|SIMPLE_SEGMENT|7996,8005|false|false|false|C0728827|transfers|transfers
Event|Event|SIMPLE_SEGMENT|8010,8018|false|false|false|||ambulate
Finding|Finding|SIMPLE_SEGMENT|8010,8018|false|false|false|C4036205|Ambulate|ambulate
Event|Event|SIMPLE_SEGMENT|8043,8049|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|8058,8067|false|false|false|||neurology
Event|Event|SIMPLE_SEGMENT|8072,8084|false|false|false|||neurosurgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8072,8084|false|false|false|C0524850|Neurosurgical Procedures|neurosurgery
Event|Event|SIMPLE_SEGMENT|8088,8095|false|false|false|||discuss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8103,8107|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|8103,8107|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|8103,8107|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|SIMPLE_SEGMENT|8109,8115|false|false|false|||manage
Finding|Functional Concept|SIMPLE_SEGMENT|8120,8128|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8120,8136|false|false|false|C0948008|Ischemic stroke|ischemic strokes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8129,8136|false|false|false|C0038454|Cerebrovascular accident|strokes
Event|Event|SIMPLE_SEGMENT|8129,8136|false|false|false|||strokes
Event|Event|SIMPLE_SEGMENT|8141,8148|false|false|false|||address
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8153,8163|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|SIMPLE_SEGMENT|8153,8163|false|false|false|||meningioma
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8182,8193|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8182,8193|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8182,8193|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8182,8193|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8182,8206|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8197,8206|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8197,8206|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|8208,8216|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8208,8216|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|8208,8216|false|false|false|||Coumadin
Event|Event|SIMPLE_SEGMENT|8220,8221|false|false|false|||'
Drug|Organic Chemical|SIMPLE_SEGMENT|8223,8230|false|false|false|C0722725|Prandin|prandin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8223,8230|false|false|false|C0722725|Prandin|prandin
Event|Event|SIMPLE_SEGMENT|8223,8230|false|false|false|||prandin
Drug|Organic Chemical|SIMPLE_SEGMENT|8239,8248|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8239,8248|false|false|false|C0017642|glipizide|glipizide
Event|Event|SIMPLE_SEGMENT|8239,8248|false|false|false|||glipizide
Drug|Organic Chemical|SIMPLE_SEGMENT|8254,8264|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8254,8264|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|8254,8264|false|false|false|||isosorbide
Event|Event|SIMPLE_SEGMENT|8266,8275|false|false|false|||dinitrate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8282,8292|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8282,8292|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|8282,8292|false|false|false|||lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|8297,8308|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8297,8308|false|false|false|C0002144|allopurinol|allopurinol
Event|Event|SIMPLE_SEGMENT|8297,8308|false|false|false|||allopurinol
Drug|Organic Chemical|SIMPLE_SEGMENT|8314,8323|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8314,8323|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|8314,8323|false|false|false|||torsemide
Drug|Organic Chemical|SIMPLE_SEGMENT|8328,8338|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8328,8338|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8328,8338|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8346,8353|false|false|false|C0593906|Lipitor|lipitor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8346,8353|false|false|false|C0593906|Lipitor|lipitor
Event|Event|SIMPLE_SEGMENT|8346,8353|false|false|false|||lipitor
Event|Event|SIMPLE_SEGMENT|8361,8370|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8361,8370|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8361,8382|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8371,8382|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8371,8382|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8371,8382|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8371,8382|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8387,8397|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8387,8397|false|false|false|C0022251|isosorbide|Isosorbide
Event|Event|SIMPLE_SEGMENT|8387,8397|false|false|false|||Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8387,8407|false|false|false|C0022252|isosorbide dinitrate|Isosorbide Dinitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8387,8407|false|false|false|C0022252|isosorbide dinitrate|Isosorbide Dinitrate
Event|Event|SIMPLE_SEGMENT|8398,8407|false|false|false|||Dinitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8414,8420|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8434,8440|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8434,8440|false|false|false|||Tablet
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8444,8447|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8444,8447|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8444,8447|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8444,8447|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8444,8447|false|false|false|C1332410|BID gene|BID
Finding|Finding|SIMPLE_SEGMENT|8450,8457|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8452,8457|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|8460,8463|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8460,8463|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8471,8481|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8471,8481|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8488,8494|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8508,8514|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8508,8514|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|8539,8549|false|false|false|||Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8565,8571|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8585,8591|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8585,8591|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8595,8598|false|false|false|||TID
Finding|Finding|SIMPLE_SEGMENT|8601,8608|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8603,8608|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|8603,8608|false|false|false|||times
Finding|Idea or Concept|SIMPLE_SEGMENT|8611,8614|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8611,8614|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|8622,8633|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8622,8633|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8640,8646|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8660,8666|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8667,8669|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|8691,8702|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8691,8702|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8710,8716|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8730,8736|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8730,8736|false|false|false|||Tablet
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8777,8783|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8797,8803|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8804,8806|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|8834,8843|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8834,8843|false|false|false|C0076840|torsemide|Torsemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8849,8855|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8869,8875|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8869,8875|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|8899,8908|false|false|false|C0017642|glipizide|Glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8899,8908|false|false|false|C0017642|glipizide|Glipizide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8915,8921|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8935,8941|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8935,8941|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8942,8944|false|false|false|||PO
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8945,8948|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8945,8948|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8945,8948|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8945,8948|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8945,8948|false|false|false|C1332410|BID gene|BID
Finding|Finding|SIMPLE_SEGMENT|8950,8957|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8952,8957|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|8952,8957|false|false|false|||times
Finding|Idea or Concept|SIMPLE_SEGMENT|8961,8964|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8961,8964|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|8972,8981|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8972,8981|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8972,8993|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8972,8993|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8982,8993|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8982,8993|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8982,8993|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|8995,9003|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8995,9003|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|8995,9008|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|9004,9008|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|9004,9008|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|9004,9008|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|9004,9008|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|9011,9019|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9011,9019|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|9025,9034|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9025,9034|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9025,9044|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9035,9044|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9035,9044|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9035,9044|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9035,9044|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9035,9044|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9046,9050|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9059,9069|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|SIMPLE_SEGMENT|9059,9069|false|false|false|||meningioma
Finding|Functional Concept|SIMPLE_SEGMENT|9071,9075|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|9095,9102|false|false|false|||infarct
Finding|Pathologic Function|SIMPLE_SEGMENT|9095,9102|false|false|false|C0021308|Infarction|infarct
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9105,9113|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|9105,9113|false|false|false|||Diabetes
Event|Event|SIMPLE_SEGMENT|9117,9126|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9117,9126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9117,9126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9117,9126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9117,9126|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9127,9136|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9127,9136|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9127,9136|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9127,9136|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9138,9144|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9138,9151|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9138,9151|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9145,9151|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9145,9151|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9153,9161|false|false|false|C0009676|Confusion|Confused
Event|Event|SIMPLE_SEGMENT|9153,9161|false|false|false|||Confused
Finding|Finding|SIMPLE_SEGMENT|9153,9161|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|9153,9161|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Event|SIMPLE_SEGMENT|9175,9180|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9175,9197|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9175,9197|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9184,9197|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9184,9197|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9184,9197|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9199,9204|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|9199,9204|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9199,9204|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|9199,9204|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|9209,9220|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|9209,9220|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|9222,9230|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9222,9230|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9222,9230|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9231,9237|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9231,9237|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9231,9237|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9239,9249|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9252,9260|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|9261,9271|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|9261,9271|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9275,9278|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|9275,9278|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|SIMPLE_SEGMENT|9275,9278|false|false|false|||aid
Finding|Gene or Genome|SIMPLE_SEGMENT|9275,9278|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9275,9278|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|SIMPLE_SEGMENT|9280,9286|false|false|false|||walker
Event|Event|SIMPLE_SEGMENT|9301,9310|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9301,9310|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9301,9323|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9301,9323|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9301,9323|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9311,9323|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9311,9323|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9311,9323|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|9336,9340|false|false|false|||take
Drug|Organic Chemical|SIMPLE_SEGMENT|9346,9354|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9346,9354|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|9346,9354|false|false|false|||coumadin
Event|Event|SIMPLE_SEGMENT|9358,9368|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|9381,9385|true|false|false|||need
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9399,9410|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9399,9410|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9399,9410|true|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9399,9410|true|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9434,9440|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|9469,9475|false|false|false|||listed
Event|Event|SIMPLE_SEGMENT|9492,9496|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|9499,9505|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|9499,9505|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|9499,9508|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|9499,9508|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|9509,9512|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|9509,9512|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9509,9512|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|9509,9512|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|9516,9524|false|false|false|||evaluate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9536,9542|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|9536,9542|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|9536,9542|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Functional Concept|SIMPLE_SEGMENT|9558,9562|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9576,9581|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9576,9581|false|false|false|C0006111|Brain Diseases|brain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9593,9604|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9593,9604|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9593,9604|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9593,9604|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9608,9618|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|9623,9629|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|9652,9656|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|9660,9665|false|false|false|||check
Finding|Classification|SIMPLE_SEGMENT|9671,9678|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|9671,9678|false|false|false|C3812897|General medical service|General
Finding|Idea or Concept|SIMPLE_SEGMENT|9671,9691|false|false|false|C1549999|General Instructions|General Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9679,9691|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9679,9691|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9679,9691|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Idea or Concept|SIMPLE_SEGMENT|9692,9703|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|Information
Finding|Intellectual Product|SIMPLE_SEGMENT|9692,9703|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|Information
Event|Event|SIMPLE_SEGMENT|9705,9709|false|false|false|||Take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9715,9719|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9715,9719|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9715,9719|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9715,9719|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|SIMPLE_SEGMENT|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9720,9728|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|SIMPLE_SEGMENT|9720,9728|false|false|false|||medicine
Event|Event|SIMPLE_SEGMENT|9732,9742|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|9745,9753|false|false|false|||Exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9745,9753|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9745,9753|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|SIMPLE_SEGMENT|9764,9771|false|false|false|||limited
Event|Event|SIMPLE_SEGMENT|9775,9782|false|false|false|||walking
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|SIMPLE_SEGMENT|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|SIMPLE_SEGMENT|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Activity|SIMPLE_SEGMENT|9787,9794|true|false|false|C0206244|Lifting|lifting
Event|Event|SIMPLE_SEGMENT|9787,9794|true|false|false|||lifting
Event|Event|SIMPLE_SEGMENT|9796,9805|true|false|false|||straining
Finding|Physiologic Function|SIMPLE_SEGMENT|9796,9805|true|false|false|C0442694|Straining (finding)|straining
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9821,9828|false|false|false|C0011119|Decompression Sickness|bending
Event|Event|SIMPLE_SEGMENT|9821,9828|false|false|false|||bending
Finding|Finding|SIMPLE_SEGMENT|9821,9828|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|SIMPLE_SEGMENT|9821,9828|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|SIMPLE_SEGMENT|9831,9839|false|false|false|||Increase
Event|Event|SIMPLE_SEGMENT|9845,9851|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|9845,9851|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|9845,9851|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Substance|SIMPLE_SEGMENT|9855,9861|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|9855,9861|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|9855,9861|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9855,9861|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Tissue|SIMPLE_SEGMENT|9866,9871|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|SIMPLE_SEGMENT|9866,9871|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9866,9871|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9876,9884|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9876,9884|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9885,9889|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9885,9889|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9885,9889|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9885,9889|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9891,9899|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|SIMPLE_SEGMENT|9891,9899|false|false|false|||medicine
Event|Event|SIMPLE_SEGMENT|9904,9909|false|false|false|||cause
Event|Event|SIMPLE_SEGMENT|9910,9922|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9910,9922|false|false|false|C0009806|Constipation|constipation
Event|Event|SIMPLE_SEGMENT|9937,9946|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|9947,9953|false|false|false|||taking
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9958,9974|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9967,9974|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|SIMPLE_SEGMENT|9967,9974|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|SIMPLE_SEGMENT|9975,9980|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|9975,9989|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9975,9989|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|SIMPLE_SEGMENT|9981,9989|false|false|false|||softener
Drug|Organic Chemical|SIMPLE_SEGMENT|9999,10007|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9999,10007|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|10009,10015|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10009,10015|false|false|false|C0282139|Colace|Colace
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10031,10039|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10031,10039|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10040,10044|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10040,10044|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10040,10044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10040,10044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10045,10055|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|10045,10055|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10045,10055|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|10065,10073|true|false|false|||directed
Event|Event|SIMPLE_SEGMENT|10082,10088|true|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|10082,10088|true|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|10097,10101|true|false|false|||take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10107,10124|true|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10125,10134|true|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|SIMPLE_SEGMENT|10125,10134|true|false|false|||medicines
Drug|Organic Chemical|SIMPLE_SEGMENT|10143,10149|true|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10143,10149|true|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|SIMPLE_SEGMENT|10151,10158|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10151,10158|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|10151,10158|false|false|false|||Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|10160,10165|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10160,10165|false|false|false|C0593507|Advil|Advil
Event|Event|SIMPLE_SEGMENT|10160,10165|false|false|false|||Advil
Finding|Gene or Genome|SIMPLE_SEGMENT|10160,10165|false|false|false|C1422473|AVIL gene|Advil
Drug|Organic Chemical|SIMPLE_SEGMENT|10172,10181|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10172,10181|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Idea or Concept|SIMPLE_SEGMENT|10182,10185|false|false|false|C1548556|Etc.|etc
Event|Event|SIMPLE_SEGMENT|10208,10212|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|10213,10217|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10213,10217|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10213,10217|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10213,10217|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|10221,10228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10221,10228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10229,10239|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|10229,10239|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10229,10239|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|10246,10250|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|10246,10250|false|false|false|C4724437|SURE Test|sure
Event|Event|SIMPLE_SEGMENT|10260,10266|false|false|false|||taking
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10269,10279|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|10269,10279|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10269,10279|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|10283,10290|false|false|false|||protect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10296,10303|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10296,10303|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10296,10303|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|10296,10303|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|10296,10303|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10296,10303|false|false|false|C0872393|Procedure on stomach|stomach
Drug|Organic Chemical|SIMPLE_SEGMENT|10305,10313|false|false|false|C0700777|Prilosec|Prilosec
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10305,10313|false|false|false|C0700777|Prilosec|Prilosec
Drug|Organic Chemical|SIMPLE_SEGMENT|10316,10324|false|false|false|C0876139|Protonix|Protonix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10316,10324|false|false|false|C0876139|Protonix|Protonix
Drug|Organic Chemical|SIMPLE_SEGMENT|10329,10335|false|false|false|C0678119|Pepcid|Pepcid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10329,10335|false|false|false|C0678119|Pepcid|Pepcid
Event|Event|SIMPLE_SEGMENT|10329,10335|false|false|false|||Pepcid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10347,10358|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10347,10358|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10347,10358|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10347,10358|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|10363,10368|false|false|false|||cause
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10369,10376|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10369,10376|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10369,10376|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|10369,10376|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|10369,10376|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10369,10376|false|false|false|C0872393|Procedure on stomach|stomach
Event|Event|SIMPLE_SEGMENT|10378,10388|false|false|false|||irritation
Finding|Intellectual Product|SIMPLE_SEGMENT|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|SIMPLE_SEGMENT|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|SIMPLE_SEGMENT|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10378,10388|false|false|false|C0441723|Irritation|irritation
Finding|Functional Concept|SIMPLE_SEGMENT|10391,10395|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|SIMPLE_SEGMENT|10391,10395|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|SIMPLE_SEGMENT|10396,10400|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|10396,10400|false|false|false|C4724437|SURE Test|sure
Event|Event|SIMPLE_SEGMENT|10404,10408|false|false|false|||take
Drug|Organic Chemical|SIMPLE_SEGMENT|10414,10421|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10414,10421|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10422,10432|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|10422,10432|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10422,10432|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|10439,10444|false|false|false|||meals
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10439,10444|false|false|false|C1998602|Meal (occasion for eating)|meals
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10451,10456|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10451,10456|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|SIMPLE_SEGMENT|10451,10456|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10451,10456|false|false|false|C0025611|methamphetamine|glass
Event|Event|SIMPLE_SEGMENT|10451,10456|false|false|false|||glass
Drug|Food|SIMPLE_SEGMENT|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Immunologic Factor|SIMPLE_SEGMENT|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Substance|SIMPLE_SEGMENT|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Event|Event|SIMPLE_SEGMENT|10460,10464|false|false|false|||milk
Finding|Body Substance|SIMPLE_SEGMENT|10460,10464|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Finding|Intellectual Product|SIMPLE_SEGMENT|10460,10464|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Event|Event|SIMPLE_SEGMENT|10467,10468|false|false|false|||
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10468,10477|false|false|false|C1382187|Clearance of substance|Clearance
Event|Event|SIMPLE_SEGMENT|10468,10477|false|false|false|||Clearance
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10468,10477|false|false|false|C2825073|Clearance [PK]|Clearance
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10468,10477|false|false|false|C4554548|Clearance procedure|Clearance
Event|Event|SIMPLE_SEGMENT|10481,10486|false|false|false|||drive
Event|Event|SIMPLE_SEGMENT|10491,10497|false|false|false|||return
Event|Occupational Activity|SIMPLE_SEGMENT|10501,10505|false|false|false|C0043227|Work|work
Event|Event|SIMPLE_SEGMENT|10514,10523|false|false|false|||addressed
Event|Event|SIMPLE_SEGMENT|10548,10554|false|false|false|||office
Finding|Idea or Concept|SIMPLE_SEGMENT|10548,10554|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|SIMPLE_SEGMENT|10548,10560|false|false|false|C0028900|Office Visits|office visit
Event|Event|SIMPLE_SEGMENT|10555,10560|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|10555,10560|false|false|false|C0545082|Visit|visit
Event|Event|SIMPLE_SEGMENT|10563,10567|false|false|false|||Make
Finding|Functional Concept|SIMPLE_SEGMENT|10563,10567|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|SIMPLE_SEGMENT|10563,10567|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|SIMPLE_SEGMENT|10568,10572|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|10568,10572|false|false|false|C4724437|SURE Test|sure
Event|Event|SIMPLE_SEGMENT|10576,10584|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|10576,10584|false|false|false|C0549178|Continuous|continue
Event|Event|SIMPLE_SEGMENT|10588,10591|false|false|false|||use
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10597,10617|false|false|false|C0454512|Incentive spirometry|incentive spirometer
Finding|Finding|SIMPLE_SEGMENT|10625,10632|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|10628,10632|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10628,10632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10628,10632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10628,10632|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|10634,10638|false|false|false|||CALL
Finding|Functional Concept|SIMPLE_SEGMENT|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Gene or Genome|SIMPLE_SEGMENT|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Intellectual Product|SIMPLE_SEGMENT|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Mental Process|SIMPLE_SEGMENT|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10644,10651|false|false|false|C5444295||SURGEON
Event|Event|SIMPLE_SEGMENT|10644,10651|false|false|false|||SURGEON
Event|Event|SIMPLE_SEGMENT|10671,10681|true|false|false|||EXPERIENCE
Finding|Mental Process|SIMPLE_SEGMENT|10671,10681|true|false|false|C0237607;C0596545|Experience;Experience (Practice)|EXPERIENCE
Event|Event|SIMPLE_SEGMENT|10682,10685|false|false|false|||ANY
Finding|Finding|SIMPLE_SEGMENT|10706,10709|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|10706,10709|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|SIMPLE_SEGMENT|10706,10715|false|false|false|C0746890|new onset|New onset
Event|Event|SIMPLE_SEGMENT|10710,10715|false|false|false|||onset
Event|Event|SIMPLE_SEGMENT|10719,10726|false|false|false|||tremors
Finding|Sign or Symptom|SIMPLE_SEGMENT|10719,10726|false|false|false|C0040822|Tremor|tremors
Event|Event|SIMPLE_SEGMENT|10730,10738|false|false|false|||seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|10730,10738|false|false|false|C0036572|Seizures|seizures
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10745,10754|true|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|10745,10754|true|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|10745,10754|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|10758,10764|true|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|10758,10764|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10758,10764|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|10758,10767|true|false|false|C0392747|Changing|change in
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10758,10781|true|false|false|C5774124||change in mental status
Finding|Finding|SIMPLE_SEGMENT|10758,10781|true|false|false|C0856054|Mental status changes|change in mental status
Finding|Mental Process|SIMPLE_SEGMENT|10768,10774|true|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10768,10781|true|false|false|C0488568;C0488569||mental status
Finding|Finding|SIMPLE_SEGMENT|10768,10781|true|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10775,10781|true|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|10775,10781|true|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|10775,10781|true|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|10789,10797|true|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|10789,10797|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10789,10797|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10799,10807|true|false|false|C0030554|Paresthesia|tingling
Event|Event|SIMPLE_SEGMENT|10799,10807|true|false|false|||tingling
Finding|Sign or Symptom|SIMPLE_SEGMENT|10799,10807|true|false|false|C2242996|Has tingling sensation|tingling
Event|Event|SIMPLE_SEGMENT|10809,10817|true|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10809,10817|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10826,10837|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10840,10844|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|10840,10844|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|10840,10844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10840,10844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|SIMPLE_SEGMENT|10848,10856|true|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|10848,10856|true|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|10877,10887|true|false|false|||increasing
Event|Event|SIMPLE_SEGMENT|10897,10905|true|false|false|||relieved
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10909,10913|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10909,10913|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10909,10913|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10914,10924|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|10914,10924|true|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10914,10924|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|SIMPLE_SEGMENT|10927,10932|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|10927,10932|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Event|Event|SIMPLE_SEGMENT|10949,10954|false|false|false|||equal
Finding|Intellectual Product|SIMPLE_SEGMENT|10949,10954|false|false|false|C1549782|Relational Operator - Equal|equal
Procedure|Health Care Activity|SIMPLE_SEGMENT|10969,10977|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10978,10990|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10978,10990|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10978,10990|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

