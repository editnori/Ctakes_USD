CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Structure of left hand|Anatomy|false|false||Left handnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Numbness of face|Finding|false|false||face numbnessnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|left hand weakness|Finding|false|false||left hand weaknessnull|Structure of left hand|Anatomy|false|false||left handnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Weakness of hand|Finding|false|false||hand weaknessnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Clumsiness|Finding|false|false||clumsinessnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Headache|Finding|false|false||headachenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Parietal|Modifier|false|false||parietalnull|Craniotomy|Procedure|false|false||craniotomynull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Incision and drainage|Procedure|false|false||incision and drainagenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Headache|Finding|false|false||headachesnull|Structure of left hand|Anatomy|false|false||left handnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Clumsiness|Finding|false|false||clumsinessnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Headache|Finding|false|false||headachesnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Much|Finding|false|false||muchnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Clumsiness|Finding|false|false||clumsinessnull|Difficult (qualifier value)|Finding|false|false||difficulty withnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|grasp|Finding|false|false||graspingnull|Physical object|Entity|false|false||objectsnull|Fingers|Anatomy|false|false||fingersnull|Fingers, unit of measurement|LabModifier|false|false||fingersnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Once - dosing instruction fragment|Finding|false|false||Oncenull|Once (schedule frequency)|Time|false|false||Oncenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Neurology speciality|Title|false|false||neurologynull|MRI of head|Procedure|false|false||MRI headnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|MRI of head|Procedure|false|false||MRI headnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Parietal|Modifier|false|false||parietalnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||metastatic diseasenull|Metastatic Lesion|Finding|false|false||metastatic diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Disease|Disorder|false|false||diseasenull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Neurosurgical Procedures|Procedure|false|false||Neurosurgerynull|Science of neurosurgery|Title|false|false||Neurosurgerynull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Headache|Finding|false|false||headachenull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Left side of face|Anatomy|false|false||left side of facenull|LEFT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE LEFT SIDE OF THE BODY)|Modifier|false|false||left side
null|Left|Modifier|false|false||left sidenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Side of face|Anatomy|false|false||side of facenull|Side|Modifier|false|false||sidenull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Structure of left hand|Anatomy|false|false||left handnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Recent|Time|false|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Airway Resistance Test|Procedure|true|false||rawnull|Raw|Modifier|false|false||rawnull|Meat|Drug|false|false||meatsnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Dysarthria|Disorder|false|false||dysarthrianull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Chills|Finding|true|false||chillsnull|Multiple Sclerosis|Disorder|false|false||Multiple sclerosisnull|Numerous|LabModifier|false|false||Multiplenull|Sclerosis|Finding|false|false||sclerosisnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Pancreatic carcinoma|Disorder|false|false||pancreatic cancer
null|Malignant neoplasm of pancreas|Disorder|false|false||pancreatic cancernull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false||pancreaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Brother - courtesy title|Finding|false|false||brother
null|Relationship - Brother|Finding|false|false||brothernull|Brothers|Subject|false|false||brothernull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|true||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|true||cancernull|Sister|Subject|false|false||sistersnull|Malignant neoplasm of brain|Disorder|false|false||brain cancer
null|Brain Neoplasms|Disorder|false|false||brain cancernull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Mental Recall|Finding|false|false||Recallnull|Recall (activity)|Event|false|false||Recallnull|Physical object|Entity|false|false||objectsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|false|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|examination of extraocular movements|Procedure|false|false||Extraocular movementsnull|Extraocular|Finding|false|false||Extraocularnull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Nystagmus|Disorder|false|false||nystagmusnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Palate|Anatomy|false|false||Palatalnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|false|false||Tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false||Tonguenull|Procedure on tongue|Procedure|false|false||Tonguenull|Tongue|Anatomy|false|false||Tonguenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Muscular fasciculation|Finding|true|false||fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Dyskinetic syndrome|Disorder|true|false||abnormal movementsnull|Abnormal movement|Finding|true|false||abnormal movementsnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|true|false||movementsnull|Tremor|Finding|false|false||tremorsnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Power (Psychology)|Finding|false|false||powernull|Power|LabModifier|false|false||powernull|Pronator drift|Finding|true|false||pronator driftnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Craniotomy|Procedure|false|false||craniotomynull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Mental Recall|Finding|false|false||Recallnull|Recall (activity)|Event|false|false||Recallnull|Physical object|Entity|false|false||objectsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|false|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|examination of extraocular movements|Procedure|false|false||Extraocular movementsnull|Extraocular|Finding|false|false||Extraocularnull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Nystagmus|Disorder|false|false||nystagmusnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Palate|Anatomy|false|false||Palatalnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|false|false||Tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false||Tonguenull|Procedure on tongue|Procedure|false|false||Tonguenull|Tongue|Anatomy|false|false||Tonguenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Muscular fasciculation|Finding|true|false||fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Observation Interpretation - Abnormal|Finding|true|false||abnormal
null|Abnormal|Finding|true|false||abnormalnull|Movement|Finding|false|false||movementsnull|Tremor|Finding|false|false||tremorsnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Power (Psychology)|Finding|false|false||powernull|Power|LabModifier|false|false||powernull|Pronator drift|Finding|true|false||pronator driftnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|MRI of head|Procedure|false|false||MRI HEADnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||HEADnull|Procedure on head|Procedure|false|false||HEADnull|Structure of head of caudate nucleus|Anatomy|false|false||HEAD
null|Head|Anatomy|false|false||HEADnull|Head Device|Device|false|false||HEADnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Ring Dosage Form|Drug|false|false||Ringnull|Ring device|Device|false|false||Ringnull|Annular shape|Modifier|false|false||Ringnull|Ring Dosing Unit|LabModifier|false|false||Ringnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|dinoflagellate sulcus|Anatomy|false|false||sulcus
null|Groove|Anatomy|false|false||sulcusnull|malignant neoplasm of frontal lobe|Disorder|false|false||frontal lobenull|frontal lobe|Anatomy|false|false||frontal lobenull|Coronal (qualifier value)|Modifier|false|false||frontalnull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Associated with|Modifier|false|false||associatednull|Vasogenic Edema|Finding|false|false||vasogenic edemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Document Confidentiality Status - Restricted|Finding|false|false||restricted
null|Confidentiality - restricted|Finding|false|false||restricted
null|Confidentiality code - Restricted|Finding|false|false||restricted
null|Restricted|Finding|false|false||restrictednull|Diffusion - RouteOfAdministration|Finding|false|false||diffusionnull|Diffusion|Phenomenon|false|false||diffusionnull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Completely - dosing instruction fragment|Finding|true|false||completelynull|Complete|Modifier|false|false||completelynull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Brain Neoplasms|Disorder|false|false||brain neoplasmnull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Neoplastic disease|Disorder|false|false||neoplasm
null|Neoplasms|Disorder|false|false||neoplasmnull|Numerous|LabModifier|false|false||Multiplenull|FLAIR (product)|Drug|false|false||FLAIR
null|FLAIR (product)|Drug|false|false||FLAIRnull|Fluid Attenuated Inversion Recovery|Procedure|false|false||FLAIRnull|Lesion|Finding|false|false||lesionsnull|Subcortical|Anatomy|false|false||subcorticalnull|White matter|Anatomy|false|false||white matternull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Protein Domain|Drug|false|false||regionnull|Geographic Locations|Entity|false|false||regionnull|regional|Modifier|false|false||regionnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Known|Modifier|false|false||knownnull|Multiple Sclerosis|Disorder|false|false||multiple sclerosisnull|Numerous|LabModifier|false|false||multiplenull|Sclerosis|Finding|false|false||sclerosisnull|Disease|Disorder|false|false||diseasenull|MRI of head|Procedure|false|false||MRI HEADnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||HEADnull|Procedure on head|Procedure|false|false||HEADnull|Structure of head of caudate nucleus|Anatomy|false|false||HEAD
null|Head|Anatomy|false|false||HEADnull|Head Device|Device|false|false||HEADnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|null|Finding|false|false||Unchangednull|About The Same|Modifier|false|false||Unchangednull|Ring Dosage Form|Drug|false|false||ringnull|Ring device|Device|false|false||ringnull|Annular shape|Modifier|false|false||ringnull|Ring Dosing Unit|LabModifier|false|false||ringnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Right precentral sulcus|Anatomy|false|false||right precentral sulcusnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of precentral sulcus|Anatomy|false|false||precentral sulcusnull|dinoflagellate sulcus|Anatomy|false|false||sulcus
null|Groove|Anatomy|false|false||sulcusnull|malignant neoplasm of frontal lobe|Disorder|false|false||frontal lobenull|frontal lobe|Anatomy|false|false||frontal lobenull|Coronal (qualifier value)|Modifier|false|false||frontalnull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Associated with|Modifier|false|false||associatednull|Vasogenic Edema|Finding|false|false||vasogenic edemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Differential Diagnosis|Procedure|false|false||differential diagnosisnull|null|Attribute|false|false||differential diagnosisnull|Amount type - Differential|Finding|false|false||differentialnull|Differential (qualifier value)|Modifier|false|false||differential
null|Different|Modifier|false|false||differential
null|Differential - view|Modifier|false|false||differentialnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Including (qualifier)|Finding|false|false||includesnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Computerized axial tomography of brain with radiopaque contrast|Procedure|false|false||CONTRAST HEAD CTnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|CAT scan of head|Procedure|false|false||HEAD CTnull|Problems with head|Disorder|false|false||HEADnull|Procedure on head|Procedure|false|false||HEADnull|Structure of head of caudate nucleus|Anatomy|false|false||HEAD
null|Head|Anatomy|false|false||HEADnull|Head Device|Device|false|false||HEADnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Craniotomy|Procedure|false|false||craniotomynull|density|LabModifier|false|false||densitynull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Right precentral sulcus|Anatomy|false|false||right precentral sulcusnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of precentral sulcus|Anatomy|false|false||precentral sulcusnull|dinoflagellate sulcus|Anatomy|false|false||sulcus
null|Groove|Anatomy|false|false||sulcusnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|null|Time|false|false||priornull|Different|Modifier|false|false||differencenull|Delta (difference)|LabModifier|false|false||differencenull|Techniques|Finding|false|false||techniquenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Intracranial Hemorrhage|Finding|true|false||intracranial hemorrhagenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Hemorrhage|Finding|true|false||hemorrhagenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||majornull|Major <Sympycninae>|Entity|false|false||majornull|Major|Modifier|false|false||majornull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Infarction|Finding|false|false||infarctnull|bifrontal|Modifier|false|false||Bifrontalnull|Subcortical|Anatomy|false|false||subcorticalnull|White matter|Anatomy|false|false||white matternull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|Multiple Sclerosis|Disorder|false|false||multiple sclerosisnull|Numerous|LabModifier|false|false||multiplenull|Sclerosis|Finding|false|false||sclerosisnull|Recombinant Colony-Stimulating Factors|Drug|false|false||CSF
null|Colony-Stimulating Factors|Drug|false|false||CSF
null|Colony-Stimulating Factors|Drug|false|false||CSF
null|CSF2 protein, human|Drug|false|false||CSF
null|CSF2 protein, human|Drug|false|false||CSF
null|Recombinant Colony-Stimulating Factors|Drug|false|false||CSF
null|Recombinant Colony-Stimulating Factors|Drug|false|false||CSFnull|Isolated femoral agenesis/hypoplasia|Disorder|false|false||CSFnull|In Cerebrospinal Fluid|Finding|false|false||CSF
null|LAMC2 wt Allele|Finding|false|false||CSF
null|Cerebrospinal Fluid|Finding|false|false||CSFnull|Circumferential Supracrestal Fiberotomy|Procedure|false|false||CSFnull|Cerebrospinal Fluid|Finding|false|false||SPINAL FLUIDnull|Spinal|Modifier|false|false||SPINALnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Unspecified tube|Finding|false|false||TUBE
null|TUBE1 gene|Finding|false|false||TUBEnull|biomedical tube device|Device|false|false||TUBE
null|Packaging Tube|Device|false|false||TUBEnull|tube|Modifier|false|false||TUBEnull|Tube (unit of presentation)|LabModifier|false|false||TUBE
null|Tube Dosing Unit|LabModifier|false|false||TUBEnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|granulocyte|Anatomy|false|false||POLYMORPHONUCLEAR LEUKOCYTES
null|neutrophil|Anatomy|false|false||POLYMORPHONUCLEAR LEUKOCYTESnull|Specimen Type - Leukocytes|Finding|true|false||LEUKOCYTES
null|null|Finding|true|false||LEUKOCYTESnull|Leukocytes|Anatomy|false|false||LEUKOCYTESnull|Microorganisms seen|Finding|false|false||MICROORGANISMS SEENnull|Microorganism|Entity|true|false||MICROORGANISMSnull|Smearing technique|Finding|false|false||smearnull|Smear test|Procedure|false|false||smearnull|Smear - instruction imperative|Event|false|false||smearnull|Method, LOINC Axis 6|Finding|false|false||method
null|Techniques|Finding|false|false||method
null|Methods|Finding|false|false||methodnull|Diagnostic Service Section ID - Hematology|Finding|false|false||hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||hematology
null|Hematology procedure|Procedure|false|false||hematology
null|Hematologic Tests|Procedure|false|false||hematologynull|hematology (field)|Title|false|false||hematologynull|Quantitative (qualifier value)|LabModifier|false|false||quantitativenull|White Blood Cell Count procedure|Procedure|false|false||white blood cell countnull|null|Lab|false|false||white blood cell countnull|Leukocytes|Anatomy|false|false||white blood cellnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Blood Cell Count|Procedure|false|false||blood cell count
null|Complete Blood Count|Procedure|false|false||blood cell countnull|Blood Cells|Anatomy|false|false||blood cellnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Cell Count|Procedure|false|false||cell countnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Accident and Emergency department|Device|false|false||Emergency Departmentnull|interventional services emergency department|Entity|false|false||Emergency Department
null|Accident and Emergency department|Entity|false|false||Emergency Departmentnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Department - No suggested values defined|Finding|false|false||Department
null|Organization Unit Type - Department|Finding|false|false||Department
null|Department - Charge type|Finding|false|false||Departmentnull|Department|Entity|false|false||Departmentnull|Patient location type - Department|Modifier|false|false||Department
null|Department - Person location type|Modifier|false|false||Departmentnull|Left sided|Modifier|false|false||left-sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|Clumsiness|Finding|false|false||clumsinessnull|Initially|Time|false|false||initiallynull|Flare|Finding|false|false||flare
null|Exacerbation of cGVHD|Finding|false|false||flarenull|Neurology speciality|Title|false|false||Neurologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Recommendation|Finding|false|false||recommendationnull|Nuclear magnetic resonance imaging brain|Procedure|false|false||MRI brainnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||metastatic diseasenull|Metastatic Lesion|Finding|false|false||metastatic diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Disease|Disorder|false|false||diseasenull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Neurosurgical Procedures|Procedure|false|false||Neurosurgerynull|Science of neurosurgery|Title|false|false||Neurosurgerynull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Craniotomy|Procedure|false|false||craniotomynull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Irrigation Route of Administration|Finding|false|false||irrigation
null|Irrigation [MoA]|Finding|false|false||irrigationnull|Irrigation|Procedure|false|false||irrigationnull|Brain Abscess|Disorder|false|false||brain abscess
null|Cerebral abscess|Disorder|false|false||brain abscessnull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Recovering from|Modifier|false|false||recovernull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Inventory of Callous-Unemotional Traits|Finding|false|false||ICUnull|Structure of intraculminate fissure|Anatomy|false|false||ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||Meropenem
null|meropenem|Drug|false|false||Meropenem
null|meropenem|Drug|false|false||Meropenemnull|Gram's stain|Drug|false|false||Gram stain
null|Gram's stain|Drug|false|false||Gram stainnull|Bacterial stain, routine|Procedure|false|false||Gram stainnull|gram|LabModifier|false|false||Gramnull|Stains|Drug|false|false||stainnull|Staining method|Procedure|false|false||stainnull|Gram-negative bacillus|Entity|false|false||gram negative rodsnull|gram|LabModifier|false|false||gramnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Rod Photoreceptors|Anatomy|false|false||rodsnull|Gram-Positive Cocci|Entity|false|false||gram positive coccinull|gram|LabModifier|false|false||gramnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Cocci bacteria|Entity|false|false||coccinull|Chain device|Device|false|false||chainsnull|post operative (finding)|Finding|false|false||Post operativenull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Operative|Time|false|false||operativenull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|post operative (finding)|Finding|false|false||post operativenull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Operative|Time|false|false||operativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|post operative (finding)|Finding|false|false||post operativenull|Operative|Time|false|false||operativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Left upper arm structure|Anatomy|false|false||left arm
null|Left arm|Anatomy|false|false||left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Extremity Paresis|Finding|false|false||arm weaknessnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||Meropenem
null|meropenem|Drug|false|false||Meropenem
null|meropenem|Drug|false|false||Meropenemnull|Leukocytes|Anatomy|false|false||WBCnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Left upper arm structure|Anatomy|false|false||Left arm
null|Left arm|Anatomy|false|false||Left armnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper Extremity Paresis|Finding|false|false||arm weaknessnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Lethargy|Finding|false|false||lethargynull|Structure of left lower leg|Anatomy|false|false||left leg
null|Left lower extremity|Anatomy|false|false||left legnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Muscle Weakness Lower Limb|Finding|false|false||leg weakness
null|Monoparesis of lower limb|Finding|false|false||leg weaknessnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Drowsiness|Finding|false|false||sleepynull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Right sided|Modifier|false|false||right sided
null|Right|Modifier|false|false||right sidednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Extremity|Anatomy|false|false||upper extremitynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Limb structure|Anatomy|false|false||extremitynull|Left lower extremity|Anatomy|false|false||left lower extremitynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Full|Modifier|false|false||fullnull|STAT protein|Drug|false|false||stat
null|STAT protein|Drug|false|false||statnull|Extended Priority Codes - Stat|Finding|false|false||stat
null|Report priority - Stat|Finding|false|false||stat
null|SOAT1 gene|Finding|false|false||stat
null|STAT family gene|Finding|false|false||stat
null|Referral priority - STAT|Finding|false|false||statnull|Stat (do immediately)|Time|false|false||statnull|National Center for Health Care Technology, U.S.|Entity|false|false||NCHCTnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Consent (record artifact)|Finding|false|false||consent
null|ActClass - consent|Finding|false|false||consent
null|Consent|Finding|false|false||consentnull|null|Attribute|false|false||consentnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||picc line placementnull|Peripherally inserted central catheter (physical object)|Device|false|false||picc linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||piccnull|Peripherally inserted central catheter (physical object)|Device|false|false||piccnull|Vascular Access Device Placement|Procedure|false|false||line placementnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Peripherally inserted central catheter (physical object)|Device|false|false||picc linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||piccnull|Peripherally inserted central catheter (physical object)|Device|false|false||piccnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Nurses|Subject|false|false||nursenull|vancomycin|Drug|false|false||vanco
null|vancomycin|Drug|false|false||vanconull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Specimen Type - Abscess|Finding|false|false||abcessnull|culture result|Lab|false|false||culture resultnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|Still|Disorder|false|false||stillnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Gait, Unsteady|Finding|false|false||unsteady gaitnull|Unsteady|Modifier|false|false||unsteadynull|Gait|Finding|false|false||gaitnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|re-evaluation|Procedure|false|false||re-evaluationnull|Stair (equipment)|Device|false|false||stairnull|Staircase|Entity|false|false||stairnull|Diagnosis Type - Final|Finding|false|false||finalnull|Final|Time|false|false||finalnull|End-stage|Modifier|false|false||finalnull|Specimen Type - Abscess|Finding|false|false||abcessnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Streptococcus milleri|Entity|false|false||streptococcus Millerinull|Streptococcus|Entity|false|false||streptococcusnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Recommendation|Finding|false|false||recommendationsnull|vancomycin|Drug|false|false||Vanco
null|vancomycin|Drug|false|false||Vanconull|ceftriaxone|Drug|false|false||Ceftriaxone
null|ceftriaxone|Drug|false|false||Ceftriaxonenull|gram|LabModifier|false|false||gramsnull|Flagyl|Drug|false|false||Flagyl
null|Flagyl|Drug|false|false||Flagylnull|three times a day at institution-specified times|Time|false|false||Tid
null|Three times daily|Time|false|false||Tidnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Headache|Finding|false|false||headachenull|CAT scan of head|Procedure|false|false||head CTnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Postoperative Period|Time|false|false||post-operativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Home visit (procedure)|Procedure|false|false||Home servicesnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|ceftriaxone|Drug|false|false||CeftriaXONE
null|ceftriaxone|Drug|false|false||CeftriaXONEnull|Every twelve hours|Time|false|false||Q12Hnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|gram|LabModifier|false|false||gramnull|Hour|Time|false|false||hoursnull|Vial device|Device|false|false||Vialnull|Vial (unit of presentation)|LabModifier|false|false||Vial
null|Vial Dosing Unit|LabModifier|false|false||Vialnull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|levetiracetam|Drug|false|false||LeVETiracetam
null|levetiracetam|Drug|false|false||LeVETiracetamnull|Measurement of levetiracetam|Procedure|false|false||LeVETiracetamnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|levetiracetam|Drug|false|false||levetiracetam
null|levetiracetam|Drug|false|false||levetiracetamnull|Measurement of levetiracetam|Procedure|false|false||levetiracetamnull|Keppra|Drug|false|false||Keppra
null|Keppra|Drug|false|false||Keppranull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|metronidazole|Drug|true|false||MetRONIDAZOLE
null|metronidazole|Drug|true|false||MetRONIDAZOLEnull|Flagyl|Drug|false|false||FLagyl
null|Flagyl|Drug|false|false||FLagylnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|metronidazole|Drug|false|false||metronidazole
null|metronidazole|Drug|false|false||metronidazolenull|Flagyl|Drug|false|false||Flagyl
null|Flagyl|Drug|false|false||Flagylnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Oxecta|Drug|false|false||Oxecta
null|Oxecta|Drug|false|false||Oxectanull|TABLET, ORAL ONLY|Drug|false|false||tablet, oral onlynull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|heparin flush|Drug|false|false||Heparin Flush
null|heparin flush|Drug|false|false||Heparin Flushnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Flush - RouteOfAdministration|Finding|false|false||Flush
null|Flushing|Finding|false|false||Flushnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|per milliliter|LabModifier|false|false||/mlnull|Mucolipidosis Type IV|Disorder|false|false||mL IVnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|null|Attribute|false|false||line flushnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Flush - RouteOfAdministration|Finding|false|false||flush
null|Flushing|Finding|false|false||flushnull|Heparin Lock Flush|Drug|false|false||heparin lock flush
null|Heparin Lock Flush|Drug|false|false||heparin lock flushnull|Heparin lock (physical object)|Device|false|false||heparin lock
null|Vascular Access Ports|Device|false|false||heparin locknull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Lock - Remote control command|Finding|false|false||locknull|Lock Device|Device|false|false||locknull|Flush - RouteOfAdministration|Finding|false|false||flush
null|Flushing|Finding|false|false||flushnull|Porcine prosthetic valve|Finding|false|false||porcinenull|Porcine species|Entity|false|false||porcine
null|Family suidae|Entity|false|false||porcinenull|Heparin Lock Flush|Drug|false|false||heparin lock flush
null|Heparin Lock Flush|Drug|false|false||heparin lock flushnull|Heparin lock (physical object)|Device|false|false||heparin lock
null|Vascular Access Ports|Device|false|false||heparin locknull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Lock - Remote control command|Finding|false|false||locknull|Lock Device|Device|false|false||locknull|Flush - RouteOfAdministration|Finding|false|false||flush
null|Flushing|Finding|false|false||flushnull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Mucolipidosis Type IV|Disorder|false|false||ml IVnull|Hour|Time|false|false||hoursnull|Vial device|Device|false|false||Vialnull|Vial (unit of presentation)|LabModifier|false|false||Vial
null|Vial Dosing Unit|LabModifier|false|false||Vialnull|refill|Finding|false|false||Refillsnull|sodium chloride|Drug|false|false||Sodium Chloridenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|Flush - RouteOfAdministration|Finding|false|false||Flush
null|Flushing|Finding|false|false||Flushnull|Mucolipidosis Type IV|Disorder|false|false||mL IVnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|null|Attribute|false|false||line flushnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Flush - RouteOfAdministration|Finding|false|false||flush
null|Flushing|Finding|false|false||flushnull|Flush - RouteOfAdministration|Finding|false|false||Flush
null|Flushing|Finding|false|false||Flushnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|sodium chloride|Drug|false|false||sodium chloridenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|chloride ion|Drug|false|false||chloride
null|Chlorides|Drug|false|false||chloridenull|Chloride metabolic function|Finding|false|false||chloridenull|Chloride measurement|Procedure|false|false||chloridenull|Saline Flush|Procedure|false|false||Saline Flushnull|Saline Solution|Drug|false|false||Saline
null|Saline Solution|Drug|false|false||Salinenull|Saline method|Procedure|false|false||Salinenull|Flush - RouteOfAdministration|Finding|false|false||Flush
null|Flushing|Finding|false|false||Flushnull|Mucolipidosis Type IV|Disorder|false|false||ml IVnull|Syringes|Device|false|false||Syringenull|Syringe (unit of presentation)|LabModifier|false|false||Syringe
null|Syringe Dosing Unit|LabModifier|false|false||Syringenull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Brain Abscess|Disorder|false|false||Brain abscess
null|Cerebral abscess|Disorder|false|false||Brain abscessnull|Brain Diseases|Disorder|false|false||Brainnull|Head>Brain|Anatomy|false|false||Brain
null|Brain|Anatomy|false|false||Brainnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Relationship - Friend|Finding|false|false||friendnull|friend|Subject|false|false||friendnull|Family member|Subject|false|false||family membernull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Member Organization|Subject|false|false||member
null|Role Class - member|Subject|false|false||member
null|member|Subject|false|false||membernull|Surgical wound|Disorder|false|true||incisionnull|Surgical incisions|Procedure|false|true||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Daily|Time|false|false||dailynull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Lifting|Event|true|false||liftingnull|Straining (finding)|Finding|true|false||strainingnull|Excessive (qualifier value)|Modifier|false|false||excessivenull|Decompression Sickness|Disorder|false|false||bendingnull|Bending - Changing basic body position|Finding|false|false||bending
null|Does bend|Finding|false|false||bendingnull|Bent|Modifier|false|false||bendingnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Suture Joint|Anatomy|false|false||suturesnull|Surgical sutures|Device|false|false||suturesnull|Hair Specimen Code|Finding|false|false||hair
null|Hair Specimen|Finding|false|false||hairnull|Hair|Anatomy|false|false||hairnull|Suture Joint|Anatomy|false|false||suturesnull|Surgical sutures|Device|false|false||suturesnull|Staple, Surgical|Device|false|false||staplesnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|shower cap|Device|false|false||shower capnull|Shower (physical object)|Device|false|false||showernull|capsule (pharmacologic)|Drug|false|false||capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||capnull|BRD4 wt Allele|Finding|false|false||cap
null|HACD1 gene|Finding|false|false||cap
null|SERPINB6 gene|Finding|false|false||cap
null|BRD4 gene|Finding|false|false||cap
null|CAP1 gene|Finding|false|false||cap
null|SORBS1 gene|Finding|false|false||cap
null|LNPEP gene|Finding|false|false||capnull|CAP Regimen|Procedure|false|false||cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||capnull|Cap (physical object)|Device|false|false||cap
null|Syringe Caps|Device|false|false||cap
null|Cap device|Device|false|false||capnull|College of American Pathologists|Subject|false|false||capnull|Controlled Attenuation Parameter|Modifier|false|false||capnull|Capsule Dosing Unit|LabModifier|false|false||capnull|null|Finding|false|false||covernull|Cover (physical object)|Device|false|false||cover
null|Cover Device|Device|false|false||covernull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Fiber brand of calcium polycarbophil|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false||fibernull|Tissue fiber|Anatomy|false|false||fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||over the counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Anti-Inflammatory Agents|Drug|false|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|false|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Etc.|Finding|false|false||etcnull|Keppra|Drug|false|false||Keppra
null|Keppra|Drug|false|false||Keppranull|levetiracetam|Drug|false|false||Levetiracetam
null|levetiracetam|Drug|false|false||Levetiracetamnull|Measurement of levetiracetam|Procedure|false|false||Levetiracetamnull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||blood
null|In Blood|Finding|true|false||bloodnull|Work|Event|true|false||worknull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Clearance procedure|Procedure|false|false||Clearancenull|Clearance of substance|Attribute|false|false||Clearancenull|Clearance [PK]|Phenomenon|false|false||Clearancenull|Clearance|Modifier|false|false||Clearancenull|Work|Event|false|false||worknull|Postoperative Period|Time|false|false||post-operativenull|Office Visits|Procedure|false|false||office visitnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Visit|Finding|false|false||visitnull|Make - Instruction Imperative|Finding|false|false||Make
null|Manufacturer Name|Finding|false|false||Makenull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Continuous|Finding|false|false||continuenull|Incentive spirometry|Procedure|false|false||incentive spirometernull|Incentive Spirometers (device)|Device|false|false||incentive spirometernull|Incentives|Modifier|false|false||incentivenull|Spirometer Device|Device|false|false||spirometernull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions