 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Antibiotic|Allergies|180,191|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|Allergies|180,191|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|Allergies|180,191|false|false|false|||amoxicillin
Event|Event|Allergies|194,203|false|false|false|||Attending
Finding|Functional Concept|Allergies|194,203|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|229,237|false|false|false|||Weakness
Finding|Sign or Symptom|Chief Complaint|229,237|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Event|Event|Chief Complaint|242,250|false|false|false|||lethargy
Finding|Sign or Symptom|Chief Complaint|242,250|false|false|false|C0023380|Lethargy|lethargy
Finding|Classification|Chief Complaint|254,259|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|272,290|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|281,290|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|281,290|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|281,290|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|281,290|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,290|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Body Substance|History of Present Illness|328,335|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|328,335|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|328,335|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|345,349|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|345,349|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|350,353|false|false|false|||old
Event|Event|History of Present Illness|366,373|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|366,376|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|377,384|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|377,384|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|377,384|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Location or Region|History of Present Illness|385,394|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|385,399|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|395,399|false|false|false|C2598155||pain
Event|Event|History of Present Illness|395,399|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|395,399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|395,399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|404,410|false|false|false|C0002871|Anemia|anemia
Event|Event|History of Present Illness|404,410|false|false|false|||anemia
Drug|Biologically Active Substance|History of Present Illness|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Drug|Organic Chemical|History of Present Illness|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Drug|Pharmacologic Substance|History of Present Illness|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Event|Event|History of Present Illness|432,440|false|false|false|||infusion
Finding|Functional Concept|History of Present Illness|432,440|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|432,440|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|History of Present Illness|447,458|false|false|false|||complicated
Finding|Functional Concept|History of Present Illness|462,470|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|462,470|false|false|false|C0574032|Infusion procedures|infusion
Finding|Pathologic Function|History of Present Illness|462,479|false|false|false|C2368034|Infusion reaction|infusion reaction
Event|Event|History of Present Illness|471,479|false|false|false|||reaction
Finding|Functional Concept|History of Present Illness|471,479|false|false|false|C0443286|Reaction|reaction
Event|Event|History of Present Illness|481,489|false|false|false|||mottling
Finding|Finding|History of Present Illness|481,489|false|false|false|C0302133|Mottling|mottling
Event|Event|History of Present Illness|494,507|false|false|false|||discoloration
Finding|Finding|History of Present Illness|494,507|false|false|false|C0332572|Abnormal color|discoloration
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|511,515|false|false|false|C0016504|Foot|feet
Drug|Organic Chemical|History of Present Illness|524,532|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|History of Present Illness|524,532|false|false|false|C0038317|Steroids|steroids
Event|Event|History of Present Illness|524,532|false|false|false|||steroids
Event|Event|History of Present Illness|537,545|false|false|false|||presents
Event|Event|History of Present Illness|562,570|false|false|false|||lethargy
Finding|Sign or Symptom|History of Present Illness|562,570|false|false|false|C0023380|Lethargy|lethargy
Event|Event|History of Present Illness|575,583|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|575,583|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|586,593|false|false|false|||History
Finding|Conceptual Entity|History of Present Illness|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|History of Present Illness|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|History of Present Illness|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|History of Present Illness|602,609|false|false|false|||records
Finding|Idea or Concept|History of Present Illness|602,609|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|History of Present Illness|602,609|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|History of Present Illness|622,626|true|false|false|||Aunt
Finding|Body Substance|History of Present Illness|630,637|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|630,637|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|630,637|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|645,652|true|false|false|||provide
Finding|Finding|History of Present Illness|653,657|true|false|false|C4281574|Much|much
Event|Event|History of Present Illness|658,665|true|false|false|||history
Finding|Conceptual Entity|History of Present Illness|658,665|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|658,665|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|658,665|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|700,704|true|false|false|||well
Finding|Finding|History of Present Illness|700,704|true|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|726,733|true|false|false|||illness
Finding|Sign or Symptom|History of Present Illness|726,733|true|false|false|C0221423|Illness (finding)|illness
Finding|Behavior|History of Present Illness|735,745|true|false|false|C0004927|Behavior|behavioral
Finding|Individual Behavior|History of Present Illness|735,752|true|false|false|C0542299|Behavioral change|behavioral change
Event|Event|History of Present Illness|746,752|true|false|false|||change
Finding|Functional Concept|History of Present Illness|746,752|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|746,752|true|false|false|C4319952|Change - procedure|change
Disorder|Disease or Syndrome|History of Present Illness|764,768|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|History of Present Illness|764,768|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|History of Present Illness|764,768|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|History of Present Illness|764,768|false|false|false|||cold
Finding|Organism Function|History of Present Illness|764,768|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|History of Present Illness|764,768|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|764,768|false|false|false|C0010412|Cold Therapy|cold
Event|Event|History of Present Illness|777,784|false|false|false|||getting
Event|Event|History of Present Illness|810,814|false|false|false|||well
Finding|Finding|History of Present Illness|810,814|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|830,841|false|false|false|||transfusion
Finding|Functional Concept|History of Present Illness|830,841|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|830,841|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Event|History of Present Illness|882,893|false|false|false|||accompanied
Event|Event|History of Present Illness|905,910|false|false|false|||visit
Finding|Social Behavior|History of Present Illness|905,910|false|false|false|C0545082|Visit|visit
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|924,927|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|History of Present Illness|924,927|false|false|false|C0082420|Endoglin, human|end
Event|Event|History of Present Illness|924,927|false|false|false|||end
Finding|Functional Concept|History of Present Illness|924,927|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|History of Present Illness|924,927|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Event|Event|History of Present Illness|935,943|false|false|false|||infusion
Finding|Functional Concept|History of Present Illness|935,943|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|935,943|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|History of Present Illness|949,958|false|false|false|||developed
Anatomy|Body Location or Region|History of Present Illness|973,978|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|973,978|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|973,990|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|979,990|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|History of Present Illness|1006,1012|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1006,1012|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1006,1012|false|false|false|C0027497|Nausea|nausea
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1014,1019|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|History of Present Illness|1014,1019|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|History of Present Illness|1014,1019|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Finding|History of Present Illness|1014,1026|false|false|false|C0039231|Tachycardia|heart racing
Event|Event|History of Present Illness|1020,1026|false|false|false|||racing
Finding|Intellectual Product|History of Present Illness|1020,1026|false|false|false|C1561444|Racing - Production Class Code|racing
Event|Event|History of Present Illness|1036,1040|false|false|false|||sent
Attribute|Clinical Attribute|History of Present Illness|1062,1065|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1062,1065|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|1062,1065|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|History of Present Illness|1062,1065|false|false|false|||SBP
Finding|Gene or Genome|History of Present Illness|1062,1065|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|1062,1065|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|History of Present Illness|1081,1085|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|1081,1085|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1081,1085|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|1094,1101|false|false|false|||records
Finding|Idea or Concept|History of Present Illness|1094,1101|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|History of Present Illness|1094,1101|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|History of Present Illness|1115,1124|true|false|false|||shivering
Finding|Finding|History of Present Illness|1115,1124|true|false|false|C0036973|Shivering|shivering
Event|Event|History of Present Illness|1136,1140|true|false|false|||open
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1145,1149|true|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|History of Present Illness|1145,1149|true|false|false|C5848506||eyes
Finding|Finding|History of Present Illness|1152,1159|true|false|false|C0302133|Mottling|mottled
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1160,1165|true|false|false|C0018563|Hand|hands
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1170,1174|false|false|false|C0016504|Foot|feet
Event|Event|History of Present Illness|1190,1197|true|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1190,1197|true|false|false|C2699424|Concern|concern
Attribute|Clinical Attribute|History of Present Illness|1202,1213|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|1202,1213|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|1202,1213|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|1202,1213|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|History of Present Illness|1202,1222|true|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|History of Present Illness|1214,1222|true|false|false|||distress
Finding|Finding|History of Present Illness|1214,1222|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|History of Present Illness|1214,1222|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|History of Present Illness|1232,1237|false|false|false|||given
Drug|Organic Chemical|History of Present Illness|1247,1255|false|false|false|C0700899|Benadryl|Benadryl
Drug|Pharmacologic Substance|History of Present Illness|1247,1255|false|false|false|C0700899|Benadryl|Benadryl
Drug|Hormone|History of Present Illness|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Drug|Organic Chemical|History of Present Illness|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Drug|Pharmacologic Substance|History of Present Illness|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Event|Event|History of Present Illness|1267,1281|false|false|false|||hydrocortisone
Procedure|Laboratory Procedure|History of Present Illness|1267,1281|false|false|false|C0201968|Cortisol Measurement|hydrocortisone
Event|Event|History of Present Illness|1286,1294|false|false|false|||observed
Finding|Intellectual Product|History of Present Illness|1311,1315|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|1316,1326|false|false|false|||discharged
Finding|Finding|History of Present Illness|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1361,1370|false|false|false|||lethargic
Finding|Sign or Symptom|History of Present Illness|1361,1370|false|false|false|C0023380|Lethargy|lethargic
Event|Event|History of Present Illness|1372,1379|false|false|false|||meaning
Event|Event|History of Present Illness|1380,1388|false|false|false|||sleeping
Event|Event|History of Present Illness|1404,1408|true|false|false|||able
Finding|Finding|History of Present Illness|1404,1408|true|false|false|C1299581|Able (qualifier value)|able
Finding|Finding|History of Present Illness|1404,1415|true|false|false|C0560880|Able to sit|able to sit
Finding|Finding|History of Present Illness|1404,1418|true|false|false|C0560835|Able to sit up|able to sit up
Finding|Finding|History of Present Illness|1412,1415|true|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Gene or Genome|History of Present Illness|1412,1415|true|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Finding|History of Present Illness|1412,1418|true|false|false|C0560837|Does sit up|sit up
Finding|Daily or Recreational Activity|History of Present Illness|1423,1427|true|false|false|C0080331|Walking (function)|walk
Event|Activity|History of Present Illness|1436,1441|true|false|false|C5966184|Issue (action)|issue
Event|Event|History of Present Illness|1436,1441|true|false|false|||issue
Finding|Finding|History of Present Illness|1436,1441|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|History of Present Illness|1436,1441|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|History of Present Illness|1448,1455|false|false|false|||arrived
Event|Event|History of Present Illness|1456,1460|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1456,1460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1456,1460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1456,1460|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|1469,1473|false|false|false|||went
Disorder|Disease or Syndrome|History of Present Illness|1477,1480|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|History of Present Illness|1477,1480|false|false|false|||bed
Finding|Intellectual Product|History of Present Illness|1477,1480|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|History of Present Illness|1494,1496|false|false|false|||AM
Event|Event|History of Present Illness|1514,1519|false|false|false|||check
Disorder|Disease or Syndrome|History of Present Illness|1539,1544|false|false|false|C1410088|Still|still
Event|Event|History of Present Illness|1545,1553|false|false|false|||sleeping
Event|Event|History of Present Illness|1563,1572|false|false|false|||reporting
Event|Event|History of Present Illness|1575,1583|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|1575,1583|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|1595,1606|false|false|false|||transfusion
Finding|Functional Concept|History of Present Illness|1595,1606|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1595,1606|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Activity|History of Present Illness|1607,1612|false|false|false|C1882509|put - instruction imperative|place
Event|Event|History of Present Illness|1607,1612|false|false|false|||place
Finding|Functional Concept|History of Present Illness|1607,1612|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|History of Present Illness|1607,1612|false|false|false|C1533810||place
Event|Event|History of Present Illness|1613,1617|false|false|false|||said
Event|Event|History of Present Illness|1624,1630|false|false|false|||happen
Event|Event|History of Present Illness|1644,1651|true|false|false|||mention
Event|Event|History of Present Illness|1658,1672|true|false|false|||characteristic
Event|Event|History of Present Illness|1684,1688|false|false|false|||gave
Drug|Organic Chemical|History of Present Illness|1693,1706|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|History of Present Illness|1693,1706|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|History of Present Illness|1693,1706|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|History of Present Illness|1693,1706|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Inorganic Chemical|History of Present Illness|1711,1716|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|History of Present Illness|1711,1716|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|History of Present Illness|1711,1716|false|false|false|||water
Finding|Intellectual Product|History of Present Illness|1711,1716|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1711,1716|false|false|false|C0020311|Hydrotherapy|water
Event|Event|History of Present Illness|1725,1729|false|false|false|||went
Drug|Organic Chemical|History of Present Illness|1738,1743|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|History of Present Illness|1738,1743|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|History of Present Illness|1738,1743|false|false|false|||sleep
Finding|Organism Function|History of Present Illness|1738,1743|false|false|false|C0037313|Sleep|sleep
Finding|Idea or Concept|History of Present Illness|1754,1758|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|History of Present Illness|1774,1779|false|false|false|||heard
Finding|Finding|History of Present Illness|1784,1789|false|false|false|C0234422|Awake (finding)|awake
Disorder|Disease or Syndrome|History of Present Illness|1798,1803|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|1798,1803|false|false|false|||times
Event|Event|History of Present Illness|1808,1811|false|false|false|||use
Event|Event|History of Present Illness|1816,1824|false|false|false|||bathroom
Finding|Intellectual Product|History of Present Illness|1826,1830|false|false|false|C1720594|Then - dosing instruction fragment|Then
Event|Event|History of Present Illness|1837,1840|false|false|false|||got
Finding|Idea or Concept|History of Present Illness|1866,1869|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1866,1869|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|1913,1919|false|false|false|||became
Event|Event|History of Present Illness|1920,1927|false|false|false|||worried
Finding|Finding|History of Present Illness|1920,1927|false|false|false|C0233481|Worried|worried
Event|Event|History of Present Illness|1933,1937|false|false|false|||told
Event|Event|History of Present Illness|1972,1976|false|false|false|||able
Finding|Finding|History of Present Illness|1972,1976|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|1980,1982|false|false|false|||do
Event|Event|History of Present Illness|1999,2003|false|false|false|||said
Event|Event|History of Present Illness|2008,2017|false|false|false|||continued
Event|Event|History of Present Illness|2028,2036|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2028,2036|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|2041,2045|false|false|false|||felt
Event|Event|History of Present Illness|2046,2052|false|false|false|||sleepy
Finding|Finding|History of Present Illness|2046,2052|false|false|false|C0013144|Drowsiness|sleepy
Event|Event|History of Present Illness|2062,2072|false|false|false|||instructed
Event|Event|History of Present Illness|2076,2078|false|false|false|||go
Event|Event|History of Present Illness|2096,2100|false|false|false|||went
Event|Event|History of Present Illness|2122,2132|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|2122,2132|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|2122,2132|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|History of Present Illness|2213,2219|false|false|false|||drowsy
Finding|Finding|History of Present Illness|2213,2219|false|false|false|C0013144|Drowsiness|drowsy
Event|Event|History of Present Illness|2236,2241|false|false|false|||voice
Finding|Idea or Concept|History of Present Illness|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|History of Present Illness|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|History of Present Illness|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Attribute|Clinical Attribute|History of Present Illness|2244,2249|false|false|false|C5890168||alert
Drug|Organic Chemical|History of Present Illness|2244,2249|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|History of Present Illness|2244,2249|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|History of Present Illness|2244,2249|false|false|false|||alert
Finding|Finding|History of Present Illness|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|History of Present Illness|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|History of Present Illness|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Finding|History of Present Illness|2250,2258|false|false|false|C1961028|Oriented to place|oriented
Event|Event|History of Present Illness|2259,2261|false|false|false|||x3
Finding|Idea or Concept|History of Present Illness|2264,2274|false|false|false|C0332290|Consistent with|consistent
Anatomy|Body Location or Region|History of Present Illness|2275,2278|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2275,2278|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|History of Present Illness|2275,2278|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|History of Present Illness|2275,2278|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|History of Present Illness|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|History of Present Illness|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|History of Present Illness|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|History of Present Illness|2279,2289|false|false|false|||fluttering
Finding|Pathologic Function|History of Present Illness|2279,2289|false|false|false|C0016385|Cardiac Flutter|fluttering
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2291,2297|false|false|false|C0034121|Pupil|pupils
Event|Event|History of Present Illness|2298,2306|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2298,2306|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|History of Present Illness|2298,2315|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2310,2315|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|History of Present Illness|2310,2315|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|History of Present Illness|2310,2315|false|false|false|||light
Finding|Finding|History of Present Illness|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|History of Present Illness|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|History of Present Illness|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2310,2315|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2310,2315|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|History of Present Illness|2320,2331|false|false|false|C0241886|Extraocular|extraocular
Finding|Finding|History of Present Illness|2320,2345|false|false|false|C0702182|Extraocular eye movement|extraocular eye movements
Anatomy|Body Location or Region|History of Present Illness|2332,2335|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2332,2335|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|History of Present Illness|2332,2335|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|History of Present Illness|2332,2335|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|History of Present Illness|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|History of Present Illness|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|History of Present Illness|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Physiologic Function|History of Present Illness|2332,2345|false|false|false|C0015413|Eye Movements|eye movements
Event|Event|History of Present Illness|2336,2345|false|false|false|||movements
Finding|Organism Function|History of Present Illness|2336,2345|false|false|false|C0026649|Movement|movements
Event|Event|History of Present Illness|2346,2350|false|false|false|||full
Event|Event|History of Present Illness|2380,2384|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|2380,2384|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|2380,2384|false|false|false|C0582103|Medical Examination|exam
Finding|Gene or Genome|History of Present Illness|2387,2390|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|History of Present Illness|2387,2390|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|History of Present Illness|2391,2395|false|false|false|||work
Event|Occupational Activity|History of Present Illness|2391,2395|false|false|false|C0043227|Work|work
Anatomy|Cell|History of Present Illness|2408,2411|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2417,2420|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|2417,2420|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|History of Present Illness|2417,2420|false|false|false|||Hgb
Finding|Gene or Genome|History of Present Illness|2417,2420|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|2417,2420|false|false|false|C0019029|Hemoglobin concentration|Hgb
Drug|Organic Chemical|History of Present Illness|2435,2441|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|History of Present Illness|2435,2441|false|false|false|C0074722|sodium bicarbonate|bicarb
Event|Event|History of Present Illness|2435,2441|false|false|false|||bicarb
Event|Event|History of Present Illness|2469,2473|false|false|false|||LFTs
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Drug|Biologically Active Substance|History of Present Illness|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Drug|Pharmacologic Substance|History of Present Illness|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Event|Event|History of Present Illness|2483,2491|false|false|false|||Ferritin
Procedure|Laboratory Procedure|History of Present Illness|2483,2491|false|false|false|C0373607|Ferritin measurement|Ferritin
Event|Event|History of Present Illness|2501,2503|false|false|false|||pH
Lab|Laboratory or Test Result|History of Present Illness|2514,2518|false|false|false|C0391839|Carbon dioxide, partial pressure|PCO2
Procedure|Laboratory Procedure|History of Present Illness|2514,2518|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|PCO2
Anatomy|Cell|History of Present Illness|2559,2562|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|History of Present Illness|2571,2580|true|false|false|C0026473|Monocytes|monocytes
Drug|Biologically Active Substance|History of Present Illness|2581,2588|true|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|History of Present Illness|2581,2588|true|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|History of Present Illness|2581,2588|true|false|false|C0017725|glucose|glucose
Event|Event|History of Present Illness|2581,2588|true|false|false|||glucose
Lab|Laboratory or Test Result|History of Present Illness|2581,2588|true|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|History of Present Illness|2581,2588|true|false|false|C0337438|Glucose measurement|glucose
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2593,2600|true|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|History of Present Illness|2593,2600|true|false|false|C0033684|Proteins|protein
Event|Event|History of Present Illness|2593,2600|true|false|false|||protein
Finding|Conceptual Entity|History of Present Illness|2593,2600|true|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|History of Present Illness|2593,2600|true|false|false|C0202202|Protein measurement|protein
Event|Event|History of Present Illness|2608,2621|true|false|false|||xanthochromia
Finding|Finding|History of Present Illness|2608,2621|true|false|false|C0863146|Yellow color (finding)|xanthochromia
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|History of Present Illness|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|History of Present Illness|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Event|Event|History of Present Illness|2642,2645|false|false|false|||MRA
Lab|Laboratory or Test Result|History of Present Illness|2642,2645|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|History of Present Illness|2642,2645|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Drug|Immunologic Factor|History of Present Illness|2650,2653|false|false|false|C0876081|MRV|MRV
Drug|Pharmacologic Substance|History of Present Illness|2650,2653|false|false|false|C0876081|MRV|MRV
Event|Event|History of Present Illness|2650,2653|false|false|false|||MRV
Event|Event|History of Present Illness|2660,2666|true|false|false|||showed
Event|Event|History of Present Illness|2670,2678|true|false|false|||thrombus
Finding|Pathologic Function|History of Present Illness|2670,2678|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|History of Present Illness|2682,2689|true|false|false|||venoous
Event|Event|History of Present Illness|2690,2700|true|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|2690,2700|true|false|false|C0040053|Thrombosis|thrombosis
Event|Event|History of Present Illness|2710,2721|false|false|false|||transferred
Event|Event|History of Present Illness|2741,2751|false|false|false|||management
Event|Occupational Activity|History of Present Illness|2741,2751|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|2741,2751|false|false|false|C0376636|Disease Management|management
Event|Activity|History of Present Illness|2760,2769|false|false|false|C0021822|Interview|interview
Event|Event|History of Present Illness|2760,2769|false|false|false|||interview
Finding|Intellectual Product|History of Present Illness|2760,2769|false|false|false|C0935630|Published Interview|interview
Event|Event|History of Present Illness|2781,2788|true|false|false|||provide
Finding|Finding|History of Present Illness|2789,2793|true|true|false|C4281574|Much|much
Event|Event|History of Present Illness|2794,2801|true|false|false|||history
Finding|Conceptual Entity|History of Present Illness|2794,2801|true|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|2794,2801|true|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|2794,2801|true|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|2817,2820|false|false|false|||say
Event|Event|History of Present Illness|2846,2851|false|false|false|||tired
Finding|Finding|History of Present Illness|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|History of Present Illness|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|History of Present Illness|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|History of Present Illness|2858,2863|false|false|false|||keeps
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2868,2872|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|History of Present Illness|2868,2872|false|false|false|C5848506||eyes
Event|Event|History of Present Illness|2873,2879|false|false|false|||closed
Event|Event|History of Present Illness|2888,2899|false|false|false|||questioning
Finding|Mental Process|History of Present Illness|2888,2899|false|false|false|C0876928|Sexual Orientation - Questioning|questioning
Event|Event|History of Present Illness|2905,2912|false|false|false|||reports
Event|Event|History of Present Illness|2913,2921|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2913,2921|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|2933,2941|true|false|false|||describe
Event|Event|History of Present Illness|2958,2966|false|false|false|||features
Event|Event|History of Present Illness|2979,2990|false|false|false|||photophobia
Finding|Sign or Symptom|History of Present Illness|2979,2990|false|false|false|C0085636|Photophobia|photophobia
Event|Event|History of Present Illness|2999,3005|false|false|false|||unable
Finding|Finding|History of Present Illness|2999,3005|false|false|false|C1299582|Unable|unable
Event|Activity|History of Present Illness|3010,3021|false|false|false|C5909499|Participate|participate
Event|Event|History of Present Illness|3031,3042|false|false|false|||questioning
Finding|Mental Process|History of Present Illness|3031,3042|false|false|false|C0876928|Sexual Orientation - Questioning|questioning
Finding|Intellectual Product|History of Present Illness|3044,3049|false|false|false|C4050225|Often - answer to question|often
Event|Event|History of Present Illness|3058,3065|false|false|false|||tearful
Finding|Finding|History of Present Illness|3058,3065|false|false|false|C0424109|Weepiness|tearful
Event|Event|History of Present Illness|3070,3076|false|false|false|||saying
Event|Event|History of Present Illness|3082,3091|false|false|false|||questions
Event|Event|History of Present Illness|3096,3100|false|false|false|||hard
Event|Event|History of Present Illness|3113,3119|false|false|false|||father
Finding|Conceptual Entity|History of Present Illness|3113,3119|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|History of Present Illness|3113,3119|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|History of Present Illness|3141,3148|true|false|false|||history
Finding|Conceptual Entity|History of Present Illness|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3141,3151|true|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|3152,3160|true|false|false|||seizures
Finding|Sign or Symptom|History of Present Illness|3152,3160|true|false|false|C0036572|Seizures|seizures
Anatomy|Body System|History of Present Illness|3165,3168|true|false|false|C3714787|Central Nervous System|CNS
Disorder|Disease or Syndrome|History of Present Illness|3169,3178|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|History of Present Illness|3169,3178|false|false|false|||infection
Finding|Pathologic Function|History of Present Illness|3169,3178|false|false|false|C3714514|Infection|infection
Disorder|Injury or Poisoning|History of Present Illness|3195,3205|false|false|false|C0006107|Brain Concussion|concussion
Event|Event|History of Present Illness|3195,3205|false|false|false|||concussion
Event|Event|History of Present Illness|3219,3222|false|false|false|||old
Disorder|Disease or Syndrome|Past Medical History|3249,3255|false|false|false|C0002871|Anemia|Anemia
Event|Event|Past Medical History|3249,3255|false|false|false|||Anemia
Event|Event|Family Medical History|3295,3301|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|3295,3301|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|3309,3315|false|false|false|C0007570|Celiac Disease|celiac
Disorder|Disease or Syndrome|Family Medical History|3309,3323|false|false|false|C0007570|Celiac Disease|celiac disease
Finding|Gene or Genome|Family Medical History|3309,3323|false|false|false|C1332802|CTLA4 gene|celiac disease
Disorder|Disease or Syndrome|Family Medical History|3316,3323|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|3316,3323|false|false|false|||disease
Finding|Functional Concept|Family Medical History|3328,3338|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Finding|Pathologic Function|Family Medical History|3328,3338|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Disorder|Disease or Syndrome|Family Medical History|3328,3353|false|false|false|C0342158|Hypothyroidism, Autoimmune|autoimmune hypothyroidism
Disorder|Disease or Syndrome|Family Medical History|3339,3353|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Event|Event|Family Medical History|3339,3353|false|false|false|||hypothyroidism
Disorder|Disease or Syndrome|Family Medical History|3355,3358|false|false|false|C1262020|Diffuse alveolar damage|Dad
Event|Event|Family Medical History|3355,3358|false|false|false|||Dad
Finding|Intellectual Product|Family Medical History|3355,3358|false|false|false|C3641946|Disability Assessment for Dementia Questionnaire|Dad
Event|Event|Family Medical History|3362,3369|false|false|false|||healthy
Event|Event|Family Medical History|3381,3387|false|false|false|||cousin
Event|Event|Family Medical History|3393,3401|false|false|false|||seizures
Finding|Sign or Symptom|Family Medical History|3393,3401|false|false|false|C0036572|Seizures|seizures
Procedure|Health Care Activity|General Exam|3420,3429|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|General Exam|3430,3434|false|false|false|||exam
Finding|Functional Concept|General Exam|3430,3434|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3430,3434|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|3462,3469|false|false|false|||General
Finding|Classification|General Exam|3462,3469|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3462,3469|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|3485,3493|false|false|false|||sleeping
Anatomy|Body Location or Region|General Exam|3506,3509|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|General Exam|3506,3509|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|General Exam|3506,3509|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|General Exam|3506,3509|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|General Exam|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|General Exam|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|General Exam|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Anatomy|Body Part, Organ, or Organ Component|General Exam|3506,3513|false|false|false|C2706046|Eye lid|eye lid
Event|Event|General Exam|3514,3524|false|false|false|||fluttering
Finding|Pathologic Function|General Exam|3514,3524|false|false|false|C0016385|Cardiac Flutter|fluttering
Anatomy|Body Part, Organ, or Organ Component|General Exam|3526,3529|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|General Exam|3526,3529|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|General Exam|3526,3529|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|General Exam|3526,3529|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Event|Event|General Exam|3530,3539|false|false|false|||movements
Finding|Organism Function|General Exam|3530,3539|false|false|false|C0026649|Movement|movements
Finding|Sign or Symptom|General Exam|3552,3566|false|false|false|C0233565|Bradykinesia|slow movements
Event|Event|General Exam|3557,3566|false|false|false|||movements
Finding|Organism Function|General Exam|3557,3566|false|false|false|C0026649|Movement|movements
Anatomy|Body Location or Region|General Exam|3570,3574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|3570,3574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|General Exam|3570,3574|false|false|false|C0362076|Problems with head|head
Event|Event|General Exam|3570,3574|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|General Exam|3570,3574|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|General Exam|3593,3598|false|false|false|C1512338|HEENT|HEENT
Disorder|Injury or Poisoning|General Exam|3603,3609|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|General Exam|3603,3609|true|false|false|||trauma
Procedure|Health Care Activity|General Exam|3603,3609|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|General Exam|3614,3622|true|false|false|||jaundice
Finding|Finding|General Exam|3614,3622|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|General Exam|3614,3622|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|General Exam|3627,3634|true|false|false|||lesions
Finding|Finding|General Exam|3627,3634|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|General Exam|3638,3648|true|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|General Exam|3654,3657|false|false|false|||RRR
Event|Event|General Exam|3663,3667|false|false|false|||Pulm
Procedure|Health Care Activity|General Exam|3663,3667|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Event|Event|General Exam|3669,3678|false|false|false|||breathing
Disorder|Congenital Abnormality|General Exam|3698,3701|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|3698,3701|false|false|false|||Ext
Finding|Gene or Genome|General Exam|3698,3701|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|3703,3709|true|false|false|||clammy
Finding|Finding|General Exam|3703,3709|true|false|false|C0392162|Clammy skin|clammy
Event|Event|General Exam|3711,3715|true|false|false|||warm
Finding|Finding|General Exam|3711,3715|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3711,3715|true|false|false|C0687712|warming process|warm
Disorder|Disease or Syndrome|General Exam|3723,3727|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|3723,3727|true|false|false|||rash
Finding|Pathologic Function|General Exam|3723,3727|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|3723,3727|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Mental Process|General Exam|3743,3749|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|3743,3756|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|General Exam|3743,3756|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|General Exam|3750,3756|false|false|false|C5889824||Status
Event|Event|General Exam|3750,3756|false|false|false|||Status
Finding|Idea or Concept|General Exam|3750,3756|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|General Exam|3778,3783|false|false|false|||upset
Finding|Mental Process|General Exam|3778,3783|false|false|false|C3887804|Feeling upset|upset
Event|Event|General Exam|3791,3795|false|false|false|||exam
Finding|Functional Concept|General Exam|3791,3795|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3791,3795|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|3803,3810|false|false|false|||tearful
Finding|Finding|General Exam|3803,3810|false|false|false|C0424109|Weepiness|tearful
Disorder|Disease or Syndrome|General Exam|3814,3819|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Intellectual Product|General Exam|3821,3825|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|General Exam|3826,3832|false|false|false|||abulic
Disorder|Disease or Syndrome|General Exam|3842,3847|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|General Exam|3842,3847|false|false|false|||times
Anatomy|Body Part, Organ, or Organ Component|General Exam|3849,3853|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|General Exam|3849,3853|false|false|false|C5848506||Eyes
Disorder|Congenital Abnormality|General Exam|3849,3858|false|false|false|C0266574|Ablepharon|Eyes open
Event|Event|General Exam|3854,3858|false|false|false|||open
Event|Event|General Exam|3875,3880|false|false|false|||voice
Finding|Idea or Concept|General Exam|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Event|Event|General Exam|3889,3897|false|false|false|||oriented
Event|Event|General Exam|3913,3917|true|false|false|||full
Event|Event|General Exam|3924,3929|false|false|false|||Knows
Finding|Idea or Concept|General Exam|3943,3951|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|General Exam|3965,3969|true|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Event|Event|General Exam|3975,3979|false|false|false|||says
Finding|Idea or Concept|General Exam|3995,4003|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|General Exam|4018,4023|false|false|false|||tired
Finding|Finding|General Exam|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|General Exam|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|General Exam|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|General Exam|4033,4039|false|false|false|||unable
Finding|Finding|General Exam|4033,4039|false|false|false|C1299582|Unable|unable
Drug|Food|General Exam|4044,4051|false|false|false|C0359589|Provide (product)|provide
Event|Activity|General Exam|4044,4051|false|false|false|C1999230|Providing (action)|provide
Event|Event|General Exam|4044,4051|false|false|false|||provide
Event|Event|General Exam|4052,4059|false|false|false|||history
Finding|Conceptual Entity|General Exam|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|General Exam|4061,4067|true|false|false|||Speech
Finding|Organism Function|General Exam|4061,4067|true|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|4061,4067|true|false|false|C0846595|Speech assessment|Speech
Event|Event|General Exam|4075,4085|true|false|false|||dysarthric
Event|Event|General Exam|4087,4091|true|false|false|||says
Event|Event|General Exam|4096,4101|true|false|false|||words
Event|Event|General Exam|4107,4112|true|false|false|||asked
Event|Event|General Exam|4113,4122|true|false|false|||questions
Finding|Functional Concept|General Exam|4127,4138|true|false|false|C0205359|Spontaneous|spontaneous
Event|Event|General Exam|4139,4145|true|false|false|||speech
Finding|Organism Function|General Exam|4139,4145|true|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|General Exam|4139,4145|true|false|false|C0846595|Speech assessment|speech
Event|Event|General Exam|4146,4152|true|false|false|||output
Finding|Conceptual Entity|General Exam|4146,4152|true|false|false|C1709366|system output|output
Procedure|Health Care Activity|General Exam|4146,4152|true|false|false|C3251815|Measurement of fluid output|output
Event|Event|General Exam|4154,4161|false|false|false|||Follows
Finding|Gene or Genome|General Exam|4162,4168|false|false|false|C1424587|LITAF gene|simple
Event|Event|General Exam|4169,4177|false|false|false|||commands
Anatomy|Body Part, Organ, or Organ Component|General Exam|4188,4192|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|4188,4192|false|false|false|C5848506||eyes
Event|Activity|General Exam|4194,4198|false|false|false|C0206244|Lifting|lift
Anatomy|Body Part, Organ, or Organ Component|General Exam|4199,4203|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|General Exam|4199,4203|false|false|false|C5781420||legs
Event|Event|General Exam|4212,4216|false|false|false|||able
Finding|Finding|General Exam|4212,4216|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|General Exam|4220,4224|false|false|false|||name
Finding|Intellectual Product|General Exam|4220,4224|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Event|Event|General Exam|4226,4229|false|false|false|||key
Finding|Conceptual Entity|General Exam|4226,4229|false|false|false|C1554080;C1706198|Key - HL7UpdateMode;Key - value|key
Finding|Intellectual Product|General Exam|4226,4229|false|false|false|C1554080;C1706198|Key - HL7UpdateMode;Key - value|key
Anatomy|Body Part, Organ, or Organ Component|General Exam|4236,4243|false|false|false|C0015731;C1744713|Feathers|feather
Drug|Immunologic Factor|General Exam|4236,4243|false|false|false|C3486460|Feathers (allergen)|feather
Disorder|Disease or Syndrome|General Exam|4248,4254|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|General Exam|4248,4254|false|false|false|||stroke
Finding|Finding|General Exam|4248,4254|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|General Exam|4255,4259|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|General Exam|4255,4259|false|false|false|C0018799|Heart Diseases|card
Event|Event|General Exam|4255,4259|false|false|false|||card
Finding|Intellectual Product|General Exam|4255,4259|false|false|false|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|General Exam|4255,4259|false|false|false|C5202809|CaRD Regimen|card
Finding|Intellectual Product|General Exam|4264,4268|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|General Exam|4269,4274|false|false|false|||stops
Event|Event|General Exam|4275,4281|false|false|false|||naming
Event|Event|General Exam|4286,4292|false|false|false|||closes
Anatomy|Body Part, Organ, or Organ Component|General Exam|4297,4301|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|4297,4301|false|false|false|C5848506||eyes
Event|Event|General Exam|4307,4312|false|false|false|||reads
Event|Event|General Exam|4323,4331|false|false|false|||sentence
Finding|Intellectual Product|General Exam|4323,4331|false|false|false|C0876929|Sentence|sentence
Disorder|Disease or Syndrome|General Exam|4335,4341|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|General Exam|4335,4341|false|false|false|||stroke
Finding|Finding|General Exam|4335,4341|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|General Exam|4342,4346|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|General Exam|4342,4346|false|false|false|C0018799|Heart Diseases|card
Event|Event|General Exam|4342,4346|false|false|false|||card
Finding|Intellectual Product|General Exam|4342,4346|false|false|false|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|General Exam|4342,4346|false|false|false|C5202809|CaRD Regimen|card
Finding|Intellectual Product|General Exam|4351,4355|true|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|General Exam|4368,4374|true|false|false|||closes
Anatomy|Body Part, Organ, or Organ Component|General Exam|4379,4383|true|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|4379,4383|true|false|false|C5848506||eyes
Event|Event|General Exam|4390,4395|false|false|false|||asked
Event|Event|General Exam|4399,4407|false|false|false|||describe
Disorder|Disease or Syndrome|General Exam|4408,4414|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|General Exam|4408,4414|false|false|false|||stroke
Finding|Finding|General Exam|4408,4414|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|General Exam|4415,4419|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|General Exam|4415,4419|false|false|true|C0018799|Heart Diseases|card
Event|Event|General Exam|4415,4419|false|false|false|||card
Finding|Intellectual Product|General Exam|4415,4419|false|false|true|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|General Exam|4415,4419|false|false|true|C5202809|CaRD Regimen|card
Event|Event|General Exam|4432,4436|false|false|false|||says
Event|Event|General Exam|4461,4472|true|false|false|||participate
Event|Event|General Exam|4484,4488|true|false|false|||exam
Finding|Functional Concept|General Exam|4484,4488|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4484,4488|true|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|General Exam|4492,4499|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4492,4506|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|4492,4506|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|4500,4506|false|false|false|C0027740|Nerve|Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|4527,4533|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|4546,4550|true|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|4559,4568|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|4559,4568|true|false|false|||nystagmus
Event|Event|General Exam|4578,4591|false|false|false|||confrontation
Finding|Finding|General Exam|4578,4591|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|4578,4591|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|4578,4591|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Diagnostic Procedure|General Exam|4594,4610|true|false|false|C0029090|Ophthalmoscopy|Fundoscopic exam
Event|Event|General Exam|4606,4610|true|false|false|||exam
Finding|Functional Concept|General Exam|4606,4610|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4606,4610|true|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|4611,4619|true|false|false|||revealed
Disorder|Disease or Syndrome|General Exam|4623,4634|true|false|false|C0030353|Papilledema|papilledema
Event|Event|General Exam|4623,4634|true|false|false|||papilledema
Event|Event|General Exam|4636,4644|true|false|false|||exudates
Finding|Body Substance|General Exam|4636,4644|true|false|false|C0015388|Exudate|exudates
Event|Event|General Exam|4649,4660|true|false|false|||hemorrhages
Finding|Pathologic Function|General Exam|4649,4660|true|false|false|C0019080|Hemorrhage|hemorrhages
Anatomy|Body Part, Organ, or Organ Component|General Exam|4663,4666|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|4663,4666|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|4671,4677|true|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|General Exam|4671,4683|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|General Exam|4671,4683|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|General Exam|4678,4683|true|false|false|||droop
Anatomy|Body Location or Region|General Exam|4685,4691|true|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4692,4703|true|false|false|C1995013|Set of muscles|musculature
Event|Event|General Exam|4704,4713|true|false|false|||symmetric
Finding|Conceptual Entity|General Exam|4704,4713|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|4704,4713|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|General Exam|4720,4727|false|false|false|||grimace
Finding|Sign or Symptom|General Exam|4720,4727|false|false|false|C0239779|Grimaces|grimace
Anatomy|Body Part, Organ, or Organ Component|General Exam|4730,4734|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|4730,4734|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|4730,4734|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|General Exam|4736,4743|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|4736,4743|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|4744,4750|false|false|false|||intact
Finding|Finding|General Exam|4744,4750|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|4754,4758|false|false|false|||exam
Finding|Functional Concept|General Exam|4754,4758|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4754,4758|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|General Exam|4767,4773|false|false|false|C0700374|Palate|Palate
Event|Event|General Exam|4774,4782|false|false|false|||elevates
Anatomy|Body Part, Organ, or Organ Component|General Exam|4804,4810|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|4804,4810|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Event|Event|General Exam|4804,4810|false|false|false|||Tongue
Procedure|Health Care Activity|General Exam|4804,4810|false|false|false|C0872394|Procedure on tongue|Tongue
Event|Event|General Exam|4811,4820|false|false|false|||protrudes
Anatomy|Cell Component|General Exam|4824,4831|false|false|false|C1660780|midline cell component|midline
Finding|Functional Concept|General Exam|4835,4840|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|4849,4853|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|4849,4853|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|4849,4853|false|false|false|||bulk
Event|Event|General Exam|4855,4859|false|false|false|||tone
Event|Event|General Exam|4876,4880|false|false|false|||says
Event|Event|General Exam|4892,4896|true|false|false|||move
Anatomy|Body Part, Organ, or Organ Component|General Exam|4901,4905|true|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|4901,4905|true|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|4901,4905|true|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|General Exam|4901,4905|true|false|false|||arms
Finding|Gene or Genome|General Exam|4901,4905|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|4901,4905|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|General Exam|4912,4916|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|4912,4916|false|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|4912,4916|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|General Exam|4912,4916|false|false|false|||arms
Finding|Gene or Genome|General Exam|4912,4916|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|4912,4916|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|General Exam|4917,4923|false|false|false|||placed
Anatomy|Body Location or Region|General Exam|4933,4937|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|4933,4937|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|General Exam|4933,4937|false|false|false|C0362076|Problems with head|head
Event|Event|General Exam|4933,4937|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|General Exam|4933,4937|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|4943,4947|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|4943,4947|false|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|4943,4947|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|General Exam|4943,4947|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|4943,4947|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Location or Region|General Exam|4964,4968|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|General Exam|4964,4968|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|General Exam|4964,4968|false|false|false|||face
Finding|Gene or Genome|General Exam|4964,4968|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Drug|Biomedical or Dental Material|General Exam|4980,4985|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|General Exam|4980,4985|false|false|false|||drops
Disorder|Disease or Syndrome|General Exam|4993,4996|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|4993,4996|false|false|false|||bed
Finding|Intellectual Product|General Exam|4993,4996|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|General Exam|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Functional Concept|General Exam|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Idea or Concept|General Exam|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Event|Event|General Exam|5013,5020|false|false|false|||fashion
Event|Event|General Exam|5032,5036|false|false|false|||lift
Anatomy|Body Part, Organ, or Organ Component|General Exam|5041,5045|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|5041,5045|false|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|5041,5045|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|General Exam|5041,5045|false|false|false|||arms
Finding|Gene or Genome|General Exam|5041,5045|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|5041,5045|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|General Exam|5049,5053|false|false|false|||hold
Event|Event|General Exam|5063,5068|false|false|false|||rails
Disorder|Disease or Syndrome|General Exam|5076,5079|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|5076,5079|false|false|false|||bed
Finding|Intellectual Product|General Exam|5076,5079|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|General Exam|5099,5104|false|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|General Exam|5109,5113|true|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|General Exam|5109,5113|true|false|false|C5781420||legs
Event|Event|General Exam|5114,5125|true|false|false|||antigravity
Event|Event|General Exam|5176,5187|false|false|false|||withdrawals
Anatomy|Body Part, Organ, or Organ Component|General Exam|5191,5208|false|false|false|C1140618|Upper Extremity|upper extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|5197,5208|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|5234,5245|false|false|false|||withdrawals
Anatomy|Body Location or Region|General Exam|5249,5254|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5249,5254|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5249,5266|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|5255,5266|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|5278,5285|false|false|false|||stimuli
Phenomenon|Phenomenon or Process|General Exam|5278,5285|false|false|false|C0234402|Stimulus|stimuli
Event|Event|General Exam|5290,5294|false|false|false|||says
Event|Event|General Exam|5304,5308|false|false|false|||DTRs
Finding|Gene or Genome|General Exam|5317,5320|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|5317,5320|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Disorder|Disease or Syndrome|General Exam|5325,5328|false|false|false|C0030587|Paroxysmal atrial tachycardia|Pat
Drug|Organic Chemical|General Exam|5325,5328|false|false|false|C2825250|Fenamole|Pat
Drug|Pharmacologic Substance|General Exam|5325,5328|false|false|false|C2825250|Fenamole|Pat
Event|Event|General Exam|5325,5328|false|false|false|||Pat
Finding|Molecular Function|General Exam|5325,5328|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|Pat
Procedure|Diagnostic Procedure|General Exam|5325,5328|false|false|false|C3897364|Thermoacoustic Computed Tomography|Pat
Disorder|Congenital Abnormality|General Exam|5329,5332|false|false|false|C0001080|Achondroplasia|Ach
Drug|Biologically Active Substance|General Exam|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Drug|Organic Chemical|General Exam|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Drug|Pharmacologic Substance|General Exam|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Event|Event|General Exam|5329,5332|false|false|false|||Ach
Finding|Gene or Genome|General Exam|5329,5332|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Finding|Sign or Symptom|General Exam|5329,5332|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Anatomy|Body Location or Region|General Exam|5380,5387|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|Plantar
Event|Event|General Exam|5388,5396|false|false|false|||response
Finding|Finding|General Exam|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|General Exam|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|General Exam|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Anatomy|Body Location or Region|General Exam|5401,5407|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Event|Event|General Exam|5423,5435|false|false|false|||Coordination
Finding|Functional Concept|General Exam|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Body Substance|General Exam|5437,5444|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5437,5444|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5437,5444|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5455,5466|true|false|false|||participate
Finding|Finding|General Exam|5469,5473|true|false|false|C0016928|Gait|Gait
Event|Event|General Exam|5485,5491|true|false|false|||assess
Finding|Body Substance|General Exam|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5513,5516|true|false|false|||get
Disorder|Disease or Syndrome|General Exam|5524,5527|true|true|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|5524,5527|true|false|false|||bed
Finding|Intellectual Product|General Exam|5524,5527|true|true|false|C2346952|Bachelor of Education|bed
Event|Event|General Exam|5529,5538|true|false|false|||Discharge
Finding|Body Substance|General Exam|5529,5538|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|5529,5538|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|5529,5538|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|5529,5538|true|false|false|C0030685|Patient Discharge|Discharge
Event|Event|General Exam|5539,5543|false|false|false|||Exam
Finding|Functional Concept|General Exam|5539,5543|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|5539,5543|false|false|false|C0582103|Medical Examination|Exam
Event|Event|General Exam|5545,5552|false|false|false|||General
Finding|Classification|General Exam|5545,5552|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|5545,5552|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|5554,5561|false|false|false|||sitting
Anatomy|Body Part, Organ, or Organ Component|General Exam|5583,5587|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|5583,5587|false|false|false|C5848506||eyes
Event|Event|General Exam|5588,5594|false|false|false|||closed
Anatomy|Body Location or Region|General Exam|5595,5600|false|false|false|C1512338|HEENT|HEENT
Disorder|Injury or Poisoning|General Exam|5605,5611|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|General Exam|5605,5611|true|false|false|||trauma
Procedure|Health Care Activity|General Exam|5605,5611|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|General Exam|5616,5624|true|false|false|||jaundice
Finding|Finding|General Exam|5616,5624|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|General Exam|5616,5624|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|General Exam|5629,5636|true|false|false|||lesions
Finding|Finding|General Exam|5629,5636|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|General Exam|5640,5650|true|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Space or Junction|General Exam|5656,5661|true|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|5656,5661|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|5656,5661|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|5656,5661|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|General Exam|5656,5673|true|false|false|C0085610;C2108107;C5235162|Sinus Bradycardia by ECG Finding;Sinus bradycardia;continuous electrocardiogram sinus bradycardia|sinus bradycardia
Finding|Pathologic Function|General Exam|5656,5673|true|false|false|C0085610;C2108107;C5235162|Sinus Bradycardia by ECG Finding;Sinus bradycardia;continuous electrocardiogram sinus bradycardia|sinus bradycardia
Event|Event|General Exam|5662,5673|true|false|false|||bradycardia
Finding|Finding|General Exam|5662,5673|true|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|General Exam|5684,5688|true|false|false|||Pulm
Procedure|Health Care Activity|General Exam|5684,5688|true|false|false|C1315068|Pulmonary ventilator management|Pulm
Disorder|Congenital Abnormality|General Exam|5719,5722|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|5719,5722|false|false|false|||Ext
Finding|Gene or Genome|General Exam|5719,5722|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|5724,5728|true|false|false|||Warm
Finding|Finding|General Exam|5724,5728|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|5724,5728|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|5733,5737|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|5738,5746|true|false|false|||perfused
Disorder|Disease or Syndrome|General Exam|5751,5755|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|5751,5755|true|false|false|||rash
Finding|Pathologic Function|General Exam|5751,5755|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|5751,5755|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|General Exam|5759,5767|true|false|false|||mottling
Finding|Finding|General Exam|5759,5767|true|false|false|C0302133|Mottling|mottling
Finding|Mental Process|General Exam|5783,5789|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|5783,5796|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|General Exam|5783,5796|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|General Exam|5790,5796|false|false|false|C5889824||Status
Event|Event|General Exam|5790,5796|false|false|false|||Status
Finding|Idea or Concept|General Exam|5790,5796|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|General Exam|5808,5817|false|false|false|||questions
Event|Event|General Exam|5834,5842|false|false|false|||sentence
Finding|Intellectual Product|General Exam|5834,5842|false|false|false|C0876929|Sentence|sentence
Event|Event|General Exam|5849,5854|false|false|false|||humor
Finding|Intellectual Product|General Exam|5849,5854|false|false|false|C0020168|Humor|humor
Procedure|Therapeutic or Preventive Procedure|General Exam|5849,5854|false|false|false|C0597811|Humor therapy|humor
Drug|Chemical Viewed Structurally|General Exam|5859,5866|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|General Exam|5867,5876|false|false|false|||sentences
Finding|Intellectual Product|General Exam|5867,5876|false|false|false|C0876929|Sentence|sentences
Event|Event|General Exam|5877,5885|false|false|false|||observed
Anatomy|Body Part, Organ, or Organ Component|General Exam|5893,5897|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|General Exam|5893,5897|false|false|false|C5848506||Eyes
Event|Event|General Exam|5913,5918|false|false|false|||close
Finding|Finding|General Exam|5913,5918|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|General Exam|5913,5918|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|General Exam|5932,5939|false|false|false|||talking
Event|Event|General Exam|5941,5947|true|false|false|||Speech
Finding|Organism Function|General Exam|5941,5947|true|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|5941,5947|true|false|false|C0846595|Speech assessment|Speech
Event|Event|General Exam|5955,5965|true|false|false|||dysarthric
Finding|Functional Concept|General Exam|5970,5981|true|false|false|C0205359|Spontaneous|spontaneous
Event|Event|General Exam|5982,5988|true|false|false|||speech
Finding|Organism Function|General Exam|5982,5988|true|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|General Exam|5982,5988|true|false|false|C0846595|Speech assessment|speech
Event|Event|General Exam|5989,5995|true|false|false|||output
Finding|Conceptual Entity|General Exam|5989,5995|true|false|false|C1709366|system output|output
Procedure|Health Care Activity|General Exam|5989,5995|true|false|false|C3251815|Measurement of fluid output|output
Finding|Gene or Genome|General Exam|6005,6011|false|false|false|C1424587|LITAF gene|simple
Event|Event|General Exam|6012,6020|false|false|false|||commands
Anatomy|Body Part, Organ, or Organ Component|General Exam|6024,6031|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|6024,6038|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|6024,6038|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|6032,6038|false|false|false|C0027740|Nerve|Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|6057,6063|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|6076,6080|true|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|6089,6098|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|6089,6098|true|false|false|||nystagmus
Anatomy|Body Location or Region|General Exam|6104,6110|false|false|false|C0015450|Face|facial
Finding|Finding|General Exam|6104,6120|false|false|false|C0517999|facial sensation|facial sensation
Event|Event|General Exam|6111,6120|false|false|false|||sensation
Finding|Finding|General Exam|6111,6120|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|6111,6120|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|6111,6120|false|false|false|C2229507|sensory exam|sensation
Finding|Finding|General Exam|6121,6127|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|6139,6142|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|6139,6142|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|6147,6153|true|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|General Exam|6147,6159|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|General Exam|6147,6159|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|General Exam|6154,6159|true|false|false|||droop
Anatomy|Body Location or Region|General Exam|6161,6167|true|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|General Exam|6168,6179|true|false|false|C1995013|Set of muscles|musculature
Event|Event|General Exam|6180,6189|true|false|false|||symmetric
Finding|Conceptual Entity|General Exam|6180,6189|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|6180,6189|true|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|General Exam|6195,6202|false|false|false|||grimace
Finding|Sign or Symptom|General Exam|6195,6202|false|false|false|C0239779|Grimaces|grimace
Finding|Functional Concept|General Exam|6207,6214|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|General Exam|6207,6214|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Anatomy|Body Location or Region|General Exam|6215,6221|false|false|false|C0015450|Face|facial
Event|Event|General Exam|6222,6231|false|false|false|||movements
Finding|Organism Function|General Exam|6222,6231|false|false|false|C0026649|Movement|movements
Anatomy|Body Part, Organ, or Organ Component|General Exam|6245,6251|false|false|false|C0700374|Palate|palate
Event|Event|General Exam|6252,6260|false|false|false|||elevates
Anatomy|Body Part, Organ, or Organ Component|General Exam|6276,6282|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|6276,6282|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|General Exam|6276,6282|false|false|false|C0872394|Procedure on tongue|tongue
Finding|Finding|General Exam|6276,6290|false|false|false|C3693372|tongue midline|tongue midline
Anatomy|Cell Component|General Exam|6283,6290|false|false|false|C1660780|midline cell component|midline
Finding|Functional Concept|General Exam|6293,6298|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|6307,6311|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|6307,6311|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|6307,6311|false|false|false|||bulk
Event|Event|General Exam|6313,6317|false|false|false|||tone
Event|Activity|General Exam|6330,6337|false|false|false|C0206244|Lifting|Lifting
Anatomy|Body Part, Organ, or Organ Component|General Exam|6338,6342|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|6338,6342|false|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|6338,6342|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|General Exam|6338,6342|false|false|false|||arms
Finding|Gene or Genome|General Exam|6338,6342|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|6338,6342|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|General Exam|6338,6351|false|false|false|C0015385|Limb structure|arms and legs
Anatomy|Body Part, Organ, or Organ Component|General Exam|6347,6351|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|General Exam|6347,6351|false|false|false|C5781420||legs
Phenomenon|Natural Phenomenon or Process|General Exam|6360,6367|true|false|false|C0282189|Gravity (physical force)|gravity
Attribute|Clinical Attribute|General Exam|6384,6394|true|false|false|C1442099|Resistance|resistance
Event|Event|General Exam|6384,6394|true|false|false|||resistance
Finding|Mental Process|General Exam|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Physiologic Function|General Exam|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Social Behavior|General Exam|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Event|Event|General Exam|6412,6421|false|false|false|||Sensation
Finding|Finding|General Exam|6412,6421|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|6412,6421|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|6412,6421|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|6422,6428|false|false|false|||intact
Finding|Finding|General Exam|6422,6428|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|6432,6437|false|false|false|||touch
Finding|Mental Process|General Exam|6432,6437|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|6432,6437|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|6432,6437|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|6442,6453|false|false|false|||temperature
Procedure|Health Care Activity|General Exam|6442,6453|false|false|false|C0886414|Body temperature measurement|temperature
Event|Event|General Exam|6467,6471|false|false|false|||DTRs
Anatomy|Body Part, Organ, or Organ Component|General Exam|6476,6484|false|false|false|C0030647|Patella|patellar
Anatomy|Body Part, Organ, or Organ Component|General Exam|6486,6492|false|false|false|C0559499|Biceps brachii muscle structure|biceps
Anatomy|Body Part, Organ, or Organ Component|General Exam|6494,6509|false|false|false|C0224264|Structure of brachioradialis muscle|brachioradialis
Event|Event|General Exam|6523,6535|false|false|false|||Coordination
Finding|Functional Concept|General Exam|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|General Exam|6540,6549|true|false|false|||dysmetria
Finding|Finding|General Exam|6540,6549|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Event|Event|General Exam|6553,6559|true|false|false|||tremor
Finding|Sign or Symptom|General Exam|6553,6559|true|false|false|C0040822|Tremor|tremor
Finding|Finding|General Exam|6564,6568|false|false|false|C0016928|Gait|Gait
Finding|Finding|General Exam|6580,6584|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|General Exam|6618,6627|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|General Exam|6628,6632|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|General Exam|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|6664,6671|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|6664,6671|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|6664,6671|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|6675,6679|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|6675,6679|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|6675,6679|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|6675,6679|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|6675,6679|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|6694,6700|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|6694,6700|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|6694,6700|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|6706,6715|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|6706,6715|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|6706,6715|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|6720,6728|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|6720,6728|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|6720,6728|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|6720,6728|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|6739,6742|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|6739,6742|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|6739,6742|false|false|false|||CO2
Finding|Finding|General Exam|6739,6742|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|6739,6742|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|6746,6751|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|6746,6755|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|6746,6755|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|6746,6755|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|6752,6755|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|6752,6755|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|6752,6755|false|false|false|||GAP
Finding|Gene or Genome|General Exam|6752,6755|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|General Exam|6773,6776|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|6773,6776|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|6773,6776|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|6773,6776|false|false|false|||ALT
Finding|Gene or Genome|General Exam|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|6773,6776|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|6777,6781|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|6777,6781|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|General Exam|6777,6781|false|false|false|||SGPT
Finding|Gene or Genome|General Exam|6777,6781|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|6777,6781|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|6785,6788|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|6785,6788|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|6785,6788|false|false|false|||AST
Finding|Gene or Genome|General Exam|6785,6788|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|6789,6793|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|6789,6793|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|General Exam|6789,6793|false|false|false|||SGOT
Finding|Gene or Genome|General Exam|6789,6793|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|6789,6793|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|6798,6801|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|6798,6801|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|General Exam|6798,6801|false|false|false|||ALK
Finding|Gene or Genome|General Exam|6798,6801|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|6798,6801|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|General Exam|6798,6806|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|General Exam|6798,6806|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|General Exam|6798,6806|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|General Exam|6802,6806|false|false|false|||PHOS
Drug|Biologically Active Substance|General Exam|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|General Exam|6838,6845|false|false|false|||CALCIUM
Finding|Physiologic Function|General Exam|6838,6845|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|6838,6845|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Event|Event|General Exam|6850,6859|false|false|false|||PHOSPHATE
Procedure|Laboratory Procedure|General Exam|6850,6859|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|6864,6873|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|General Exam|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Drug|Enzyme|General Exam|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Drug|Pharmacologic Substance|General Exam|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Event|Event|General Exam|6892,6895|false|false|false|||tTG
Finding|Gene or Genome|General Exam|6892,6895|false|false|false|C5575307|TGM2 wt Allele|tTG
Drug|Amino Acid, Peptide, or Protein|General Exam|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Immunologic Factor|General Exam|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Pharmacologic Substance|General Exam|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Event|Event|General Exam|6896,6899|false|false|false|||IgA
Finding|Gene or Genome|General Exam|6896,6899|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|IgA
Procedure|Laboratory Procedure|General Exam|6896,6899|false|false|false|C0202083|Immunoglobulin A measurement|IgA
Anatomy|Cell|General Exam|6916,6919|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6924,6927|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6924,6927|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6924,6927|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6934,6937|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|6934,6937|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|6934,6937|false|false|false|||HGB
Finding|Gene or Genome|General Exam|6934,6937|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|6934,6937|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|General Exam|6943,6946|false|false|false|||HCT
Procedure|Laboratory Procedure|General Exam|6943,6946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|6943,6946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|6952,6955|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|6952,6955|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|6952,6955|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6952,6955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6952,6955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6960,6963|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6960,6963|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6960,6963|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6960,6963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6960,6963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6960,6963|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6969,6973|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6969,6973|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|7013,7016|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|7013,7016|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Body Substance|General Exam|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|7052,7058|false|false|false|||RANDOM
Finding|Body Substance|General Exam|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Classification|General Exam|7082,7090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|7082,7090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|7082,7090|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Body Substance|General Exam|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|7119,7122|false|false|false|||NEG
Finding|Finding|General Exam|7119,7122|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|7132,7135|false|false|false|C5848551|Neg - answer|NEG
Drug|Hazardous or Poisonous Substance|General Exam|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Organic Chemical|General Exam|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Pharmacologic Substance|General Exam|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Event|Event|General Exam|7136,7143|false|false|false|||opiates
Procedure|Laboratory Procedure|General Exam|7136,7143|false|false|false|C0242401|Opiate Measurement|opiates
Event|Event|General Exam|7144,7147|false|false|false|||NEG
Finding|Finding|General Exam|7144,7147|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|General Exam|7149,7156|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|General Exam|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|General Exam|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|General Exam|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|General Exam|7149,7156|false|false|false|C0009170|cocaine|cocaine
Event|Event|General Exam|7149,7156|false|false|false|||cocaine
Procedure|Laboratory Procedure|General Exam|7149,7156|false|false|false|C0202362|Cocaine measurement|cocaine
Event|Event|General Exam|7157,7160|false|false|false|||NEG
Finding|Finding|General Exam|7157,7160|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|7170,7173|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|7182,7185|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|7194,7197|false|false|false|||NEG
Finding|Finding|General Exam|7194,7197|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|7210,7222|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|7217,7222|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|7217,7222|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|General Exam|7217,7222|false|false|false|||COLOR
Drug|Organic Chemical|General Exam|7223,7228|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|General Exam|7236,7241|false|false|false|||Clear
Finding|Idea or Concept|General Exam|7236,7241|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|7261,7273|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|7268,7273|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7268,7273|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7268,7273|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|7274,7276|false|false|false|||LG
Drug|Biologically Active Substance|General Exam|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Event|Event|General Exam|7286,7289|false|false|false|||NEG
Finding|Finding|General Exam|7286,7289|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|7290,7297|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|7290,7297|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|General Exam|7290,7297|false|false|false|||PROTEIN
Finding|Conceptual Entity|General Exam|7290,7297|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|7290,7297|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|General Exam|7298,7301|false|false|false|||NEG
Finding|Finding|General Exam|7298,7301|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|7303,7310|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|7303,7310|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|7303,7310|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|General Exam|7311,7314|false|false|false|||NEG
Finding|Finding|General Exam|7311,7314|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|7315,7321|false|false|false|C0022634|Ketones|KETONE
Drug|Biologically Active Substance|General Exam|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|7326,7335|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|General Exam|7336,7339|false|false|false|||NEG
Finding|Finding|General Exam|7336,7339|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|7350,7353|false|false|false|||NEG
Finding|Finding|General Exam|7350,7353|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|7367,7370|false|false|false|||NEG
Finding|Finding|General Exam|7367,7370|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|7383,7393|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|General Exam|7390,7393|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7390,7393|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7390,7393|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|7397,7400|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|General Exam|7403,7411|true|false|false|C1510439|bacteria aspects|BACTERIA
Event|Event|General Exam|7412,7415|true|false|false|||FEW
Drug|Food|General Exam|7417,7422|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|7417,7422|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|7417,7422|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|7417,7422|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|General Exam|7423,7427|false|false|false|||NONE
Disorder|Disease or Syndrome|General Exam|7429,7432|true|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|7429,7432|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|7429,7432|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|7429,7432|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|7429,7432|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|7429,7432|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|General Exam|7429,7432|true|false|false|||EPI
Finding|Gene or Genome|General Exam|7429,7432|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|7429,7432|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|7429,7432|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|General Exam|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|7447,7460|false|false|false|C0455910|Mucus in urine (finding)|URINE  MUCOUS
Finding|Body Substance|General Exam|7454,7460|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|MUCOUS
Event|Event|General Exam|7461,7465|false|false|false|||RARE
Finding|Gene or Genome|General Exam|7461,7465|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Disorder|Neoplastic Process|General Exam|7485,7488|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|7485,7488|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|7485,7488|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Anatomy|Cell|General Exam|7512,7515|false|false|false|C0023516|Leukocytes|WBC
Event|Event|General Exam|7512,7515|false|false|false|||WBC
Anatomy|Cell|General Exam|7520,7523|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7520,7523|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7520,7523|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|7529,7532|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|7529,7532|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|7529,7532|false|false|false|||HGB
Finding|Gene or Genome|General Exam|7529,7532|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|7529,7532|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|General Exam|7538,7541|false|false|false|||HCT
Procedure|Laboratory Procedure|General Exam|7538,7541|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|7538,7541|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|7547,7550|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|7547,7550|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|7547,7550|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|7547,7550|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|7547,7550|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|7555,7558|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|7555,7558|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|7555,7558|false|false|false|||MCH
Finding|Gene or Genome|General Exam|7555,7558|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|7555,7558|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|7555,7558|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|7564,7568|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|7564,7568|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|7608,7613|false|false|false|||NEUTS
Drug|Antibiotic|General Exam|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|7633,7636|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|General Exam|7633,7636|false|false|false|||EOS
Finding|Gene or Genome|General Exam|7633,7636|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|General Exam|7740,7743|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|7740,7743|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Classification|General Exam|7772,7775|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|PO2
Finding|Molecular Function|General Exam|7772,7775|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|PO2
Procedure|Laboratory Procedure|General Exam|7772,7775|false|false|false|C1283004|PO2 measurement|PO2
Lab|Laboratory or Test Result|General Exam|7780,7784|false|false|false|C0391839|Carbon dioxide, partial pressure|PCO2
Procedure|Laboratory Procedure|General Exam|7780,7784|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|PCO2
Drug|Biologically Active Substance|General Exam|7804,7807|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|7804,7807|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|7804,7807|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|7804,7807|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Anatomy|Body Location or Region|General Exam|7811,7815|false|false|false|C2987514|Anatomical base|BASE
Drug|Biomedical or Dental Material|General Exam|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Chemical Viewed Functionally|General Exam|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Finding|Gene or Genome|General Exam|7811,7815|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Finding|Idea or Concept|General Exam|7811,7815|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Event|Event|General Exam|7821,7829|false|false|false|||COMMENTS
Finding|Intellectual Product|General Exam|7821,7829|false|false|false|C0282411;C0947611|Comment;Published Comment|COMMENTS
Event|Event|General Exam|7836,7839|false|false|false|||TOP
Drug|Biologically Active Substance|General Exam|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|7854,7861|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|7854,7861|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|7854,7861|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|7865,7869|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|7865,7869|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|7865,7869|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|7865,7869|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|7865,7869|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|7884,7890|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|7884,7890|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|7884,7890|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|7896,7905|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|7896,7905|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|7896,7905|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|7910,7918|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|7910,7918|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|7910,7918|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|7910,7918|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|7929,7932|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|7929,7932|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|7929,7932|false|false|false|||CO2
Finding|Finding|General Exam|7929,7932|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|7929,7932|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|7936,7941|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|7936,7945|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|7936,7945|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|7936,7945|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|7942,7945|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|7942,7945|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|7942,7945|false|false|false|||GAP
Finding|Gene or Genome|General Exam|7942,7945|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|General Exam|7995,7998|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|7995,7998|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|7995,7998|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|7995,7998|false|false|false|||ALT
Finding|Gene or Genome|General Exam|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|7995,7998|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|7999,8003|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|7999,8003|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|General Exam|7999,8003|false|false|false|||SGPT
Finding|Gene or Genome|General Exam|7999,8003|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|7999,8003|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|8007,8010|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|8007,8010|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|8007,8010|false|false|false|||AST
Finding|Gene or Genome|General Exam|8007,8010|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|8011,8015|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|8011,8015|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|General Exam|8011,8015|false|false|false|||SGOT
Finding|Gene or Genome|General Exam|8011,8015|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|8011,8015|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|8023,8026|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|8023,8026|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|8023,8026|false|false|false|||CPK
Finding|Gene or Genome|General Exam|8023,8026|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|8023,8026|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|8031,8034|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|8031,8034|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|General Exam|8031,8034|false|false|false|||ALK
Finding|Gene or Genome|General Exam|8031,8034|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|8031,8034|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|General Exam|8071,8076|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|8071,8076|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|8071,8076|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|8071,8076|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|General Exam|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|General Exam|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|General Exam|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|General Exam|8094,8101|false|false|false|||ALBUMIN
Finding|Gene or Genome|General Exam|8094,8101|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|General Exam|8094,8101|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|General Exam|8094,8101|false|false|false|C0201838|Albumin measurement|ALBUMIN
Drug|Biologically Active Substance|General Exam|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|General Exam|8106,8113|false|false|false|||CALCIUM
Finding|Physiologic Function|General Exam|8106,8113|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|8106,8113|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|8118,8127|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|8133,8142|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Event|Event|General Exam|8161,8164|false|false|false|||VIT
Finding|Gene or Genome|General Exam|8161,8164|false|false|false|C1421454;C5401427;C5401428|AML Vitals Table;EWS Vitals Table;VIT gene|VIT
Finding|Intellectual Product|General Exam|8161,8164|false|false|false|C1421454;C5401427;C5401428|AML Vitals Table;EWS Vitals Table;VIT gene|VIT
Procedure|Therapeutic or Preventive Procedure|General Exam|8161,8164|false|false|false|C1831721|VIT Regimen|VIT
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Organic Chemical|General Exam|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Pharmacologic Substance|General Exam|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Vitamin|General Exam|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Event|Event|General Exam|8165,8168|false|false|false|||B12
Finding|Gene or Genome|General Exam|8165,8168|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Attribute|Clinical Attribute|General Exam|8188,8191|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Event|Event|General Exam|8188,8191|false|false|false|||TSH
Procedure|Laboratory Procedure|General Exam|8188,8191|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Attribute|Clinical Attribute|General Exam|8210,8213|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Event|Event|General Exam|8210,8213|false|false|false|||TSH
Procedure|Laboratory Procedure|General Exam|8210,8213|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|8250,8253|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|General Exam|8250,8253|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Event|Event|General Exam|8250,8253|false|false|false|||CRP
Finding|Gene or Genome|General Exam|8250,8253|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Event|Event|General Exam|8259,8264|false|false|false|||dsDNA
Event|Event|General Exam|8265,8273|false|false|false|||NEGATIVE
Finding|Classification|General Exam|8265,8273|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|8265,8273|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|8265,8273|false|false|false|C5237010|Expression Negative|NEGATIVE
Drug|Amino Acid, Peptide, or Protein|General Exam|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|General Exam|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|General Exam|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|General Exam|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|General Exam|8315,8318|false|false|false|||ASA
Finding|Gene or Genome|General Exam|8315,8318|false|false|false|C1412553|ARSA gene|ASA
Event|Event|General Exam|8319,8322|false|false|false|||NEG
Finding|Finding|General Exam|8319,8322|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|General Exam|8323,8330|false|false|false|C0161679|Toxic effect of ethyl alcohol|ETHANOL
Drug|Organic Chemical|General Exam|8323,8330|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Drug|Pharmacologic Substance|General Exam|8323,8330|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Event|Event|General Exam|8323,8330|false|false|false|||ETHANOL
Procedure|Laboratory Procedure|General Exam|8323,8330|false|false|false|C0202304|Ethanol measurement|ETHANOL
Event|Event|General Exam|8331,8334|false|false|false|||NEG
Finding|Finding|General Exam|8331,8334|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|8345,8348|false|false|false|||NEG
Finding|Finding|General Exam|8345,8348|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|8360,8363|false|false|false|||NEG
Finding|Finding|General Exam|8360,8363|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|8365,8368|false|false|false|||EEG
Procedure|Diagnostic Procedure|General Exam|8365,8368|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|General Exam|8389,8399|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|8389,8399|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|8389,8399|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|General Exam|8406,8415|true|false|false|||telemetry
Procedure|Diagnostic Procedure|General Exam|8406,8415|true|false|false|C0039451|Telemetry|telemetry
Event|Event|General Exam|8416,8424|true|false|false|||captured
Event|Event|General Exam|8439,8450|true|false|false|||activations
Event|Event|General Exam|8457,8467|false|false|false|||background
Finding|Conceptual Entity|General Exam|8457,8467|false|false|false|C1706907|Background|background
Event|Event|General Exam|8468,8474|false|false|false|||showed
Event|Event|General Exam|8482,8488|false|false|false|||waking
Finding|Physiologic Function|General Exam|8482,8488|false|false|false|C0442696|Waking|waking
Drug|Organic Chemical|General Exam|8493,8498|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|General Exam|8493,8498|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|General Exam|8493,8498|false|false|false|C0037313|Sleep|sleep
Event|Event|General Exam|8499,8507|false|false|false|||patterns
Disorder|Congenital Abnormality|General Exam|8530,8543|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|8530,8543|true|false|false|||abnormalities
Finding|Functional Concept|General Exam|8530,8543|true|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|8558,8566|true|false|false|||features
Event|Event|General Exam|8587,8595|false|false|false|||seizures
Finding|Sign or Symptom|General Exam|8587,8595|false|false|false|C0036572|Seizures|seizures
Event|Event|General Exam|8599,8610|false|false|false|||bradycardia
Finding|Finding|General Exam|8599,8610|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|General Exam|8615,8620|false|false|false|||noted
Event|Event|General Exam|8624,8631|false|false|false|||IMAGING
Finding|Finding|General Exam|8624,8631|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|8624,8631|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|8642,8645|true|false|false|||MRI
Finding|Gene or Genome|General Exam|8642,8645|true|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|General Exam|8642,8645|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|General Exam|8642,8645|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|General Exam|8642,8651|true|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI BRAIN
Anatomy|Body Part, Organ, or Organ Component|General Exam|8646,8651|true|false|false|C0006104;C4266577|Brain;Head>Brain|BRAIN
Disorder|Disease or Syndrome|General Exam|8646,8651|true|false|false|C0006111|Brain Diseases|BRAIN
Event|Event|General Exam|8646,8651|true|false|false|||BRAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|8665,8673|true|false|false|C0009924|Contrast Media|CONTRAST
Drug|Organic Chemical|Findings|8701,8706|false|false|false|C0309093|FLAIR (product)|FLAIR
Drug|Pharmacologic Substance|Findings|8701,8706|false|false|false|C0309093|FLAIR (product)|FLAIR
Procedure|Diagnostic Procedure|Findings|8701,8706|false|false|false|C2826145|Fluid Attenuated Inversion Recovery|FLAIR
Event|Event|Findings|8707,8718|false|false|false|||hypointense
Finding|Idea or Concept|Findings|8726,8736|false|false|false|C1517605|Isointense|isointense
Event|Event|Findings|8737,8743|false|false|false|||lesion
Finding|Finding|Findings|8737,8743|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Findings|8737,8743|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Cell Component|Findings|8747,8754|false|false|false|C1660780|midline cell component|midline
Disorder|Disease or Syndrome|Findings|8769,8777|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Findings|8769,8777|false|false|false|||anterior
Disorder|Disease or Syndrome|Findings|8782,8791|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|Findings|8782,8801|false|false|false|C0032009;C0447640|Pituitary Gland, Posterior;pars nervosa of hypophysis|posterior pituitary
Drug|Amino Acid, Peptide, or Protein|Findings|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Hormone|Findings|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Pharmacologic Substance|Findings|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Anatomy|Body Part, Organ, or Organ Component|Findings|8792,8801|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|Findings|8792,8801|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|Findings|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|Findings|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|Findings|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Event|Event|Findings|8792,8801|false|false|false|||pituitary
Event|Event|Findings|8805,8810|false|false|false|||noted
Event|Event|Findings|8824,8832|true|false|false|||evidence
Finding|Idea or Concept|Findings|8824,8832|true|false|false|C3887511|Evidence|evidence
Event|Event|Findings|8838,8848|true|false|false|||hemorrhage
Finding|Pathologic Function|Findings|8838,8848|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|Findings|8850,8855|true|false|false|C1717255||edema
Event|Event|Findings|8850,8855|true|false|false|||edema
Finding|Pathologic Function|Findings|8850,8855|true|false|false|C0013604|Edema|edema
Finding|Finding|Findings|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Findings|8857,8868|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|Findings|8862,8868|false|false|false|||effect
Anatomy|Cell Component|Findings|8870,8877|false|false|false|C1660780|midline cell component|midline
Finding|Finding|Findings|8870,8883|false|false|false|C4086580|Midline Shift|midline shift
Event|Event|Findings|8878,8883|false|false|false|||shift
Finding|Functional Concept|Findings|8878,8883|false|false|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|Findings|8878,8883|false|false|false|C2347509|Physical Shift|shift
Event|Event|Findings|8887,8897|false|false|false|||infarction
Finding|Pathologic Function|Findings|8887,8897|false|false|false|C0021308|Infarction|infarction
Anatomy|Body Part, Organ, or Organ Component|Findings|8904,8914|false|false|false|C0018827|Heart Ventricle|ventricles
Event|Event|Findings|8919,8924|false|false|false|||sulci
Event|Event|Findings|8929,8935|false|false|false|||normal
Event|Event|Findings|8939,8946|false|false|false|||caliber
Event|Event|Findings|8951,8964|false|false|false|||configuration
Finding|Conceptual Entity|Findings|8951,8964|false|false|false|C2827597|Computer Configuration|configuration
Finding|Finding|Findings|8979,8987|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Findings|8979,8987|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Activity|Findings|8988,8999|true|false|false|C2349975|Enhance (action)|enhancement
Event|Event|Findings|8988,8999|true|false|false|||enhancement
Procedure|Therapeutic or Preventive Procedure|Findings|8988,8999|true|false|false|C1627358|Refractive surgery enhancement|enhancement
Drug|Indicator, Reagent, or Diagnostic Aid|Findings|9006,9014|true|false|false|C0009924|Contrast Media|contrast
Event|Event|Findings|9015,9029|true|false|false|||administration
Event|Occupational Activity|Findings|9015,9029|true|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Findings|9015,9029|true|false|false|C1533734|Administration (procedure)|administration
Drug|Organic Chemical|Impression|9059,9064|false|false|false|C0309093|FLAIR (product)|FLAIR
Drug|Pharmacologic Substance|Impression|9059,9064|false|false|false|C0309093|FLAIR (product)|FLAIR
Procedure|Diagnostic Procedure|Impression|9059,9064|false|false|false|C2826145|Fluid Attenuated Inversion Recovery|FLAIR
Event|Event|Impression|9065,9076|false|false|false|||hypointense
Finding|Idea or Concept|Impression|9084,9094|false|false|false|C1517605|Isointense|isointense
Event|Event|Impression|9095,9101|false|false|false|||lesion
Finding|Finding|Impression|9095,9101|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|9095,9101|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Cell Component|Impression|9105,9112|false|false|false|C1660780|midline cell component|midline
Disorder|Disease or Syndrome|Impression|9127,9135|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Impression|9127,9135|false|false|false|||anterior
Disorder|Disease or Syndrome|Impression|9140,9149|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|Impression|9140,9159|false|false|false|C0032009;C0447640|Pituitary Gland, Posterior;pars nervosa of hypophysis|posterior pituitary
Drug|Amino Acid, Peptide, or Protein|Impression|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Hormone|Impression|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Pharmacologic Substance|Impression|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Anatomy|Body Part, Organ, or Organ Component|Impression|9150,9159|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|Impression|9150,9159|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|Impression|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|Impression|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|Impression|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Finding|Finding|Impression|9160,9166|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Impression|9160,9166|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Impression|9167,9177|false|false|false|||represents
Disorder|Anatomical Abnormality|Impression|9196,9200|false|false|false|C0010709|Cyst|cyst
Event|Event|Impression|9196,9200|false|false|false|||cyst
Finding|Body Substance|Impression|9196,9200|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Impression|9196,9200|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|Impression|9212,9222|false|false|false|||evaluation
Finding|Idea or Concept|Impression|9212,9222|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Impression|9212,9222|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|Impression|9226,9232|false|false|false|||needed
Event|Event|Impression|9234,9243|false|false|false|||dedicated
Anatomy|Body Part, Organ, or Organ Component|Impression|9244,9253|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|Impression|9244,9253|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|Impression|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|Impression|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|Impression|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Event|Event|Impression|9254,9256|false|false|false|||MR
Event|Event|Impression|9265,9273|false|false|false|||obtained
Finding|Intellectual Product|Hospital Course|9309,9318|false|false|false|C2349155|Worksheet|worksheet
Attribute|Clinical Attribute|Hospital Course|9321,9332|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9321,9332|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9321,9332|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9321,9332|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|9321,9345|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|9336,9345|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|9336,9345|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|9347,9357|false|false|false|C0015620|famotidine|famotidine
Drug|Pharmacologic Substance|Hospital Course|9347,9357|false|false|false|C0015620|famotidine|famotidine
Event|Event|Hospital Course|9347,9357|false|false|false|||famotidine
Finding|Finding|Hospital Course|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Finding|Intellectual Product|Hospital Course|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Finding|Organism Function|Hospital Course|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9370,9383|false|false|false|C0700589|Contraceptive methods|birth control
Drug|Organic Chemical|Hospital Course|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|9376,9383|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|Hospital Course|9435,9445|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|9435,9445|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|Hospital Course|9467,9477|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|9467,9477|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|Hospital Course|9467,9477|false|false|false|||Metoprolol
Drug|Organic Chemical|Hospital Course|9467,9486|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|9467,9486|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|9478,9486|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|9478,9486|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Organic Chemical|Hospital Course|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|9510,9523|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|9526,9534|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|9526,9534|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|9537,9540|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9537,9540|false|false|false|||TAB
Finding|Intellectual Product|Hospital Course|9614,9618|false|false|false|C1720092|Once - dosing instruction fragment|ONCE
Attribute|Clinical Attribute|Hospital Course|9620,9629|false|false|false|C3854082||Prognosis
Event|Event|Hospital Course|9620,9629|false|false|false|||Prognosis
Procedure|Health Care Activity|Hospital Course|9620,9629|false|false|false|C0033325|Forecast of outcome|Prognosis
Finding|Idea or Concept|Hospital Course|9631,9635|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Event|Activity|Hospital Course|9666,9670|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|9666,9670|false|false|false|C2828567|PRSS30P gene|Disp
Event|Event|Hospital Course|9680,9687|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9680,9687|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|9695,9704|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9695,9704|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9695,9716|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9695,9716|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9705,9716|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|9705,9716|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|9705,9716|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|9718,9726|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9718,9726|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|9718,9731|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|9727,9731|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|9727,9731|false|false|false|||Care
Finding|Finding|Hospital Course|9727,9731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|9727,9731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|9734,9742|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|9734,9742|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|9750,9759|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9750,9759|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9750,9769|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9760,9769|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9760,9769|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9760,9769|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9760,9769|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9760,9769|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Conceptual Entity|Hospital Course|9771,9781|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Finding|Functional Concept|Hospital Course|9771,9781|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Disorder|Disease or Syndrome|Hospital Course|9795,9803|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|9795,9803|false|false|false|||syndrome
Finding|Mental Process|Discharge Condition|9829,9835|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9829,9842|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9829,9842|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9836,9842|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9836,9842|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9844,9849|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|9844,9849|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|9854,9862|false|false|false|||coherent
Finding|Finding|Discharge Condition|9854,9862|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|9864,9869|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|9864,9886|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9864,9886|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|9873,9886|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|9873,9886|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9873,9886|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Event|Event|Discharge Condition|9888,9897|false|false|false|||Lethargic
Finding|Sign or Symptom|Discharge Condition|9888,9897|false|false|false|C0023380|Lethargy|Lethargic
Event|Event|Discharge Condition|9902,9911|false|false|false|||arousable
Event|Activity|Discharge Condition|9913,9921|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9913,9921|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9913,9921|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9922,9928|false|false|false|C5889824||Status
Event|Event|Discharge Condition|9922,9928|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|9922,9928|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9930,9940|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9930,9940|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|9943,9954|false|false|false|||Independent
Finding|Finding|Discharge Condition|9943,9954|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|9943,9954|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|9983,9987|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|10007,10015|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|10007,10015|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|10007,10015|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|10023,10027|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|10023,10027|false|false|false|||care
Finding|Finding|Discharge Instructions|10023,10027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10023,10027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10023,10030|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|Discharge Instructions|10065,10073|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10085,10093|false|false|false|||headache
Finding|Sign or Symptom|Discharge Instructions|10085,10093|false|false|false|C0018681|Headache|headache
Event|Event|Discharge Instructions|10095,10103|false|false|false|||lethargy
Finding|Sign or Symptom|Discharge Instructions|10095,10103|false|false|false|C0023380|Lethargy|lethargy
Event|Event|Discharge Instructions|10110,10118|false|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|10110,10118|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Drug|Biologically Active Substance|Discharge Instructions|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Discharge Instructions|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Discharge Instructions|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Discharge Instructions|10128,10132|false|false|false|C0337439|Iron measurement|iron
Event|Event|Discharge Instructions|10133,10141|false|false|false|||infusion
Finding|Functional Concept|Discharge Instructions|10133,10141|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10133,10141|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|Discharge Instructions|10154,10160|false|false|false|||number
Finding|Idea or Concept|Discharge Instructions|10154,10160|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Event|Discharge Instructions|10164,10169|false|false|false|||tests
Finding|Intellectual Product|Discharge Instructions|10164,10169|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|Discharge Instructions|10164,10169|false|false|false|C0022885|Laboratory Procedures|tests
Finding|Idea or Concept|Discharge Instructions|10187,10195|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10216,10226|false|false|false|||reassuring
Procedure|Health Care Activity|Discharge Instructions|10216,10226|false|false|false|C0557055|Reassuring (procedure)|reassuring
Event|Event|Discharge Instructions|10231,10234|true|false|false|||MRI
Finding|Gene or Genome|Discharge Instructions|10231,10234|true|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Discharge Instructions|10231,10234|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Discharge Instructions|10231,10234|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10243,10248|true|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|10243,10248|true|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|10249,10255|true|false|false|||showed
Event|Event|Discharge Instructions|10259,10267|true|false|false|||evidence
Finding|Idea or Concept|Discharge Instructions|10259,10267|true|false|false|C3887511|Evidence|evidence
Disorder|Disease or Syndrome|Discharge Instructions|10272,10278|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Discharge Instructions|10272,10278|true|false|false|||stroke
Finding|Finding|Discharge Instructions|10272,10278|true|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Discharge Instructions|10282,10294|true|false|false|||inflammation
Finding|Pathologic Function|Discharge Instructions|10282,10294|true|false|false|C0021368|Inflammation|inflammation
Event|Event|Discharge Instructions|10299,10302|false|false|false|||EEG
Procedure|Diagnostic Procedure|Discharge Instructions|10299,10302|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|Discharge Instructions|10306,10313|true|false|false|||monitor
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10319,10324|true|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|10319,10324|true|false|false|C0006111|Brain Diseases|brain
Finding|Organ or Tissue Function|Discharge Instructions|10319,10330|true|false|false|C0678909|Brain Waves|brain waves
Event|Event|Discharge Instructions|10325,10330|true|false|false|||waves
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|10325,10330|true|false|false|C0678544||waves
Event|Event|Discharge Instructions|10332,10338|true|false|false|||showed
Event|Event|Discharge Instructions|10342,10350|true|false|false|||evidence
Finding|Idea or Concept|Discharge Instructions|10342,10350|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|10342,10353|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Discharge Instructions|10354,10361|true|false|false|||seizure
Finding|Sign or Symptom|Discharge Instructions|10354,10361|true|false|false|C0036572|Seizures|seizure
Event|Event|Discharge Instructions|10368,10376|false|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|10368,10376|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Discharge Instructions|10387,10395|false|false|false|||improved
Event|Event|Discharge Instructions|10421,10436|false|false|false|||hospitalization
Procedure|Health Care Activity|Discharge Instructions|10421,10436|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Discharge Instructions|10446,10454|false|false|false|||continue
Event|Event|Discharge Instructions|10459,10466|false|false|false|||improve
Event|Event|Discharge Instructions|10477,10482|false|false|false|||leave
Event|Event|Discharge Instructions|10487,10495|false|false|false|||hospital
Finding|Idea or Concept|Discharge Instructions|10487,10495|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10505,10512|false|false|false|||leaving
Finding|Idea or Concept|Discharge Instructions|10517,10525|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10538,10546|false|false|false|||continue
Event|Event|Discharge Instructions|10550,10554|false|false|false|||work
Event|Event|Discharge Instructions|10559,10568|false|false|false|||improving
Event|Event|Discharge Instructions|10574,10582|false|false|false|||strength
Finding|Idea or Concept|Discharge Instructions|10574,10582|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|Discharge Instructions|10592,10599|false|false|false|||improve
Event|Event|Discharge Instructions|10615,10619|false|false|false|||work
Disorder|Disease or Syndrome|Discharge Instructions|10644,10648|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|10644,10648|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|10644,10648|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|10659,10663|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|10659,10663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|10659,10663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|10659,10668|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|10659,10668|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|10671,10679|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10680,10692|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10680,10692|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10680,10692|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

