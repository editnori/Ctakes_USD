 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|40,49|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|40,49|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|40,54|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|74,83|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|74,83|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|74,88|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|130,133|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|141,148|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|141,148|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|150,158|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|173,181|false|false|false|C0040610|tramadol|Tramadol
Drug|Pharmacologic Substance|Allergies|173,181|false|false|false|C0040610|tramadol|Tramadol
Event|Event|Allergies|173,181|false|false|false|||Tramadol
Procedure|Laboratory Procedure|Allergies|173,181|false|false|false|C1266765|Tramadol measurement (procedure)|Tramadol
Event|Event|Allergies|184,193|false|false|false|||Attending
Finding|Functional Concept|Allergies|184,193|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|219,228|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|Chief Complaint|219,239|false|false|false|C0000731|Abdomen distended|Abdominal distention
Event|Event|Chief Complaint|229,239|false|false|false|||distention
Finding|Finding|Chief Complaint|229,239|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Chief Complaint|229,239|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Sign or Symptom|Chief Complaint|241,250|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Chief Complaint|246,250|false|false|false|C2598155||pain
Event|Event|Chief Complaint|246,250|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|246,250|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|246,250|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Chief Complaint|252,257|false|false|false|||fever
Finding|Finding|Chief Complaint|252,257|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Chief Complaint|252,257|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|Chief Complaint|259,271|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Chief Complaint|259,271|false|false|false|||leukocytosis
Finding|Finding|Chief Complaint|259,271|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Classification|Chief Complaint|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|302,311|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|302,311|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|313,325|false|false|false|||Paracentesis
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|313,325|false|false|false|C0034115|Paracentesis|Paracentesis
Event|Event|History of Present Illness|389,396|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|389,396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|389,396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|389,396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|389,399|false|false|false|C0262926|Medical History|history of
Drug|Organic Chemical|History of Present Illness|400,404|false|false|false|C0001962|ethanol|ETOH
Drug|Pharmacologic Substance|History of Present Illness|400,404|false|false|false|C0001962|ethanol|ETOH
Event|Event|History of Present Illness|400,404|false|false|false|||ETOH
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|400,410|false|false|false|C0085762|Alcohol abuse|ETOH abuse
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|405,410|false|false|false|C0013146|Drug abuse|abuse
Event|Event|History of Present Illness|405,410|false|false|false|||abuse
Event|Event|History of Present Illness|405,410|false|false|false|C1546935|Abuse|abuse
Finding|Finding|History of Present Illness|405,410|false|false|false|C0562381|Victim of abuse (finding)|abuse
Event|Event|History of Present Illness|416,424|false|false|false|||presents
Anatomy|Body Location or Region|History of Present Illness|430,439|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|430,450|false|false|false|C0000731|Abdomen distended|abdominal distention
Event|Event|History of Present Illness|440,450|false|false|false|||distention
Finding|Finding|History of Present Illness|440,450|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|440,450|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Sign or Symptom|History of Present Illness|452,461|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|History of Present Illness|457,461|false|false|false|C2598155||pain
Event|Event|History of Present Illness|457,461|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|457,461|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|457,461|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|463,468|false|false|false|||fever
Finding|Finding|History of Present Illness|463,468|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|463,468|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|490,495|false|false|false|||count
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|501,506|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|History of Present Illness|501,506|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|History of Present Illness|501,506|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|History of Present Illness|501,506|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|History of Present Illness|501,506|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|History of Present Illness|501,506|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Finding|Finding|History of Present Illness|501,506|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|History of Present Illness|501,506|false|false|false|C0872387|Procedures on liver|Liver
Event|Event|History of Present Illness|538,546|false|false|false|||admitted
Event|Event|History of Present Illness|555,563|false|false|false|||hospital
Finding|Idea or Concept|History of Present Illness|555,563|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|History of Present Illness|572,576|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|History of Present Illness|577,580|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|586,595|false|false|false|||treatment
Finding|Conceptual Entity|History of Present Illness|586,595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|History of Present Illness|586,595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|History of Present Illness|586,595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|586,595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|History of Present Illness|599,606|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|599,606|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|599,606|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|History of Present Illness|611,615|false|false|false|||work
Event|Occupational Activity|History of Present Illness|611,615|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|History of Present Illness|611,618|false|false|false|C0750430|Work-up|work-up
Disorder|Disease or Syndrome|History of Present Illness|622,641|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|History of Present Illness|632,641|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|History of Present Illness|632,641|false|false|false|||hepatitis
Finding|Finding|History of Present Illness|653,657|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|653,657|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|653,657|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|668,678|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|History of Present Illness|668,678|false|false|false|||diagnostic
Finding|Functional Concept|History of Present Illness|668,678|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|History of Present Illness|668,678|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|History of Present Illness|668,678|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Finding|Functional Concept|History of Present Illness|668,694|false|false|false|C5817574|Combined diagnostic and therapeutic intent|diagnostic and therapeutic
Drug|Organic Chemical|History of Present Illness|683,694|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|History of Present Illness|683,694|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|History of Present Illness|683,694|false|false|false|||therapeutic
Finding|Functional Concept|History of Present Illness|683,694|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|History of Present Illness|683,694|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|683,694|false|false|false|C0087111|Therapeutic procedure|therapeutic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|683,707|false|false|false|C2057774|Therapeutic abdominal paracentesis|therapeutic paracentesis
Event|Event|History of Present Illness|695,707|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|695,707|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|History of Present Illness|717,724|false|false|false|||treated
Disorder|Disease or Syndrome|History of Present Illness|731,734|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|731,734|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|History of Present Illness|731,734|false|false|false|C0077906|urinastatin|UTI
Event|Event|History of Present Illness|731,734|false|false|false|||UTI
Finding|Gene or Genome|History of Present Illness|731,734|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|History of Present Illness|745,755|false|false|false|||discharged
Event|Event|History of Present Illness|756,760|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|756,760|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|756,760|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|756,760|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|765,775|false|false|false|||instructed
Event|Event|History of Present Illness|780,786|false|false|false|||follow
Finding|Functional Concept|History of Present Illness|780,786|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|History of Present Illness|780,786|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|History of Present Illness|780,789|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|History of Present Illness|780,789|false|false|false|C1522577|follow-up|follow-up
Event|Event|History of Present Illness|787,789|false|false|false|||up
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|793,798|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|Liver
Disorder|Disease or Syndrome|History of Present Illness|793,798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Disorder|Neoplastic Process|History of Present Illness|793,798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|Liver
Drug|Organic Chemical|History of Present Illness|793,798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Pharmacologic Substance|History of Present Illness|793,798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Drug|Vitamin|History of Present Illness|793,798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|Liver
Event|Event|History of Present Illness|793,798|false|false|false|||Liver
Finding|Finding|History of Present Illness|793,798|false|false|false|C0577060|Liver problem|Liver
Procedure|Health Care Activity|History of Present Illness|793,798|false|false|false|C0872387|Procedures on liver|Liver
Finding|Intellectual Product|History of Present Illness|811,815|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|History of Present Illness|821,824|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|821,824|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|828,840|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|828,840|false|false|false|C0449450|Presentation|presentation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|845,850|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|History of Present Illness|845,850|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|History of Present Illness|845,850|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|History of Present Illness|845,850|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|History of Present Illness|845,850|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|History of Present Illness|845,850|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|History of Present Illness|845,850|false|false|false|||liver
Finding|Finding|History of Present Illness|845,850|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|History of Present Illness|845,850|false|false|false|C0872387|Procedures on liver|liver
Finding|Body Substance|History of Present Illness|859,866|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|859,866|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|859,866|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|867,877|false|false|false|||complained
Event|Event|History of Present Illness|881,890|false|false|false|||worsening
Finding|Idea or Concept|History of Present Illness|881,890|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|History of Present Illness|891,900|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|891,905|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|901,905|false|false|false|C2598155||pain
Event|Event|History of Present Illness|901,905|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|901,905|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|901,905|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|911,914|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|911,914|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Classification|History of Present Illness|915,920|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|History of Present Illness|915,920|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Event|Event|History of Present Illness|921,927|false|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|921,927|false|false|false|C0015967|Fever|fevers
Finding|Finding|History of Present Illness|928,935|false|false|false|C4534363|At home|at home
Event|Event|History of Present Illness|931,935|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|931,935|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|931,935|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|931,935|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|942,949|false|false|false|||labwork
Event|Event|History of Present Illness|959,970|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|959,970|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|1024,1032|false|false|false|||admitted
Event|Occupational Activity|History of Present Illness|1037,1041|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|History of Present Illness|1037,1044|false|false|false|C0750430|Work-up|work-up
Event|Event|History of Present Illness|1048,1053|false|false|false|||fever
Finding|Finding|History of Present Illness|1048,1053|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1048,1053|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1079,1088|false|false|false|||treatment
Finding|Conceptual Entity|History of Present Illness|1079,1088|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|History of Present Illness|1079,1088|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|History of Present Illness|1079,1088|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1079,1088|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|History of Present Illness|1103,1110|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|1103,1110|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|1103,1110|false|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Organic Chemical|Past Medical History|1138,1145|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Drug|Pharmacologic Substance|Past Medical History|1138,1145|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Finding|Intellectual Product|Past Medical History|1138,1145|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|Alcohol
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1138,1151|false|false|false|C0085762|Alcohol abuse|Alcohol abuse
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1146,1151|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Past Medical History|1146,1151|false|false|false|||abuse
Event|Event|Past Medical History|1146,1151|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Past Medical History|1146,1151|false|false|false|C0562381|Victim of abuse (finding)|abuse
Finding|Intellectual Product|Past Medical History|1154,1161|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Past Medical History|1154,1161|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|Past Medical History|1154,1171|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|Past Medical History|1162,1171|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Past Medical History|1167,1171|false|false|false|C2598155||pain
Event|Event|Past Medical History|1167,1171|false|false|false|||pain
Finding|Functional Concept|Past Medical History|1167,1171|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Past Medical History|1167,1171|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1210,1216|false|false|false|C0006141|Breast|Breast
Disorder|Neoplastic Process|Family Medical History|1210,1216|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|Breast
Event|Event|Family Medical History|1210,1216|false|false|false|||Breast
Finding|Finding|Family Medical History|1210,1216|false|false|false|C0567499|Breast problem|Breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1210,1216|false|false|false|C0191838|Procedures on breast|Breast
Disorder|Neoplastic Process|Family Medical History|1210,1223|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|Breast cancer
Disorder|Neoplastic Process|Family Medical History|1217,1223|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1217,1223|false|false|false|||cancer
Finding|Idea or Concept|Family Medical History|1227,1233|true|false|false|C1546508|Relationship - Mother|mother
Attribute|Clinical Attribute|Family Medical History|1234,1237|true|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|1234,1237|true|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|1234,1237|true|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|1234,1237|true|false|false|||age
Disorder|Disease or Syndrome|Family Medical History|1246,1249|true|false|false|C0021390;C0022104|Inflammatory Bowel Diseases;Irritable Bowel Syndrome|IBD
Drug|Organic Chemical|Family Medical History|1246,1249|true|false|false|C0123047|ibudilast|IBD
Drug|Pharmacologic Substance|Family Medical History|1246,1249|true|false|false|C0123047|ibudilast|IBD
Event|Event|Family Medical History|1246,1249|true|false|false|||IBD
Finding|Gene or Genome|Family Medical History|1246,1249|true|false|false|C5780974|ACAD8 wt Allele|IBD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1251,1256|true|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|1251,1256|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|1251,1256|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|1251,1256|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|1251,1256|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|1251,1256|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Family Medical History|1251,1256|true|false|false|||liver
Finding|Finding|Family Medical History|1251,1256|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|1251,1256|true|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|1251,1264|true|false|false|C0085605|Liver Failure|liver failure
Event|Event|Family Medical History|1257,1264|true|false|false|||failure
Finding|Functional Concept|Family Medical History|1257,1264|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Family Medical History|1257,1264|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Family Medical History|1257,1264|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Family Medical History|1277,1286|false|false|false|||relatives
Disorder|Mental or Behavioral Dysfunction|Family Medical History|1292,1302|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcoholism
Event|Event|Family Medical History|1292,1302|false|false|false|||alcoholism
Event|Event|General Exam|1356,1359|false|false|false|||GEN
Finding|Classification|General Exam|1356,1359|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|1356,1359|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Event|Event|General Exam|1368,1376|false|false|false|||pleasant
Finding|Mental Process|General Exam|1368,1376|false|false|false|C2987187|Pleasant|pleasant
Event|Event|General Exam|1378,1389|false|false|false|||appropriate
Finding|Finding|General Exam|1391,1395|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1396,1405|false|false|false|||appearing
Anatomy|Body Location or Region|General Exam|1408,1413|false|false|false|C1512338|HEENT|HEENT
Disorder|Disease or Syndrome|General Exam|1418,1434|true|false|false|C1112303|Facial wasting|temporal wasting
Finding|Finding|General Exam|1418,1434|true|false|false|C2029785|Temporal wasting|temporal wasting
Disorder|Disease or Syndrome|General Exam|1427,1434|true|false|false|C0235394|Wasting|wasting
Event|Event|General Exam|1427,1434|true|false|false|||wasting
Finding|Sign or Symptom|General Exam|1427,1434|true|false|false|C0006625|Cachexia|wasting
Event|Event|General Exam|1436,1439|true|false|false|||JVD
Finding|Finding|General Exam|1436,1439|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|General Exam|1454,1458|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|1454,1458|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|1454,1458|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|General Exam|1454,1464|true|false|false|C0226542;C4266538|Neck>Neck veins;Structure of vein of neck|neck veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|1459,1464|true|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|1459,1464|true|false|false|C0398102|Procedure on vein|veins
Event|Activity|General Exam|1465,1469|true|false|false|C1708059|Fill|fill
Finding|Idea or Concept|General Exam|1476,1481|false|false|false|C1552828|Table Frame - above|above
Event|Event|General Exam|1489,1492|true|false|false|||RRR
Event|Event|General Exam|1497,1500|true|false|false|||MRG
Finding|Gene or Genome|General Exam|1497,1500|true|false|false|C1422304|MAS1L gene|MRG
Event|Event|General Exam|1503,1507|true|false|false|||PULM
Procedure|Health Care Activity|General Exam|1503,1507|true|false|false|C1315068|Pulmonary ventilator management|PULM
Drug|Organic Chemical|General Exam|1509,1513|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|1509,1513|false|false|false|||CTAB
Event|Event|General Exam|1518,1527|false|false|false|||decreased
Finding|Finding|General Exam|1518,1527|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Anatomy|Body Location or Region|General Exam|1536,1540|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|1536,1540|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|1536,1540|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1536,1540|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|1536,1540|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|1536,1540|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Location or Region|General Exam|1544,1547|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|1544,1547|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|1544,1547|false|false|false|||ABD
Event|Event|General Exam|1549,1558|false|false|false|||Distended
Finding|Finding|General Exam|1549,1558|false|false|false|C0700124|Dilated|Distended
Event|Event|General Exam|1580,1586|false|false|false|||tender
Event|Event|General Exam|1590,1599|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|1590,1599|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|1617,1627|false|false|false|||flatulence
Finding|Sign or Symptom|General Exam|1617,1627|false|false|false|C0016204|Flatulence|flatulence
Anatomy|Body Part, Organ, or Organ Component|General Exam|1631,1636|false|false|false|C0015385|Limb structure|LIMBS
Attribute|Clinical Attribute|General Exam|1641,1646|false|false|false|C1717255||edema
Event|Event|General Exam|1641,1646|false|false|false|||edema
Finding|Pathologic Function|General Exam|1641,1646|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|1654,1657|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|General Exam|1654,1657|false|false|false|C0023595|Lewis Blood-Group System|LEs
Anatomy|Body Location or Region|General Exam|1661,1665|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|1661,1665|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|1661,1665|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|1661,1665|false|false|false|C0562271|Examination of knee joint|knee
Drug|Food|General Exam|1682,1688|false|false|false|C5890763||pulses
Event|Event|General Exam|1682,1688|false|false|false|||pulses
Finding|Physiologic Function|General Exam|1682,1688|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|1682,1688|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|1717,1726|true|false|false|||asterixis
Finding|Sign or Symptom|General Exam|1717,1726|true|false|false|C0232766|Asterixis|asterixis
Finding|Finding|General Exam|1728,1737|true|false|false|C4036115|Very mild|very mild
Finding|Intellectual Product|General Exam|1733,1737|true|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|General Exam|1738,1745|true|false|false|||general
Finding|Classification|General Exam|1738,1745|true|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|General Exam|1738,1745|true|false|false|C3812897|General medical service|general
Event|Event|General Exam|1746,1752|true|false|false|||tremor
Finding|Sign or Symptom|General Exam|1746,1752|true|false|false|C0040822|Tremor|tremor
Event|Event|General Exam|1775,1779|false|false|false|||Labs
Lab|Laboratory or Test Result|General Exam|1775,1779|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Finding|General Exam|1780,1792|false|false|false|C4533677|at admission|at Admission
Event|Event|General Exam|1783,1792|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|1783,1792|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Disorder|Disease or Syndrome|General Exam|1807,1812|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1807,1812|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1807,1812|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1813,1816|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1824,1827|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1824,1827|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1824,1827|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1834,1837|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1834,1837|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1834,1837|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1834,1837|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1843,1846|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1843,1846|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1853,1856|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|1853,1856|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|1853,1856|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1853,1856|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1853,1856|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1862,1865|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1862,1865|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|1862,1865|false|false|false|||MCH
Finding|Gene or Genome|General Exam|1862,1865|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1862,1865|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1862,1865|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|1872,1876|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|1892,1895|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|1912,1917|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1912,1917|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1912,1917|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|1936,1942|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|1946,1951|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|1946,1951|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|1946,1951|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|1954,1957|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|1954,1957|false|false|false|||Eos
Finding|Gene or Genome|General Exam|1954,1957|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|1993,1998|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1993,1998|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1993,1998|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|2015,2020|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2015,2020|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2015,2020|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Inorganic Chemical|General Exam|2060,2064|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2060,2064|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2060,2064|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2089,2094|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2089,2094|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2095,2098|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2095,2098|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2095,2098|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|2095,2098|false|false|false|||ALT
Finding|Gene or Genome|General Exam|2095,2098|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2095,2098|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2095,2098|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2095,2098|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|2103,2106|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2103,2106|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2103,2106|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2103,2106|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2103,2106|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|2103,2106|false|false|false|||AST
Finding|Gene or Genome|General Exam|2103,2106|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2115,2118|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|2115,2118|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|General Exam|2115,2118|false|false|false|||LDH
Finding|Finding|General Exam|2115,2118|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|2115,2118|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|2126,2133|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|2126,2133|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|2164,2169|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2164,2169|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2164,2169|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2164,2177|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|2170,2177|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|2170,2177|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|2170,2177|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|2170,2177|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|2170,2177|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|2170,2177|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|2170,2177|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|2183,2190|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2183,2190|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2183,2190|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2183,2190|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2183,2190|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2183,2190|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2183,2190|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2183,2190|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|2224,2229|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2224,2229|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2224,2229|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2224,2237|false|false|false|C0855900|Blood ethanol|BLOOD Ethanol
Disorder|Injury or Poisoning|General Exam|2230,2237|false|false|false|C0161679|Toxic effect of ethyl alcohol|Ethanol
Drug|Organic Chemical|General Exam|2230,2237|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Drug|Pharmacologic Substance|General Exam|2230,2237|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Event|Event|General Exam|2230,2237|false|false|false|||Ethanol
Procedure|Laboratory Procedure|General Exam|2230,2237|false|false|false|C0202304|Ethanol measurement|Ethanol
Event|Event|General Exam|2238,2241|false|false|false|||NEG
Finding|Finding|General Exam|2238,2241|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|2250,2253|false|false|false|||NEG
Finding|Finding|General Exam|2250,2253|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|2255,2259|false|false|false|||Labs
Lab|Laboratory or Test Result|General Exam|2255,2259|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|General Exam|2263,2272|false|false|false|||Discharge
Finding|Body Substance|General Exam|2263,2272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|2263,2272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|2263,2272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|2263,2272|false|false|false|C0030685|Patient Discharge|Discharge
Disorder|Disease or Syndrome|General Exam|2287,2292|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2287,2292|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2287,2292|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2293,2296|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2303,2306|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2303,2306|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2303,2306|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2313,2316|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2313,2316|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2313,2316|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2313,2316|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2323,2326|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2323,2326|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2334,2337|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2334,2337|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2334,2337|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2334,2337|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2334,2337|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2343,2346|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2343,2346|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2343,2346|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2343,2346|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2343,2346|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2343,2346|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2353,2357|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2353,2357|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2372,2375|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2392,2397|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2392,2397|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2392,2397|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2402,2405|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|2402,2405|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|2402,2405|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2428,2433|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2428,2433|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2428,2433|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2428,2441|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2428,2441|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2428,2441|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2434,2441|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2434,2441|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2434,2441|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2434,2441|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2434,2441|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2434,2441|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|2513,2518|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2513,2518|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2513,2518|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2519,2522|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2519,2522|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2519,2522|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|2519,2522|false|false|false|||ALT
Finding|Gene or Genome|General Exam|2519,2522|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2519,2522|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2519,2522|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2519,2522|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|2526,2529|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2526,2529|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2526,2529|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2526,2529|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2526,2529|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|2526,2529|false|false|false|||AST
Finding|Gene or Genome|General Exam|2526,2529|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2548,2555|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|2548,2555|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|2587,2592|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2587,2592|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2587,2592|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2587,2600|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|2593,2600|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|2593,2600|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|2593,2600|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|2593,2600|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|2593,2600|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|2593,2600|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|2593,2600|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|2606,2613|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2606,2613|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2606,2613|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2606,2613|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2606,2613|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2606,2613|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2606,2613|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2606,2613|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Conceptual Entity|General Exam|2638,2643|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|General Exam|2638,2643|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|General Exam|2638,2643|false|false|false|C0085672|Microbiology procedure|Micro
Event|Event|General Exam|2644,2648|false|false|false|||Data
Finding|Idea or Concept|General Exam|2644,2648|false|false|false|C1511726|Data|Data
Anatomy|Body Location or Region|General Exam|2655,2665|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|2655,2665|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|2655,2671|true|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|2655,2671|true|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|2655,2682|false|false|false|C2020989|peritoneal fluid Gram stain|PERITONEAL FLUID GRAM STAIN
Drug|Substance|General Exam|2666,2671|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|2666,2671|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|2666,2671|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2672,2682|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|2672,2682|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|2672,2682|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2677,2682|true|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|2677,2682|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|2677,2682|true|false|false|C0487602|Staining method|STAIN
Event|Event|General Exam|2684,2692|false|false|false|||negative
Finding|Classification|General Exam|2684,2692|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2684,2692|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2684,2692|false|false|false|C5237010|Expression Negative|negative
Drug|Substance|General Exam|2694,2699|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|2694,2699|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|2694,2699|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|2701,2708|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|2701,2708|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|2701,2708|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|2701,2708|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|2701,2708|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|2709,2716|false|false|false|||PENDING
Finding|Idea or Concept|General Exam|2709,2716|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|PENDING
Procedure|Laboratory Procedure|General Exam|2718,2735|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|2728,2735|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|2728,2735|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|2728,2735|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|2728,2735|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|2728,2735|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|2737,2745|false|false|false|||negative
Finding|Classification|General Exam|2737,2745|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2737,2745|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2737,2745|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|General Exam|2750,2755|false|false|false|C0015733|Feces|STOOL
Drug|Amino Acid, Peptide, or Protein|General Exam|2756,2783|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Biologically Active Substance|General Exam|2756,2783|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Hazardous or Poisonous Substance|General Exam|2756,2783|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Amino Acid, Peptide, or Protein|General Exam|2756,2785|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|General Exam|2756,2785|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Hazardous or Poisonous Substance|General Exam|2756,2785|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|General Exam|2778,2783|false|false|false|C0040549|Toxin|TOXIN
Drug|Hazardous or Poisonous Substance|General Exam|2778,2783|false|false|false|C0040549|Toxin|TOXIN
Event|Event|General Exam|2778,2783|false|false|false|||TOXIN
Event|Event|General Exam|2784,2785|false|false|false|||A
Anatomy|Body Location or Region|General Exam|2791,2795|false|false|false|C4318744|Test - temporal region|TEST
Event|Event|General Exam|2791,2795|false|false|false|||TEST
Finding|Functional Concept|General Exam|2791,2795|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Finding|Intellectual Product|General Exam|2791,2795|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Lab|Laboratory or Test Result|General Exam|2791,2795|false|false|false|C0456984|Test Result|TEST
Procedure|Laboratory Procedure|General Exam|2791,2795|false|false|false|C0022885|Laboratory Procedures|TEST
Event|Event|General Exam|2797,2805|false|false|false|||negative
Finding|Classification|General Exam|2797,2805|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2797,2805|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2797,2805|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|General Exam|2810,2815|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2810,2815|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2810,2815|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|General Exam|2816,2821|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2816,2821|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2816,2821|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|2816,2829|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|2822,2829|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|2822,2829|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|2822,2829|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|2822,2829|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|2822,2829|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|2831,2839|false|false|false|||negative
Finding|Classification|General Exam|2831,2839|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2831,2839|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2831,2839|false|false|false|C5237010|Expression Negative|negative
Drug|Biomedical or Dental Material|General Exam|2844,2848|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|SWAB
Drug|Substance|General Exam|2844,2848|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|SWAB
Event|Event|General Exam|2844,2848|false|false|false|||SWAB
Procedure|Diagnostic Procedure|General Exam|2844,2848|false|false|false|C0563454|Taking of swab|SWAB
Drug|Amino Acid, Peptide, or Protein|General Exam|2853,2863|false|true|false|C0042313|vancomycin|VANCOMYCIN
Drug|Antibiotic|General Exam|2853,2863|false|true|false|C0042313|vancomycin|VANCOMYCIN
Event|Event|General Exam|2853,2863|false|false|false|||VANCOMYCIN
Procedure|Laboratory Procedure|General Exam|2853,2863|false|true|false|C0489941|Vancomycin measurement|VANCOMYCIN
Finding|Functional Concept|General Exam|2864,2873|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|RESISTANT
Finding|Idea or Concept|General Exam|2864,2873|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|RESISTANT
Lab|Laboratory or Test Result|General Exam|2864,2873|false|false|false|C2827757|Antimicrobial Resistance Result|RESISTANT
Event|Event|General Exam|2889,2897|false|false|false|||negative
Finding|Classification|General Exam|2889,2897|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2889,2897|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2889,2897|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|General Exam|2902,2907|false|false|false|C0015733|Feces|STOOL
Drug|Amino Acid, Peptide, or Protein|General Exam|2908,2935|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Biologically Active Substance|General Exam|2908,2935|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Hazardous or Poisonous Substance|General Exam|2908,2935|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Amino Acid, Peptide, or Protein|General Exam|2908,2937|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|General Exam|2908,2937|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Hazardous or Poisonous Substance|General Exam|2908,2937|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|General Exam|2930,2935|false|false|false|C0040549|Toxin|TOXIN
Drug|Hazardous or Poisonous Substance|General Exam|2930,2935|false|false|false|C0040549|Toxin|TOXIN
Event|Event|General Exam|2930,2935|false|false|false|||TOXIN
Event|Event|General Exam|2936,2937|false|false|false|||A
Anatomy|Body Location or Region|General Exam|2943,2947|false|false|false|C4318744|Test - temporal region|TEST
Event|Event|General Exam|2943,2947|false|false|false|||TEST
Finding|Functional Concept|General Exam|2943,2947|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Finding|Intellectual Product|General Exam|2943,2947|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Lab|Laboratory or Test Result|General Exam|2943,2947|false|false|false|C0456984|Test Result|TEST
Procedure|Laboratory Procedure|General Exam|2943,2947|false|false|false|C0022885|Laboratory Procedures|TEST
Event|Event|General Exam|2949,2957|false|false|false|||negative
Finding|Classification|General Exam|2949,2957|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|2949,2957|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|2949,2957|false|false|false|C5237010|Expression Negative|negative
Drug|Substance|General Exam|2962,2967|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|2962,2967|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|2962,2967|false|false|false|C1546638|Fluid Specimen Code|FLUID
Event|Event|General Exam|2968,2976|false|false|false|||RECEIVED
Finding|Body Substance|General Exam|2977,2985|false|false|false|C0005768|In Blood|IN BLOOD
Disorder|Disease or Syndrome|General Exam|2980,2985|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2980,2985|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2980,2985|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2980,2993|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|2986,2993|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|2986,2993|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|2986,2993|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|2986,2993|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|2986,2993|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|2994,3001|false|false|false|||BOTTLES
Drug|Substance|General Exam|3003,3008|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|General Exam|3003,3008|false|false|false|||Fluid
Finding|Intellectual Product|General Exam|3003,3008|false|false|false|C1546638|Fluid Specimen Code|Fluid
Drug|Biomedical or Dental Material|General Exam|3009,3016|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|3009,3016|false|false|false|||Culture
Finding|Functional Concept|General Exam|3009,3016|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|3009,3016|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|3009,3016|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|General Exam|3029,3037|false|false|false|||negative
Finding|Classification|General Exam|3029,3037|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|3029,3037|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|3029,3037|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Location or Region|General Exam|3042,3052|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|3042,3052|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|3042,3058|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|3042,3058|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|3042,3069|false|false|false|C2020989|peritoneal fluid Gram stain|PERITONEAL FLUID GRAM STAIN
Drug|Substance|General Exam|3053,3058|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|3053,3058|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|3053,3058|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3059,3069|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|3059,3069|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|3059,3069|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3064,3069|false|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|3064,3069|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|3064,3069|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|3070,3075|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Drug|Substance|General Exam|3077,3082|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|3077,3082|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|3077,3082|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|3084,3091|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3084,3091|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3084,3091|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3084,3091|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3084,3091|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|3092,3097|false|false|false|||FINAL
Finding|Idea or Concept|General Exam|3092,3097|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Procedure|Laboratory Procedure|General Exam|3099,3116|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|3109,3116|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3109,3116|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3109,3116|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3109,3116|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3109,3116|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|3118,3126|false|false|false|||negative
Finding|Classification|General Exam|3118,3126|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|3118,3126|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|3118,3126|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|General Exam|3131,3136|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3131,3136|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3131,3144|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|3137,3144|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3137,3144|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3137,3144|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3137,3144|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3137,3144|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Procedure|Laboratory Procedure|General Exam|3137,3150|false|false|false|C0200949|Blood culture|CULTURE Blood
Disorder|Disease or Syndrome|General Exam|3145,3150|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|3145,3150|false|false|false|||Blood
Finding|Body Substance|General Exam|3145,3150|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|3145,3158|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|3151,3158|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|3151,3158|false|false|false|||Culture
Finding|Functional Concept|General Exam|3151,3158|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|3151,3158|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|3151,3158|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|General Exam|3160,3167|false|false|false|||Routine
Finding|Idea or Concept|General Exam|3160,3167|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|General Exam|3160,3167|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|General Exam|3160,3167|false|false|false|C1979801|Routine coag|Routine
Event|Event|General Exam|3170,3178|false|false|false|||negative
Finding|Classification|General Exam|3170,3178|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|3170,3178|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|3170,3178|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|General Exam|3184,3189|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3184,3189|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3184,3197|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|3190,3197|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3190,3197|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3190,3197|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3190,3197|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3190,3197|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Procedure|Laboratory Procedure|General Exam|3190,3203|false|false|false|C0200949|Blood culture|CULTURE Blood
Disorder|Disease or Syndrome|General Exam|3198,3203|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|3198,3203|false|false|false|||Blood
Finding|Body Substance|General Exam|3198,3203|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|3198,3211|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|3204,3211|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|3204,3211|false|false|false|||Culture
Finding|Functional Concept|General Exam|3204,3211|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|3204,3211|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|3204,3211|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Event|Event|General Exam|3214,3221|false|false|false|||Routine
Finding|Idea or Concept|General Exam|3214,3221|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|General Exam|3214,3221|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|General Exam|3214,3221|false|false|false|C1979801|Routine coag|Routine
Event|Event|General Exam|3222,3230|false|false|false|||negative
Finding|Classification|General Exam|3222,3230|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|3222,3230|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|3222,3230|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|General Exam|3236,3241|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|3236,3241|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|3236,3241|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|General Exam|3242,3247|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|3242,3247|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|3242,3247|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|3242,3255|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|3248,3255|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3248,3255|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3248,3255|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3248,3255|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3248,3255|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|General Exam|3256,3261|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Disorder|Cell or Molecular Dysfunction|General Exam|3268,3276|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Event|Event|General Exam|3268,3276|false|false|false|||POSITIVE
Finding|Classification|General Exam|3268,3276|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|General Exam|3268,3276|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Event|Event|General Exam|3278,3286|false|false|false|||BACTERIA
Finding|Functional Concept|General Exam|3278,3286|false|false|false|C1510439|bacteria aspects|BACTERIA
Event|Event|General Exam|3288,3297|false|false|false|||INPATIENT
Finding|Idea or Concept|General Exam|3288,3297|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|INPATIENT
Procedure|Health Care Activity|General Exam|3288,3297|false|false|false|C1555324|inpatient encounter|INPATIENT
Drug|Substance|General Exam|3303,3308|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|3303,3308|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|3303,3308|false|false|false|C1546638|Fluid Specimen Code|FLUID
Event|Event|General Exam|3309,3317|false|false|false|||RECEIVED
Finding|Body Substance|General Exam|3318,3326|false|false|false|C0005768|In Blood|IN BLOOD
Disorder|Disease or Syndrome|General Exam|3321,3326|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3321,3326|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3321,3326|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3321,3334|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|3327,3334|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|3327,3334|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|3327,3334|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|3327,3334|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|3327,3334|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|3335,3342|false|false|false|||BOTTLES
Event|Event|General Exam|3344,3352|false|false|false|||negative
Finding|Classification|General Exam|3344,3352|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|3344,3352|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|3344,3352|false|false|false|C5237010|Expression Negative|negative
Event|Event|General Exam|3354,3361|false|false|false|||Imaging
Finding|Finding|General Exam|3354,3361|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|3354,3361|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Drug|Amino Acid, Peptide, or Protein|General Exam|3372,3375|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|3372,3375|false|false|false|||CTA
Finding|Gene or Genome|General Exam|3372,3375|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|3372,3375|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|General Exam|3389,3397|true|false|false|||evidence
Finding|Idea or Concept|General Exam|3389,3397|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|3389,3400|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|General Exam|3401,3410|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|3401,3410|true|false|false|C2707265||pulmonary
Finding|Finding|General Exam|3401,3410|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|3401,3419|true|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|General Exam|3411,3419|true|false|false|||embolism
Finding|Finding|General Exam|3411,3419|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|General Exam|3411,3419|true|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Intellectual Product|General Exam|3425,3431|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|General Exam|3432,3443|false|false|false|||atelectasis
Finding|Pathologic Function|General Exam|3432,3443|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Functional Concept|General Exam|3451,3456|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|3451,3461|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|General Exam|3451,3466|false|false|false|C0225708|Structure of base of right lung|right lung base
Anatomy|Body Location or Region|General Exam|3457,3461|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3457,3461|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3457,3461|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3457,3461|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3457,3466|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|General Exam|3462,3466|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|3462,3466|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|3462,3466|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3462,3466|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|3462,3466|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|3462,3466|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Finding|General Exam|3472,3480|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|3472,3480|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|General Exam|3481,3486|false|false|false|||right
Finding|Functional Concept|General Exam|3481,3486|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|General Exam|3497,3501|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|General Exam|3502,3509|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|3502,3509|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|3502,3519|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|General Exam|3510,3519|false|false|false|||effusions
Finding|Pathologic Function|General Exam|3510,3519|false|false|false|C0013687|effusion|effusions
Event|Event|General Exam|3521,3530|false|false|false|||unchanged
Finding|Finding|General Exam|3521,3530|false|false|false|C0442739||unchanged
Event|Event|General Exam|3534,3538|false|false|false|||CTAP
Event|Event|General Exam|3549,3561|false|false|false|||Hepatomegaly
Finding|Finding|General Exam|3549,3561|false|false|false|C0019209|Hepatomegaly|Hepatomegaly
Finding|Gene or Genome|General Exam|3566,3571|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|General Exam|3572,3579|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|3572,3579|false|false|false|||ascites
Finding|Pathologic Function|General Exam|3572,3579|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|General Exam|3580,3590|false|false|false|||consistent
Finding|Idea or Concept|General Exam|3580,3590|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|3580,3595|false|false|false|C0332290|Consistent with|consistent with
Event|Event|General Exam|3603,3610|false|false|false|||history
Finding|Conceptual Entity|General Exam|3603,3610|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|3603,3610|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|3603,3610|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Anatomy|Body Part, Organ, or Organ Component|General Exam|3615,3620|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|3615,3620|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|3615,3620|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|3615,3620|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|3615,3620|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|3615,3620|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|3615,3620|false|false|false|||liver
Finding|Finding|General Exam|3615,3620|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|3615,3620|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|General Exam|3622,3629|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|3622,3629|false|false|false|||disease
Event|Event|General Exam|3634,3642|true|false|false|||evidence
Finding|Idea or Concept|General Exam|3634,3642|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|3634,3645|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Location or Region|General Exam|3646,3652|true|false|false|C0205054|Hepatic|portal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3653,3659|true|false|false|C0042449|Veins|venous
Finding|Finding|General Exam|3653,3670|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|General Exam|3653,3670|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|General Exam|3660,3670|true|false|false|||thrombosis
Finding|Pathologic Function|General Exam|3660,3670|true|false|false|C0040053|Thrombosis|thrombosis
Event|Event|General Exam|3671,3681|true|false|false|||suggesting
Attribute|Clinical Attribute|General Exam|3692,3700|false|false|false|C2926606||findings
Event|Event|General Exam|3692,3700|false|false|false|||findings
Finding|Functional Concept|General Exam|3692,3700|false|false|false|C2607943|findings aspects|findings
Event|Event|General Exam|3714,3724|false|false|false|||ultrasound
Finding|Functional Concept|General Exam|3714,3724|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|3714,3724|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|3714,3724|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|General Exam|3734,3742|false|false|false|||resulted
Attribute|Clinical Attribute|General Exam|3766,3778|false|false|false|C3827727|Undetectable|undetectable
Phenomenon|Natural Phenomenon or Process|General Exam|3779,3783|false|false|false|C0806140|Flow|flow
Finding|Finding|General Exam|3790,3798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|3790,3798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|General Exam|3799,3804|false|false|false|||right
Finding|Functional Concept|General Exam|3799,3804|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|General Exam|3815,3819|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|General Exam|3820,3827|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|3820,3827|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|3820,3837|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|General Exam|3828,3837|false|false|false|||effusions
Finding|Pathologic Function|General Exam|3828,3837|false|false|false|C0013687|effusion|effusions
Event|Event|General Exam|3839,3848|false|false|false|||increased
Finding|Functional Concept|General Exam|3857,3862|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|General Exam|3869,3874|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Pathologic Function|General Exam|3875,3894|false|false|false|C4049574|Basilar atelectasis|basilar atelectasis
Event|Event|General Exam|3883,3894|false|false|false|||atelectasis
Finding|Pathologic Function|General Exam|3883,3894|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Functional Concept|General Exam|3900,3908|false|false|false|C0559956;C1299987|Replaced by;Replacement|Replaced
Finding|Functional Concept|General Exam|3909,3914|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|3909,3929|false|false|false|C0226302;C1305708|Structure of right branch of hepatic artery|right hepatic artery
Anatomy|Body Location or Region|General Exam|3915,3922|false|false|false|C0205054|Hepatic|hepatic
Anatomy|Body Part, Organ, or Organ Component|General Exam|3915,3929|false|false|false|C0019145;C4037987|Abdomen>Hepatic artery;Hepatic artery|hepatic artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|3923,3929|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|3923,3929|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|General Exam|3930,3937|false|false|false|||arising
Disorder|Disease or Syndrome|General Exam|3947,3950|false|false|false|C0026847;C4024957;C5890956|Minor Salivary Gland Sclerosing Microcystic Adenocarcinoma;Proximal spinal muscular atrophy;Spinal Muscular Atrophy|SMA
Disorder|Neoplastic Process|General Exam|3947,3950|false|false|false|C0026847;C4024957;C5890956|Minor Salivary Gland Sclerosing Microcystic Adenocarcinoma;Proximal spinal muscular atrophy;Spinal Muscular Atrophy|SMA
Drug|Amino Acid, Peptide, or Protein|General Exam|3947,3950|false|false|false|C1700794|SNRPF protein, human|SMA
Drug|Immunologic Factor|General Exam|3947,3950|false|false|false|C1700794|SNRPF protein, human|SMA
Event|Event|General Exam|3947,3950|false|false|false|||SMA
Finding|Gene or Genome|General Exam|3947,3950|false|false|false|C1420257;C4284041|SMN1 gene;SMN1 wt Allele|SMA
Anatomy|Body Part, Organ, or Organ Component|General Exam|3976,3984|false|false|false|C0003842|Arteries|arterial
Anatomy|Body Part, Organ, or Organ Component|General Exam|3989,3995|false|false|false|C0042449|Veins|venous
Anatomy|Anatomical Structure|General Exam|3996,4003|false|false|false|C0700276|Anatomical structure|anatomy
Finding|Finding|Hospital Course|4055,4061|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|4055,4061|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|4062,4081|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|4072,4081|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|Hospital Course|4072,4081|false|false|false|||hepatitis
Disorder|Disease or Syndrome|Hospital Course|4097,4104|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|4097,4104|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|4097,4104|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|Hospital Course|4112,4120|false|false|false|||admitted
Finding|Finding|Hospital Course|4126,4129|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|4126,4129|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Classification|Hospital Course|4130,4135|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Hospital Course|4130,4135|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Event|Event|Hospital Course|4136,4142|false|false|false|||fevers
Finding|Sign or Symptom|Hospital Course|4136,4142|false|false|false|C0015967|Fever|fevers
Event|Event|Hospital Course|4144,4148|false|false|false|||high
Finding|Finding|Hospital Course|4144,4148|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|4144,4148|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|4144,4148|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Anatomy|Body Location or Region|Hospital Course|4167,4176|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|4167,4181|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|4177,4181|false|false|false|C2598155||pain
Event|Event|Hospital Course|4177,4181|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4177,4181|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4177,4181|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|4187,4194|false|false|false|C0003962|Ascites|ASCITES
Event|Event|Hospital Course|4187,4194|false|false|false|||ASCITES
Finding|Pathologic Function|Hospital Course|4187,4194|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Anatomy|Body Location or Region|Hospital Course|4195,4198|false|false|false|C3495964|area LC of Bonin|ALC
Finding|Gene or Genome|Hospital Course|4195,4198|false|false|false|C1424945|ALLC gene|ALC
Procedure|Laboratory Procedure|Hospital Course|4195,4198|false|false|false|C3811058|Absolute Blood Lymphocyte Count|ALC
Disorder|Disease or Syndrome|Hospital Course|4199,4208|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|HEPATITIS
Disorder|Disease or Syndrome|Hospital Course|4209,4221|false|false|false|C0023518|Leukocytosis|LEUKOCYTOSIS
Event|Event|Hospital Course|4209,4221|false|false|false|||LEUKOCYTOSIS
Finding|Finding|Hospital Course|4209,4221|false|false|false|C0750426|Blood leukocyte number above reference range|LEUKOCYTOSIS
Finding|Body Substance|Hospital Course|4223,4230|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4223,4230|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4223,4230|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|4236,4247|false|false|false|C0015695;C2711227|Fatty Liver;Steatohepatitis|fatty liver
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4242,4247|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|4242,4247|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|4242,4247|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|4242,4247|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|4242,4247|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|4242,4247|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|4242,4247|false|false|false|||liver
Finding|Finding|Hospital Course|4242,4247|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|4242,4247|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Hospital Course|4253,4260|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|4253,4260|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|4253,4260|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|Hospital Course|4264,4271|false|false|false|||setting
Finding|Mental Process|Hospital Course|4264,4271|false|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|4285,4293|false|false|false|||drinking
Finding|Individual Behavior|Hospital Course|4285,4293|false|false|false|C0001948;C0684271|Alcohol consumption;Drinking (function)|drinking
Finding|Organism Function|Hospital Course|4285,4293|false|false|false|C0001948;C0684271|Alcohol consumption;Drinking (function)|drinking
Event|Event|Hospital Course|4294,4301|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|4294,4301|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4294,4301|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|4294,4301|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Anatomy|Body Space or Junction|Hospital Course|4306,4309|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|Hospital Course|4306,4309|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4306,4309|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|Hospital Course|4306,4309|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|Hospital Course|4306,4309|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|Hospital Course|4306,4309|false|false|false|||AST
Finding|Gene or Genome|Hospital Course|4306,4309|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|Hospital Course|4310,4313|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4310,4313|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|Hospital Course|4310,4313|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|Hospital Course|4310,4313|false|false|false|||ALT
Finding|Gene or Genome|Hospital Course|4310,4313|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|Hospital Course|4310,4313|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|Hospital Course|4310,4313|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4310,4313|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Event|Event|Hospital Course|4315,4324|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4315,4324|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|Hospital Course|4342,4350|false|false|false|||function
Finding|Finding|Hospital Course|4342,4350|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|4342,4350|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|4342,4350|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|4342,4350|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Hospital Course|4354,4363|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4354,4363|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|4375,4382|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4375,4382|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4375,4382|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|4389,4401|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4389,4401|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Hospital Course|4413,4415|false|false|false|||4L
Event|Event|Hospital Course|4420,4427|false|false|false|||removed
Anatomy|Body Location or Region|Hospital Course|4430,4440|true|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|Hospital Course|4430,4440|true|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Finding|Body Substance|Hospital Course|4430,4446|true|false|false|C0003964|Peritoneal fluid (substance)|peritoneal fluid
Procedure|Laboratory Procedure|Hospital Course|4430,4446|true|false|false|C2053903|Peritoneal fluid analysis|peritoneal fluid
Drug|Substance|Hospital Course|4441,4446|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Hospital Course|4441,4446|true|false|false|||fluid
Finding|Intellectual Product|Hospital Course|4441,4446|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Hospital Course|4451,4459|false|false|false|||negative
Finding|Classification|Hospital Course|4451,4459|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|4451,4459|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|4451,4459|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|4451,4463|false|false|false|C0205160|Negative|negative for
Attribute|Clinical Attribute|Hospital Course|4464,4467|true|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4464,4467|true|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|4464,4467|true|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|4464,4467|true|false|false|||SBP
Finding|Gene or Genome|Hospital Course|4464,4467|true|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|4464,4467|true|false|false|C1306620|Systolic blood pressure measurement|SBP
Drug|Pharmacologic Substance|Hospital Course|4469,4478|false|false|false|C0012798|Diuretics|Diuretics
Event|Event|Hospital Course|4469,4478|false|false|false|||Diuretics
Event|Event|Hospital Course|4495,4499|false|false|false|||held
Finding|Mental Process|Hospital Course|4507,4514|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|4518,4530|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|4518,4530|false|false|false|||hyponatremia
Event|Event|Hospital Course|4540,4547|false|false|false|||treated
Event|Event|Hospital Course|4567,4576|false|false|false|||nutrition
Finding|Finding|Hospital Course|4567,4576|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|Hospital Course|4567,4576|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|Hospital Course|4567,4576|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|Hospital Course|4567,4576|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4567,4576|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Finding|Intellectual Product|Hospital Course|4578,4583|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Drug|Antibiotic|Hospital Course|4584,4595|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|4584,4595|false|false|false|||antibiotics
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4600,4607|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4600,4613|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|Hospital Course|4600,4613|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4608,4613|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|Hospital Course|4615,4624|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|4615,4624|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|4615,4624|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|Hospital Course|4636,4647|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|4636,4647|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|4654,4665|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Hospital Course|4654,4665|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Hospital Course|4654,4665|false|false|false|||therapeutic
Finding|Functional Concept|Hospital Course|4654,4665|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Hospital Course|4654,4665|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4654,4665|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|Hospital Course|4666,4678|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4666,4678|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|Hospital Course|4688,4696|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|4688,4696|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|4688,4696|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Cell|Hospital Course|4698,4708|false|false|false|C0023516|Leukocytes|white cell
Anatomy|Cell|Hospital Course|4704,4708|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|4704,4708|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|Hospital Course|4704,4714|false|false|false|C0007584|Cell Count|cell count
Event|Event|Hospital Course|4709,4714|false|false|false|||count
Drug|Biologically Active Substance|Hospital Course|4720,4735|false|false|false|C0005437|Bilirubin|total bilirubin
Drug|Organic Chemical|Hospital Course|4720,4735|false|false|false|C0005437|Bilirubin|total bilirubin
Finding|Physiologic Function|Hospital Course|4720,4735|false|false|false|C4553024|Total bilirubin metabolic function|total bilirubin
Lab|Laboratory or Test Result|Hospital Course|4720,4735|false|false|false|C0368753|Total bilirubin level|total bilirubin
Procedure|Laboratory Procedure|Hospital Course|4720,4735|false|false|false|C0201913|Bilirubin, total measurement|total bilirubin
Drug|Biologically Active Substance|Hospital Course|4726,4735|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Organic Chemical|Hospital Course|4726,4735|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Pharmacologic Substance|Hospital Course|4726,4735|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Event|Event|Hospital Course|4726,4735|false|false|false|||bilirubin
Procedure|Laboratory Procedure|Hospital Course|4726,4735|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|bilirubin
Event|Event|Hospital Course|4742,4751|false|false|false|||improving
Finding|Finding|Hospital Course|4755,4759|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4755,4759|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4755,4759|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|4763,4772|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4763,4772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4763,4772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4763,4772|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4763,4772|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|4783,4789|false|false|false|||follow
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4810,4815|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|4810,4815|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|4810,4815|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|4810,4815|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|4810,4815|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|4810,4815|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|4810,4815|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|4810,4815|false|false|false|C0872387|Procedures on liver|liver
Finding|Intellectual Product|Hospital Course|4836,4848|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|4836,4848|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|Hospital Course|4836,4857|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|Hospital Course|4836,4857|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|Hospital Course|4844,4848|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|4844,4848|false|false|false|||care
Finding|Finding|Hospital Course|4844,4848|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|4844,4848|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Hospital Course|4849,4857|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|4849,4857|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Disorder|Disease or Syndrome|Hospital Course|4887,4899|false|false|false|C0020625|Hyponatremia|HYPONATREMIA
Event|Event|Hospital Course|4887,4899|false|false|false|||HYPONATREMIA
Finding|Finding|Hospital Course|4901,4907|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|4901,4907|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Lab|Laboratory or Test Result|Hospital Course|4908,4919|false|true|false|C0752266|Hypovolemic|hypovolemic
Disorder|Disease or Syndrome|Hospital Course|4920,4932|false|true|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|4920,4932|false|false|false|||hyponatremia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4944,4953|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|4944,4953|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|4944,4953|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|4944,4953|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|4944,4953|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|4944,4953|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Disease or Syndrome|Hospital Course|4967,4979|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|4967,4979|false|false|false|||hyponatremia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4985,4990|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|4985,4990|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|4985,4990|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|4985,4990|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|4985,4990|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|4985,4990|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Hospital Course|4985,4990|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|4985,4990|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Hospital Course|4985,4998|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|Hospital Course|4991,4998|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|4991,4998|false|false|false|||disease
Event|Event|Hospital Course|5005,5018|false|false|false|||spironlactone
Event|Event|Hospital Course|5023,5027|false|false|false|||held
Event|Event|Hospital Course|5039,5048|false|false|false|||restarted
Event|Event|Hospital Course|5056,5066|false|false|false|||discretion
Finding|Functional Concept|Hospital Course|5056,5066|false|false|false|C5556474|Discretion|discretion
Finding|Classification|Hospital Course|5075,5085|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|5075,5085|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5086,5091|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|5086,5091|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|5086,5091|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|5086,5091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|5086,5091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|5086,5091|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|5086,5091|false|false|false|||liver
Finding|Finding|Hospital Course|5086,5091|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|5086,5091|false|false|false|C0872387|Procedures on liver|liver
Drug|Biologically Active Substance|Hospital Course|5112,5118|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|5112,5118|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|5112,5118|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|5112,5118|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|5112,5118|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|5112,5118|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Finding|Hospital Course|5122,5126|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|5122,5126|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|5122,5126|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|5131,5140|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5131,5140|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5131,5140|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5131,5140|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5131,5140|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|5163,5170|false|false|false|||advised
Event|Event|Hospital Course|5174,5182|false|false|false|||continue
Finding|Finding|Hospital Course|5185,5188|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|5185,5188|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|5185,5195|false|false|false|C0860871|Sodium decreased|low sodium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5185,5195|false|false|false|C0012169|Low sodium diet|low sodium
Drug|Biologically Active Substance|Hospital Course|5189,5195|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|5189,5195|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|5189,5195|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|5189,5195|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|5189,5195|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|5189,5195|false|false|false|C0337443|Sodium measurement|sodium
Drug|Food|Hospital Course|5197,5201|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|5197,5201|false|false|false|||diet
Finding|Functional Concept|Hospital Course|5197,5201|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5197,5201|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|5206,5210|false|false|false|||free
Finding|Functional Concept|Hospital Course|5206,5210|false|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|Hospital Course|5206,5216|false|false|false|C5572587|Free water|free water
Drug|Inorganic Chemical|Hospital Course|5211,5216|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Hospital Course|5211,5216|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Hospital Course|5211,5216|false|false|false|||water
Finding|Intellectual Product|Hospital Course|5211,5216|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5211,5216|false|false|false|C0020311|Hydrotherapy|water
Event|Event|Hospital Course|5217,5228|false|false|false|||restriction
Finding|Functional Concept|Hospital Course|5217,5228|false|false|false|C0443288|Restricted|restriction
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5254,5264|false|false|false|C0001973|Alcoholic Intoxication, Chronic|ALCOHOLISM
Event|Event|Hospital Course|5254,5264|false|false|false|||ALCOHOLISM
Finding|Body Substance|Hospital Course|5266,5273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|5266,5273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|5266,5273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|Hospital Course|5266,5277|false|false|false|C0332310|Has patient|Patient has
Event|Event|Hospital Course|5283,5289|false|false|false|||trying
Event|Event|Hospital Course|5293,5296|false|false|false|||cut
Event|Event|Hospital Course|5317,5324|false|false|false|||reports
Finding|Intellectual Product|Hospital Course|5317,5324|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|Hospital Course|5317,5324|false|false|false|C0700287|Reporting|reports
Drug|Organic Chemical|Hospital Course|5337,5344|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Hospital Course|5337,5344|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Hospital Course|5337,5344|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Individual Behavior|Hospital Course|5337,5351|false|false|false|C0001948|Alcohol consumption|alcohol intake
Event|Event|Hospital Course|5345,5351|false|false|false|||intake
Finding|Functional Concept|Hospital Course|5345,5351|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|5345,5351|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5389,5399|false|false|false|C2825032|Withdrawal (dysfunction)|withdrawal
Event|Activity|Hospital Course|5389,5399|false|false|false|C2349954|Withdraw (activity)|withdrawal
Event|Event|Hospital Course|5389,5399|false|false|false|||withdrawal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5389,5399|false|false|false|C3812880|Withdrawal - birth control|withdrawal
Finding|Sign or Symptom|Hospital Course|5389,5408|false|false|false|C0087169|Withdrawal Symptoms|withdrawal symptoms
Event|Event|Hospital Course|5400,5408|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|5400,5408|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5400,5408|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|5423,5431|true|false|false|||seizures
Finding|Sign or Symptom|Hospital Course|5423,5431|true|false|false|C0036572|Seizures|seizures
Event|Event|Hospital Course|5433,5439|false|false|false|||Shakes
Finding|Finding|Hospital Course|5433,5439|false|false|false|C0040822;C0392703|Shakes;Tremor|Shakes
Finding|Sign or Symptom|Hospital Course|5433,5439|false|false|false|C0040822;C0392703|Shakes;Tremor|Shakes
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5445,5459|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Hospital Course|5445,5459|false|false|false|||hallucinations
Event|Event|Hospital Course|5462,5469|false|false|false|||Reports
Finding|Intellectual Product|Hospital Course|5462,5469|false|false|false|C0684224|Report (document)|Reports
Procedure|Health Care Activity|Hospital Course|5462,5469|false|false|false|C0700287|Reporting|Reports
Event|Event|Hospital Course|5470,5478|false|false|false|||sobriety
Finding|Individual Behavior|Hospital Course|5470,5478|false|false|false|C0680686|sobriety|sobriety
Event|Event|Hospital Course|5491,5500|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5491,5500|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|5512,5520|false|false|false|||continue
Finding|Classification|Hospital Course|5521,5531|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|5521,5531|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|5532,5537|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5532,5537|false|false|false|C0034991|Rehabilitation therapy|rehab
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5544,5551|false|false|false|C0042027|Urinary tract|URINARY
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5544,5557|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|URINARY TRACT
Anatomy|Body System|Hospital Course|5544,5557|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|URINARY TRACT
Disorder|Disease or Syndrome|Hospital Course|5544,5567|false|false|false|C0042029|Urinary tract infection|URINARY TRACT INFECTION
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5552,5557|false|false|false|C1185740|Tract|TRACT
Disorder|Disease or Syndrome|Hospital Course|5558,5567|false|false|false|C0009450|Communicable Diseases|INFECTION
Event|Event|Hospital Course|5558,5567|false|false|false|||INFECTION
Finding|Pathologic Function|Hospital Course|5558,5567|false|false|false|C3714514|Infection|INFECTION
Event|Event|Hospital Course|5577,5584|false|false|false|||treated
Finding|Idea or Concept|Hospital Course|5598,5601|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5598,5601|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5603,5609|false|false|false|||course
Drug|Antibiotic|Hospital Course|5621,5632|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|5621,5632|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|5621,5632|false|false|false|||ceftriaxone
Event|Event|Hospital Course|5637,5644|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|5637,5644|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|5648,5651|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5648,5651|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|5648,5651|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|5648,5651|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|5648,5651|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Sign or Symptom|Hospital Course|5656,5665|false|false|false|C0004604|Back Pain|BACK PAIN
Attribute|Clinical Attribute|Hospital Course|5661,5665|false|false|false|C2598155||PAIN
Event|Event|Hospital Course|5661,5665|false|false|false|||PAIN
Finding|Functional Concept|Hospital Course|5661,5665|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Hospital Course|5661,5665|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Hospital Course|5666,5675|false|false|false|C0000726|Abdomen|ABDOMINAL
Finding|Sign or Symptom|Hospital Course|5666,5680|false|false|false|C0000737|Abdominal Pain|ABDOMINAL PAIN
Attribute|Clinical Attribute|Hospital Course|5676,5680|false|false|false|C2598155||PAIN
Event|Event|Hospital Course|5676,5680|false|false|false|||PAIN
Finding|Functional Concept|Hospital Course|5676,5680|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Hospital Course|5676,5680|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Event|Event|Hospital Course|5691,5698|false|false|false|||treated
Drug|Organic Chemical|Hospital Course|5714,5723|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|5714,5723|false|false|false|C0023660|lidocaine|lidocaine
Event|Event|Hospital Course|5714,5723|false|false|false|||lidocaine
Procedure|Laboratory Procedure|Hospital Course|5714,5723|false|false|false|C0202404|Lidocaine measurement|lidocaine
Event|Event|Hospital Course|5724,5731|false|false|false|||patches
Event|Event|Hospital Course|5735,5741|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|5746,5755|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|5746,5755|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|5746,5755|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|5746,5755|false|false|false|C0524222|Oxycodone measurement|oxycodone
Event|Event|Hospital Course|5759,5765|false|false|false|||needed
Event|Event|Hospital Course|5781,5789|false|false|false|||provided
Event|Event|Hospital Course|5803,5809|false|false|false|||course
Drug|Organic Chemical|Hospital Course|5813,5821|false|false|false|C0040610|tramadol|Tramadol
Drug|Pharmacologic Substance|Hospital Course|5813,5821|false|false|false|C0040610|tramadol|Tramadol
Event|Event|Hospital Course|5813,5821|false|false|false|||Tramadol
Procedure|Laboratory Procedure|Hospital Course|5813,5821|false|false|false|C1266765|Tramadol measurement (procedure)|Tramadol
Event|Event|Hospital Course|5825,5829|false|false|false|||take
Event|Event|Hospital Course|5833,5839|false|false|false|||needed
Finding|Functional Concept|Hospital Course|5847,5853|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|5847,5853|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|5847,5856|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|5847,5856|false|false|false|C1522577|follow-up|follow-up
Finding|Intellectual Product|Hospital Course|5866,5878|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|5866,5878|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|Hospital Course|5866,5887|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|Hospital Course|5866,5887|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|Hospital Course|5874,5878|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|5874,5878|false|false|false|||care
Finding|Finding|Hospital Course|5874,5878|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|5874,5878|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Hospital Course|5879,5887|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|5879,5887|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Event|Hospital Course|5893,5904|false|false|false|||understands
Finding|Idea or Concept|Hospital Course|5926,5935|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Finding|Intellectual Product|Hospital Course|5926,5935|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Drug|Pharmacologic Substance|Hospital Course|5936,5946|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|5936,5946|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|5936,5946|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|5960,5972|false|false|false|||discontinued
Finding|Intellectual Product|Hospital Course|5982,5987|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|5982,5997|false|false|false|C0267797|Acute hepatitis|acute hepatitis
Disorder|Disease or Syndrome|Hospital Course|5988,5997|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|Hospital Course|5988,5997|false|false|false|||hepatitis
Event|Event|Hospital Course|5998,6006|false|false|false|||resolves
Event|Event|Hospital Course|6011,6022|false|false|false|||Prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6011,6022|false|false|false|C0199176|Prophylactic treatment|Prophylaxis
Anatomy|Body Location or Region|Hospital Course|6027,6030|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|6027,6030|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|6027,6030|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|6031,6034|false|false|false|||ppx
Finding|Gene or Genome|Hospital Course|6031,6034|false|false|false|C1418850|PPP4C gene|ppx
Drug|Biologically Active Substance|Hospital Course|6043,6050|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|6043,6050|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|6043,6050|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|6043,6050|false|false|false|||heparin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6054,6059|true|false|false|C0021853|Intestines|Bowel
Procedure|Health Care Activity|Hospital Course|6054,6067|true|false|false|C5979615|Bowel Regimen|Bowel regimen
Event|Event|Hospital Course|6060,6067|true|false|false|||regimen
Finding|Intellectual Product|Hospital Course|6060,6067|true|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6060,6067|true|false|false|C0040808|Treatment Protocols|regimen
Drug|Organic Chemical|Hospital Course|6073,6082|true|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|Hospital Course|6073,6082|true|false|false|C0022957|lactulose|lactulose
Event|Event|Hospital Course|6073,6082|true|false|false|||lactulose
Drug|Pharmacologic Substance|Hospital Course|6087,6090|true|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|Hospital Course|6087,6090|true|false|false|||PPI
Finding|Physiologic Function|Hospital Course|6087,6090|true|false|false|C0871125|Prepulse Inhibition|PPI
Attribute|Clinical Attribute|Hospital Course|6094,6098|true|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|6094,6098|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|6094,6098|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6094,6109|true|false|false|C0002766|Pain management (procedure)|Pain management
Event|Event|Hospital Course|6099,6109|true|false|false|||management
Event|Occupational Activity|Hospital Course|6099,6109|true|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|6099,6109|true|false|false|C0376636|Disease Management|management
Drug|Organic Chemical|Hospital Course|6115,6124|true|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|6115,6124|true|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|6115,6124|true|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|6115,6124|true|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Hospital Course|6129,6138|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|6129,6138|false|false|false|C0023660|lidocaine|lidocaine
Event|Event|Hospital Course|6129,6138|false|false|false|||lidocaine
Procedure|Laboratory Procedure|Hospital Course|6129,6138|false|false|false|C0202404|Lidocaine measurement|lidocaine
Drug|Clinical Drug|Hospital Course|6129,6144|false|false|false|C1251704|Lidocaine Patch|lidocaine patch
Drug|Biomedical or Dental Material|Hospital Course|6139,6144|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|Hospital Course|6139,6144|false|false|false|||patch
Finding|Finding|Hospital Course|6139,6144|false|false|false|C0332461|Plaque (lesion)|patch
Event|Event|Hospital Course|6149,6162|false|false|false|||Communication
Finding|Social Behavior|Hospital Course|6149,6162|false|false|false|C0009452|Communication|Communication
Finding|Body Substance|Hospital Course|6164,6171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6164,6171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6164,6171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6176,6180|false|false|false|||Code
Event|Occupational Activity|Hospital Course|6176,6180|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|6176,6180|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Attribute|Clinical Attribute|Hospital Course|6198,6209|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6198,6209|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6198,6209|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6198,6209|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|6198,6222|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|6213,6222|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|6213,6222|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|6224,6236|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|6224,6236|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|6224,6236|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Event|Event|Hospital Course|6224,6236|false|false|false|||Multivitamin
Drug|Organic Chemical|Hospital Course|6238,6246|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Pharmacologic Substance|Hospital Course|6238,6246|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Drug|Vitamin|Hospital Course|6238,6246|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|thiamine
Event|Event|Hospital Course|6238,6246|false|false|false|||thiamine
Procedure|Laboratory Procedure|Hospital Course|6238,6246|false|false|false|C0373727|Thiamine measurement|thiamine
Drug|Organic Chemical|Hospital Course|6248,6254|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Hospital Course|6248,6254|false|false|false|C0178638|folate|folate
Drug|Vitamin|Hospital Course|6248,6254|false|false|false|C0178638|folate|folate
Event|Event|Hospital Course|6248,6254|false|false|false|||folate
Procedure|Laboratory Procedure|Hospital Course|6248,6254|false|false|false|C0523631|Folic acid measurement|folate
Drug|Organic Chemical|Hospital Course|6256,6270|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Hospital Course|6256,6270|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|Hospital Course|6256,6270|false|false|false|||spironolactone
Drug|Organic Chemical|Hospital Course|6284,6293|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|6284,6293|false|false|false|C0023660|lidocaine|lidocaine
Event|Event|Hospital Course|6284,6293|false|false|false|||lidocaine
Procedure|Laboratory Procedure|Hospital Course|6284,6293|false|false|false|C0202404|Lidocaine measurement|lidocaine
Drug|Clinical Drug|Hospital Course|6284,6299|false|false|false|C1251704|Lidocaine Patch|lidocaine patch
Drug|Biomedical or Dental Material|Hospital Course|6294,6299|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|Hospital Course|6294,6299|false|false|false|||patch
Finding|Finding|Hospital Course|6294,6299|false|false|false|C0332461|Plaque (lesion)|patch
Finding|Gene or Genome|Hospital Course|6300,6303|false|false|false|C1422467|CIAO3 gene|prn
Drug|Hazardous or Poisonous Substance|Hospital Course|6305,6313|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|Hospital Course|6305,6313|false|false|false|C0028040|nicotine|nicotine
Drug|Clinical Drug|Hospital Course|6305,6319|false|false|false|C0358855|Nicotine Transdermal Patch|nicotine patch
Drug|Biomedical or Dental Material|Hospital Course|6314,6319|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|Hospital Course|6314,6319|false|false|false|||patch
Finding|Finding|Hospital Course|6314,6319|false|false|false|C0332461|Plaque (lesion)|patch
Event|Event|Hospital Course|6323,6332|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6323,6332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6323,6332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6323,6332|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6323,6332|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6323,6344|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6333,6344|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6333,6344|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6333,6344|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6333,6344|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6349,6361|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|6349,6361|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|Hospital Course|6349,6361|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|Hospital Course|6349,6372|false|false|false|C0978787|Multivitamin tablet|Multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|6366,6372|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6366,6372|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|6386,6392|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6386,6392|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|6417,6425|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|Hospital Course|6417,6425|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|Hospital Course|6417,6425|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Event|Event|Hospital Course|6417,6425|false|false|false|||Thiamine
Procedure|Laboratory Procedure|Hospital Course|6417,6425|false|false|false|C0373727|Thiamine measurement|Thiamine
Drug|Organic Chemical|Hospital Course|6417,6429|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Pharmacologic Substance|Hospital Course|6417,6429|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Vitamin|Hospital Course|6417,6429|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Disorder|Neoplastic Process|Hospital Course|6426,6429|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|6426,6429|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|6426,6429|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|6426,6429|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|6426,6429|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|6437,6443|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6457,6463|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6457,6463|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|6488,6498|false|false|false|C0016410|folic acid|Folic Acid
Drug|Pharmacologic Substance|Hospital Course|6488,6498|false|false|false|C0016410|folic acid|Folic Acid
Drug|Vitamin|Hospital Course|6488,6498|false|false|false|C0016410|folic acid|Folic Acid
Procedure|Laboratory Procedure|Hospital Course|6488,6498|false|false|false|C0523631|Folic acid measurement|Folic Acid
Event|Event|Hospital Course|6494,6498|false|false|false|||Acid
Drug|Biomedical or Dental Material|Hospital Course|6504,6510|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6511,6514|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|6524,6530|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6524,6530|false|false|false|||Tablet
Drug|Hazardous or Poisonous Substance|Hospital Course|6555,6563|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|Hospital Course|6555,6563|false|false|false|C0028040|nicotine|Nicotine
Drug|Biomedical or Dental Material|Hospital Course|6576,6581|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|6576,6581|false|false|false|||Patch
Finding|Finding|Hospital Course|6576,6581|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Biomedical or Dental Material|Hospital Course|6601,6606|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|6601,6606|false|false|false|||Patch
Finding|Finding|Hospital Course|6601,6606|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Finding|Hospital Course|6614,6625|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Finding|Functional Concept|Hospital Course|6614,6625|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Drug|Organic Chemical|Hospital Course|6646,6655|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|6646,6655|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|Hospital Course|6646,6655|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|Hospital Course|6667,6672|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Hospital Course|6667,6672|false|false|false|C0332461|Plaque (lesion)|patch
Drug|Biomedical or Dental Material|Hospital Course|6683,6688|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|6683,6688|false|false|false|||Patch
Finding|Finding|Hospital Course|6683,6688|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Pharmacologic Substance|Hospital Course|6690,6699|false|false|false|C3812869|Medicated|Medicated
Event|Event|Hospital Course|6690,6699|false|false|false|||Medicated
Finding|Finding|Hospital Course|6690,6699|false|false|false|C3812868|Medicated (finding)|Medicated
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6700,6703|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6700,6703|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6700,6703|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6700,6703|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|6723,6728|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|6723,6728|false|false|false|||Patch
Finding|Finding|Hospital Course|6723,6728|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Pharmacologic Substance|Hospital Course|6730,6739|false|false|false|C3812869|Medicated|Medicated
Event|Event|Hospital Course|6730,6739|false|false|false|||Medicated
Finding|Finding|Hospital Course|6730,6739|false|false|false|C3812868|Medicated (finding)|Medicated
Drug|Biomedical or Dental Material|Hospital Course|6740,6747|false|false|false|C1710439|Topical Dosage Form|Topical
Finding|Functional Concept|Hospital Course|6740,6747|false|false|false|C1522168|Topical Route of Administration|Topical
Drug|Organic Chemical|Hospital Course|6768,6776|false|false|false|C0040610|tramadol|Tramadol
Drug|Pharmacologic Substance|Hospital Course|6768,6776|false|false|false|C0040610|tramadol|Tramadol
Event|Event|Hospital Course|6768,6776|false|false|false|||Tramadol
Procedure|Laboratory Procedure|Hospital Course|6768,6776|false|false|false|C1266765|Tramadol measurement (procedure)|Tramadol
Drug|Biomedical or Dental Material|Hospital Course|6783,6789|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6803,6809|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6839,6845|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|6850,6854|false|false|false|C2598155||pain
Event|Event|Hospital Course|6850,6854|false|false|false|||pain
Finding|Functional Concept|Hospital Course|6850,6854|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6850,6854|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|6865,6871|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|6876,6883|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|6891,6900|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6891,6900|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6891,6900|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6891,6900|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6891,6900|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6891,6912|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6891,6912|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6901,6912|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6901,6912|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6901,6912|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6914,6918|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6914,6918|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6914,6918|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6914,6918|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|6921,6930|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6921,6930|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6921,6930|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6921,6930|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6921,6930|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6921,6940|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6931,6940|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6931,6940|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6931,6940|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6931,6940|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6931,6940|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Hospital Course|6942,6959|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|Hospital Course|6950,6959|false|false|false|C0945731||diagnosis
Event|Event|Hospital Course|6950,6959|false|false|false|||diagnosis
Finding|Classification|Hospital Course|6950,6959|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|6950,6959|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6950,6959|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|Hospital Course|6961,6980|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|Hospital Course|6971,6980|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|Hospital Course|6971,6980|false|false|false|||hepatitis
Finding|Mental Process|Discharge Condition|7005,7011|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|7005,7018|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|7005,7018|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|7012,7018|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|7012,7018|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7020,7025|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|7020,7025|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|7030,7038|false|false|false|||coherent
Finding|Finding|Discharge Condition|7030,7038|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|7040,7045|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|7040,7062|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|7040,7062|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|7049,7062|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|7049,7062|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|7049,7062|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|7064,7069|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|7064,7069|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|7064,7069|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|7064,7069|false|false|false|||Alert
Finding|Finding|Discharge Condition|7064,7069|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|7064,7069|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|7064,7069|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|7074,7085|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|7074,7085|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|7087,7095|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|7087,7095|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|7087,7095|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|7096,7102|false|false|false|C5889824||Status
Event|Event|Discharge Condition|7096,7102|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|7096,7102|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|7104,7114|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|7104,7114|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|7104,7114|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|7104,7114|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|7104,7114|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|7117,7128|false|false|false|||Independent
Finding|Finding|Discharge Condition|7117,7128|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|7117,7128|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|7165,7173|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|7181,7189|false|false|false|C1547192|Organization unit type - Hospital|hospital
Disorder|Disease or Syndrome|Discharge Instructions|7194,7213|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|Discharge Instructions|7204,7213|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|Discharge Instructions|7204,7213|false|false|false|||hepatitis
Attribute|Clinical Attribute|Discharge Instructions|7226,7235|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|7226,7235|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|7226,7235|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|7226,7235|false|false|false|C1705253|Logical Condition|condition
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7250,7255|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|7250,7255|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|7250,7255|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|7250,7255|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|7250,7255|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|7250,7255|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Discharge Instructions|7250,7255|false|false|false|||liver
Finding|Finding|Discharge Instructions|7250,7255|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|7250,7255|false|false|false|C0872387|Procedures on liver|liver
Event|Event|Discharge Instructions|7256,7263|false|false|false|||becomes
Event|Event|Discharge Instructions|7264,7272|false|false|false|||inflamed
Drug|Organic Chemical|Discharge Instructions|7291,7298|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|7291,7298|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Discharge Instructions|7291,7298|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Individual Behavior|Discharge Instructions|7291,7305|false|false|false|C0001948|Alcohol consumption|alcohol intake
Event|Event|Discharge Instructions|7299,7305|false|false|false|||intake
Finding|Functional Concept|Discharge Instructions|7299,7305|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Discharge Instructions|7299,7305|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|Discharge Instructions|7321,7326|false|false|false|||noted
Event|Event|Discharge Instructions|7335,7337|false|false|false|||an
Anatomy|Cell|Discharge Instructions|7348,7358|false|false|false|C0023516|Leukocytes|white cell
Anatomy|Cell|Discharge Instructions|7354,7358|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Discharge Instructions|7354,7358|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|Discharge Instructions|7354,7364|false|false|false|C0007584|Cell Count|cell count
Event|Event|Discharge Instructions|7359,7364|false|false|false|||count
Event|Event|Discharge Instructions|7385,7393|false|false|false|||indicate
Disorder|Disease or Syndrome|Discharge Instructions|7395,7404|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|7395,7404|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|7395,7404|false|false|false|C3714514|Infection|infection
Event|Event|Discharge Instructions|7415,7422|false|false|false|||treated
Finding|Intellectual Product|Discharge Instructions|7430,7435|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|Discharge Instructions|7436,7442|false|false|false|||course
Drug|Antibiotic|Discharge Instructions|7446,7457|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|7446,7457|false|false|false|||antibiotics
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7465,7472|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7465,7478|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|Discharge Instructions|7465,7478|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|Discharge Instructions|7465,7488|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7473,7478|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|Discharge Instructions|7479,7488|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|7479,7488|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|7479,7488|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|Discharge Instructions|7505,7510|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7505,7510|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7505,7510|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Location or Region|Discharge Instructions|7516,7526|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|Discharge Instructions|7516,7526|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Finding|Body Substance|Discharge Instructions|7516,7532|false|false|false|C0003964|Peritoneal fluid (substance)|peritoneal fluid
Procedure|Laboratory Procedure|Discharge Instructions|7516,7532|false|false|false|C2053903|Peritoneal fluid analysis|peritoneal fluid
Drug|Substance|Discharge Instructions|7527,7532|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|7527,7532|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|7527,7532|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|7542,7548|false|false|false|||remain
Event|Event|Discharge Instructions|7549,7557|false|false|false|||negative
Finding|Classification|Discharge Instructions|7549,7557|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Discharge Instructions|7549,7557|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Discharge Instructions|7549,7557|false|false|false|C5237010|Expression Negative|negative
Event|Event|Discharge Instructions|7563,7567|false|false|false|||made
Event|Event|Discharge Instructions|7582,7589|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|7582,7589|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Discharge Instructions|7598,7609|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7598,7609|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|7598,7609|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|7598,7609|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|7615,7622|false|false|false|||stopped
Drug|Organic Chemical|Discharge Instructions|7628,7642|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|7628,7642|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|Discharge Instructions|7628,7642|false|false|false|||spironolactone
Disorder|Disease or Syndrome|Discharge Instructions|7656,7661|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7656,7661|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7656,7661|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|7656,7668|false|false|false|C0853174|Blood sodium|blood sodium
Drug|Biologically Active Substance|Discharge Instructions|7662,7668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Discharge Instructions|7662,7668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Discharge Instructions|7662,7668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Discharge Instructions|7662,7668|false|false|false|||sodium
Finding|Physiologic Function|Discharge Instructions|7662,7668|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Discharge Instructions|7662,7668|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|Discharge Instructions|7669,7675|false|false|false|||levels
Finding|Finding|Discharge Instructions|7682,7689|false|false|false|C4036057|Too low|too low
Event|Event|Discharge Instructions|7686,7689|false|false|false|||low
Finding|Finding|Discharge Instructions|7686,7689|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|7686,7689|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Discharge Instructions|7694,7699|false|false|false|||added
Drug|Organic Chemical|Discharge Instructions|7700,7708|false|false|false|C0040610|tramadol|Tramadol
Drug|Pharmacologic Substance|Discharge Instructions|7700,7708|false|false|false|C0040610|tramadol|Tramadol
Event|Event|Discharge Instructions|7700,7708|false|false|false|||Tramadol
Procedure|Laboratory Procedure|Discharge Instructions|7700,7708|false|false|false|C1266765|Tramadol measurement (procedure)|Tramadol
Event|Event|Discharge Instructions|7712,7716|false|false|false|||take
Event|Event|Discharge Instructions|7720,7726|false|false|false|||needed
Finding|Sign or Symptom|Discharge Instructions|7731,7740|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Discharge Instructions|7736,7740|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7736,7740|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7736,7740|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7736,7740|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Health Care Activity|Discharge Instructions|7745,7753|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7754,7766|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|7754,7766|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|7754,7766|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

