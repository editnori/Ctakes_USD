CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Personal History of Coronary Artery Disease|Attribute|false|false||history of coronary artery diseasenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Ischemic|Finding|false|false||ischemicnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|MDFAttributeType - Fraction|Finding|false|false||fractionnull|Fraction of|LabModifier|false|false||fractionnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Peripheral Vascular Diseases|Disorder|false|false||peripheral vascular diseasenull|Peripheral|Modifier|false|false||peripheralnull|Vascular Diseases|Disorder|false|false||vascular diseasenull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Chronic disease|Disorder|false|false||disease, chronicnull|Disease|Disorder|false|false||diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false||kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Disease|Disorder|false|false||diseasenull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|null|Time|false|false||priornull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Hypertensive disease|Disorder|false|false||HTNnull|Dyslipidemias|Disorder|false|false||dyslipidemianull|Several days|Finding|false|false||several daysnull|Several|LabModifier|false|false||severalnull|day|Time|false|false||daysnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Patients|Subject|false|false||Patientsnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||acute onsetnull|Sudden onset (attribute)|Time|false|false||acute onset
null|acute|Time|false|false||acute onsetnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Prior functioning.stairs|Finding|false|false||stairsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Does sit|Finding|false|false||sit
null|Sitting position|Finding|false|false||sit
null|HHAT gene|Finding|false|false||sit
null|SIT1 gene|Finding|false|false||sitnull|Breath|Finding|false|false||breathnull|day|Time|false|false||daysnull|null|Time|false|false||priornull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Prior functioning.stairs|Finding|false|false||stairsnull|Has difficulty doing (qualifier value)|Finding|true|false||difficultynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Associated with|Modifier|false|false||associatednull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Palpitations|Finding|true|false||palpitationsnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Lightheadedness|Finding|false|false||lightheadednessnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Further|Modifier|false|false||furthernull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Fever|Finding|false|false||feversnull|Chills|Finding|false|false||chillsnull|Chest discomfort|Finding|false|false||chest discomfortnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Discomfort|Finding|false|false||discomfortnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|True or Present Nearly Every Day|Finding|false|false||nearly every daynull|Nearly every day|Time|false|false||nearly every daynull|Nearly|Modifier|false|false||nearlynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Gain|LabModifier|false|false||gainnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|More|LabModifier|false|false||morenull|Current (present time)|Time|false|false||currentlynull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Missing|Modifier|false|false||missednull|Dosage|LabModifier|false|false||dosesnull|Abdominal bloating|Finding|false|false||abdominal bloating
null|Abdomen distended|Finding|false|false||abdominal bloatingnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Abdominal bloating|Finding|false|false||bloating
null|Abdomen distended|Finding|false|false||bloatingnull|Constipation|Finding|false|false||constipationnull|Recent|Time|false|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|husband|Subject|false|false||husbandnull|Viral|Finding|false|false||viralnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Obvious|Modifier|false|false||Obviousnull|Bilateral|Modifier|false|false||bilateralnull|Wheezing|Finding|false|false||wheezingnull|Hypervolemia (finding)|Finding|true|false||volume overloadnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|Fracture of second cervical vertebra|Disorder|false|false||axisnull|Axis vertebra|Anatomy|false|false||axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|Interval|Time|false|false||intervalsnull|Corrected QT Interval|LabModifier|false|false||QTcnull|null|Phenomenon|false|false||wavesnull|aVF|Modifier|false|false||aVFnull|aVF|Modifier|false|false||aVFnull|Lateral|Modifier|false|false||lateralnull|Sexually Transmitted Diseases|Disorder|false|false||STDsnull|Laboratory test finding|Lab|false|false||Labsnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|Bone Morphogenetic Proteins|Drug|false|false||BMP
null|Bone Morphogenetic Proteins|Drug|false|false||BMPnull|carmustine/methotrexate/procarbazine protocol|Procedure|false|false||BMPnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Urobilinogen|Drug|false|false||urobilinogen
null|Urobilinogen|Drug|false|false||urobilinogennull|Urobilinogen measurement|Procedure|false|false||urobilinogennull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|bilirubin preparation|Drug|false|false||bilirubin
null|bilirubin preparation|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubinnull|Bilirubin, total measurement|Procedure|false|false||bilirubin
null|blood bilirubin level test|Procedure|false|false||bilirubinnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||nitrite
null|Nitrites|Drug|false|false||nitrite
null|Nitrites|Drug|false|false||nitrite
null|Nitrites|Drug|false|false||nitrite
null|nitrite ion|Drug|false|false||nitrite
null|nitrite ion|Drug|false|false||nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||protein
null|Proteins|Drug|false|false||proteinnull|Protein Info|Finding|false|false||proteinnull|Protein measurement|Procedure|false|false||proteinnull|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucose
null|glucose|Drug|false|false||glucosenull|Glucose measurement|Procedure|false|false||glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||ketonesnull|Toxic effect of ketones|Disorder|false|false||ketonesnull|Ketone bodies measurement, quantitative|Procedure|false|false||ketones
null|Urine ketone test|Procedure|false|false||ketonesnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Leukocytes|Anatomy|false|false||WBCnull|bacteria aspects|Finding|false|false||bacterianull|Bacteria <walking sticks>|Entity|false|false||bacteria
null|Bacteria|Entity|false|false||bacterianull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Plain chest X-ray|Procedure|false|false||CXRnull|Lung|Anatomy|false|false||Lungsnull|Moderate Response|Finding|false|false||moderately
null|Moderate|Finding|false|false||moderately
null|Moderate Effect|Finding|false|false||moderatelynull|Moderate (severity modifier)|Modifier|false|false||moderately
null|Moderation|Modifier|false|false||moderatelynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Asymmetry (qualifier value)|Modifier|false|false||asymmetricnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Lung opacity|Finding|false|false||lung opacitynull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Enlargement procedure|Procedure|false|false||enlargednull|Enlarged|Modifier|false|false||enlargednull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary vascular congestion|Disorder|false|false||pulmonary vascular congestionnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Congestion|Finding|false|false||congestionnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Pneumothorax|Disorder|false|false||pneumothoraxnull|Structure of right lower lobe of lung|Anatomy|false|false||Right lower lobenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Pneumonia|Disorder|false|false||pneumonianull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Clinical setting|Modifier|false|false||clinical settingnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Atelectasis|Finding|false|false||atelectasisnull|Asymmetry (qualifier value)|Modifier|false|false||asymmetricnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Experimental Finding|Finding|false|false||finding
null|Signs and Symptoms|Finding|false|false||finding
null|Finding|Finding|false|false||findingnull|Lateral|Modifier|false|false||lateralnull|View|Modifier|false|false||viewsnull|Helpful|Modifier|false|false||helpfulnull|Further|Modifier|false|false||furthernull|Knowledge acquisition using a method of assessment|Finding|false|false||assessmentnull|assessment of cognitive functions|Procedure|false|false||assessment
null|Physical Examination|Procedure|false|false||assessment
null|Nutrition Assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Personal care assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Evaluation procedure|Procedure|false|false||assessment
null|Evaluation|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessmentnull|Assessed|Event|false|false||assessmentnull|Consultation|Procedure|false|false||Consultsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycinnull|ceftriaxone|Drug|false|false||CefTRIAXone
null|ceftriaxone|Drug|false|false||CefTRIAXonenull|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONEnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|ceftriaxone|Drug|false|false||CefTRIAXone
null|ceftriaxone|Drug|false|false||CefTRIAXonenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycin
null|azithromycin|Drug|false|false||Azithromycinnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Transfer - product ownership|Finding|false|false||Transfer
null|Transfer Technique|Finding|false|false||Transfer
null|ActClass - transfer|Finding|false|false||Transfer
null|null|Finding|false|false||Transfernull|Transfer (immobility management)|Procedure|false|false||Transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Aftercare|Procedure|false|false||after treatmentnull|Post-Therapy|Time|false|false||after treatmentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Continuous|Finding|false|false||ongoingnull|Dyspnea|Finding|false|false||SOBnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Reactive Oxygen Species|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|Reactive Oxygen Species|Drug|false|false||ROSnull|ROS1 wt Allele|Finding|false|false||ROS
null|ROS1 gene|Finding|false|false||ROSnull|Review of systems (procedure)|Procedure|false|false||ROSnull|rostral sulcus|Anatomy|false|false||ROSnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Peripheral Vascular Diseases|Disorder|false|false||Peripheral vascular diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false||vascular diseasenull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Disease|Disorder|false|false||diseasenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type II Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type II Diabetesnull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Diabetic Retinopathy|Disorder|false|false||diabetic retinopathynull|Diabetic|Finding|false|false||diabeticnull|Retinal Diseases|Disorder|false|false||retinopathynull|Obesity|Disorder|false|false||Obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|false|false||Obesitynull|Terminal esophageal web|Disorder|false|false||Esophageal ringnull|Esophageal Diseases|Disorder|false|false||Esophagealnull|Esophageal|Modifier|false|false||Esophagealnull|Ring Dosage Form|Drug|false|false||ringnull|Ring device|Device|false|false||ringnull|Annular shape|Modifier|false|false||ringnull|Ring Dosing Unit|LabModifier|false|false||ringnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Bilateral|Modifier|false|false||Bilateralnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false||tibialnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||Stage IVnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Hypertensive disease|Disorder|false|false||HTNnull|Hyperparathyroidism, Secondary|Disorder|false|false||secondary hyperparathyroidismnull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Hyperparathyroidism|Disorder|false|false||hyperparathyroidismnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Gout|Disorder|false|false||Goutnull|Niece|Subject|false|false||Niecenull|Sorting - Cell Movement|Finding|false|false||sort
null|Sorting (Cognition)|Finding|false|false||sortnull|Sorting|Event|false|false||sortnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Lung diseases|Disorder|false|false||lung diseasenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Disease|Disorder|false|false||diseasenull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Early|Time|false|false||earlynull|DFFB protein, human|Drug|true|false||CAD
null|DFFB protein, human|Drug|true|false||CADnull|Cold Hemagglutinin Disease|Disorder|true|false||CAD
null|Coronary heart disease|Disorder|true|false||CAD
null|Coronary Artery Disease|Disorder|true|false||CADnull|CAD gene|Finding|true|false||CAD
null|CALD1 wt Allele|Finding|true|false||CAD
null|B4GALNT2 gene|Finding|true|false||CAD
null|DFFB wt Allele|Finding|true|false||CAD
null|ACOD1 gene|Finding|true|false||CAD
null|DFFB gene|Finding|true|false||CADnull|cytarabine/daunorubicin protocol|Procedure|true|false||CAD
null|Computer Assisted Diagnosis|Procedure|true|false||CAD
null|Collision-Induced Dissociation|Procedure|true|false||CAD
null|CyADIC regimen|Procedure|true|false||CADnull|Caddo language|Entity|true|false||CADnull|Sudden Cardiac Death|Finding|true|false||sudden cardiac deathnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Cardiac Death|Finding|true|false||cardiac deathnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Event Consequence - Death|Finding|false|false||death
null|Death (finding)|Finding|false|false||death
null|Cessation of life|Finding|false|false||deathnull|Known|Modifier|false|false||knownnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Pleasant|Finding|false|false||Pleasantnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Breath|Finding|false|false||breathsnull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Jugular venous engorgement|Finding|false|false||JVDnull|Malignant neoplasm of heart|Disorder|false|false||HEART
null|benign neoplasm of heart|Disorder|false|false||HEARTnull|HEART PROBLEM|Finding|false|false||HEARTnull|Chest>Heart|Anatomy|false|false||HEART
null|Heart|Anatomy|false|false||HEARTnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||LUNGSnull|cetrimonium bromide|Drug|false|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Obese abdomen|Finding|false|false||Obese abdomennull|Obesity|Disorder|false|false||Obesenull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Protective muscle spasm|Finding|false|false||guardingnull|Hepatosplenomegaly|Finding|false|false||hepatosplenomegalynull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Cyanosis|Finding|true|false||cyanosisnull|Clubbing|Disorder|true|false||clubbingnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|PURPOSE (pharmacologic preparation)|Drug|false|false||purpose
null|PURPOSE (pharmacologic preparation)|Drug|false|false||purposenull|Purpose|Finding|false|false||purposenull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Excoriation|Disorder|true|false||excoriationsnull|Lesion|Finding|true|false||lesionsnull|Skin rash|Finding|false|false||rashes
null|Exanthema|Finding|false|false||rashesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Jugular venous engorgement|Finding|true|false||JVDnull|Carotid bruit|Finding|true|false||carotid bruitsnull|Carotid Arteries|Anatomy|false|false||carotidnull|Bruit|Finding|true|false||bruitsnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|cetrimonium bromide|Drug|false|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Symmetric Relationship|Finding|false|false||Symmetric
null|Symmetrical|Finding|false|false||Symmetricnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Pitting edema|Finding|true|false||pitting edemanull|Pitting|Finding|true|false||pittingnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB-6|Drug|false|false||MB-6null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 5|Drug|false|false||MB-5null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false||Base
null|Base|Drug|false|false||Base
null|Dental Base|Drug|false|false||Base
null|base - RoleClass|Drug|false|false||Basenull|Base - General Qualifier|Finding|false|false||Base
null|BPIFA4P gene|Finding|false|false||Base
null|Base - RX Component Type|Finding|false|false||Basenull|Anatomical base|Anatomy|false|false||Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|null|Finding|false|false||left atrial volumenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false||atrialnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Html Link Type - index|Finding|false|false||index
null|Index|Finding|false|false||index
null|Indexes|Finding|false|false||indexnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Right atrial pressure|Attribute|false|false||right atrial pressure
null|null|Attribute|false|false||right atrial pressurenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Atrial Pressure|Finding|false|false||atrial pressurenull|Heart Atrium|Anatomy|false|false||atrialnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mmHgnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Wall of ventricle|Anatomy|false|false||ventricular wallnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||left ventricular systolic dysfunctionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Basal|Modifier|false|false||basalnull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Inferolateral|Modifier|false|false||inferolateralnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Middle|Modifier|false|false||midnull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Doppler studies|Procedure|false|false||Dopplernull|Observation parameter|Finding|false|false||parametersnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Grade|Finding|false|false||with Gradenull|Clavien-Dindo Grade II|Finding|false|false||Grade II
null|G2 stage (tumor staging)|Finding|false|false||Grade II
null|Disease Grade 2|Finding|false|false||Grade II
null|Grade two rank|Finding|false|false||Grade IInull|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Diastolic dysfunction|Finding|false|false||diastolic dysfunctionnull|Diastole|Attribute|false|false||diastolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Diameter (qualifier value)|LabModifier|false|false||diametersnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Sequencing - Ascending|Finding|false|false||ascending
null|Ascend (action)|Finding|false|false||ascendingnull|Ascending|Modifier|false|false||ascendingnull|Age-Related Clonal Hematopoiesis|Finding|false|false||arch
null|ZBTB8OS gene|Finding|false|false||archnull|Arch of foot|Anatomy|false|false||arch
null|Structure of nucleus infundibularis hypothalami|Anatomy|false|false||arch
null|ARCH|Anatomy|false|false||archnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Aortic Valve Stenosis|Finding|false|false||aortic stenosisnull|Aorta|Anatomy|false|false||aorticnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|AORTIC VALVE DISEASE 3|Disorder|true|false||aortic valve stenosis
null|Stenosis of aorta|Disorder|true|false||aortic valve stenosisnull|Aortic Valve Stenosis|Finding|true|false||aortic valve stenosisnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|true|false||stenosisnull|Stenosis <Pimeliinae>|Entity|true|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Sequence Chromatogram|Finding|false|false||Tracenull|Trace Dosing Unit|LabModifier|false|false||Trace
null|trace amount|LabModifier|false|false||Trace
null|unknown - trace|LabModifier|false|false||Tracenull|Aorta|Anatomy|false|false||aorticnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Moderate Response|Finding|false|false||moderately
null|Moderate|Finding|false|false||moderately
null|Moderate Effect|Finding|false|false||moderatelynull|Moderate (severity modifier)|Modifier|false|false||moderately
null|Moderation|Modifier|false|false||moderatelynull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Tricuspid|Modifier|false|false||tricuspidnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Pericardial effusion|Disorder|true|false||pericardial effusionnull|Pericardial effusion body substance|Finding|true|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|true|false||effusion
null|null|Finding|true|false||effusion
null|effusion|Finding|true|false||effusionnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||LV systolic dysfunctionnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Old myocardial infarction|Finding|false|false||prior myocardial infarctionnull|null|Time|false|false||priornull|Myocardial Infarction|Disorder|false|false||myocardial infarctionnull|null|Attribute|false|false||myocardial infarctionnull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false||infarctionnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Clavien-Dindo Grade II|Finding|false|false||Grade II
null|G2 stage (tumor staging)|Finding|false|false||Grade II
null|Disease Grade 2|Finding|false|false||Grade II
null|Grade two rank|Finding|false|false||Grade IInull|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Left ventricular diastolic dysfunction|Disorder|false|false||LV diastolic dysfunctionnull|Diastolic dysfunction|Finding|false|false||diastolic dysfunctionnull|Diastole|Attribute|false|false||diastolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|null|Time|false|false||priornull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|regional|Modifier|false|false||Regional
null|Local|Modifier|false|false||Regionalnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Greater|LabModifier|false|false||greaternull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Plain chest X-ray|Procedure|false|false||CXRnull|LAT protein, human|Drug|false|false||LAT
null|L-Type Amino Acid Transporter|Drug|false|false||LAT
null|L-Type Amino Acid Transporter|Drug|false|false||LAT
null|ORC3 protein, human|Drug|false|false||LAT
null|ORC3 protein, human|Drug|false|false||LAT
null|LAT protein, human|Drug|false|false||LATnull|LAT gene|Finding|false|false||LAT
null|ORC3 wt Allele|Finding|false|false||LAT
null|ORC3 gene|Finding|false|false||LAT
null|SPNS1 gene|Finding|false|false||LATnull|Latin Language|Entity|false|false||LATnull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|true|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Bilateral|Modifier|false|false||BILATERALnull|Lower Extremity|Anatomy|false|false||LOWER EXTREMITYnull|Body Site Modifier - Lower|Anatomy|false|false||LOWERnull|Lower (action)|Event|false|false||LOWERnull|Lower - spatial qualifier|Modifier|false|false||LOWERnull|Limb structure|Anatomy|false|false||EXTREMITYnull|Doppler Ultrasound (procedure)|Procedure|false|false||DOPPLER ULTRASOUNDnull|Doppler studies|Procedure|false|false||DOPPLERnull|Ultrasonic|Finding|false|false||ULTRASOUNDnull|Urological ultrasound|Procedure|false|false||ULTRASOUND
null|Ultrasonography|Procedure|false|false||ULTRASOUNDnull|ultrasound device|Device|false|false||ULTRASOUNDnull|Ultrasonic Shockwave|Phenomenon|false|false||ULTRASOUND
null|Ultrasonics (sound)|Phenomenon|false|false||ULTRASOUNDnull|Thrombosis|Finding|false|false||thrombosisnull|Pair|Modifier|false|false||pairednull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false||tibialnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Deep Vein Thrombosis|Disorder|true|false||deep venous thrombosisnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous thrombosis after immobility|Finding|true|false||venous thrombosis
null|Venous Thrombosis|Finding|true|false||venous thrombosisnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|true|false||thrombosisnull|Limb structure|Anatomy|false|false||extremitynull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|Maximal (qualifier value)|Modifier|false|false||maximalnull|Maximum|LabModifier|false|false||maximalnull|Diameter (qualifier value)|LabModifier|false|false||diameternull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Enterococcus|Entity|false|false||ENTEROCOCCUS SPnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|cfu/mL|LabModifier|false|false||CFU/mLnull|Colony-forming unit|LabModifier|false|false||CFUnull|per milliliter|LabModifier|false|false||/mLnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Pending - Allergy Clinical Status|Finding|false|false||PENDING
null|Pending - referral status|Finding|false|false||PENDINGnull|Pending - status|Time|false|false||PENDINGnull|pending - ManagedParticipationStatus|Modifier|false|false||PENDING
null|pending - RoleStatus|Modifier|false|false||PENDING
null|Pending - Day type|Modifier|false|false||PENDINGnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Pending - Allergy Clinical Status|Finding|false|false||PENDING
null|Pending - referral status|Finding|false|false||PENDINGnull|Pending - status|Time|false|false||PENDINGnull|pending - ManagedParticipationStatus|Modifier|false|false||PENDING
null|pending - RoleStatus|Modifier|false|false||PENDING
null|Pending - Day type|Modifier|false|false||PENDINGnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Ischemic|Finding|false|false||ischemicnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||LV systolic dysfunctionnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Pad Dosage Form|Drug|false|false||PADnull|Pad Mass|Disorder|false|false||PAD
null|Peripheral Arterial Diseases|Disorder|false|false||PADnull|PADI4 wt Allele|Finding|false|false||PAD
null|PADI4 gene|Finding|false|false||PAD
null|DHX40 gene|Finding|false|false||PADnull|PAD Regimen|Procedure|false|false||PADnull|Strucure of thick cushion of skin|Anatomy|false|false||PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|null|Time|false|false||priornull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Subacute|Time|false|false||subacutenull|Dyspnea|Finding|false|false||SOBnull|Weight Gain|Finding|false|false||weight gain
null|Gaining Weight question|Finding|false|false||weight gainnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Gain|LabModifier|false|false||gainnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exacerbation|Finding|false|false||exacerbationnull|Diuresis|Finding|false|false||diuresisnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Rapid|Modifier|false|false||rapidnull|Improvement|Finding|false|false||improvementnull|subjective (symptom)|Finding|false|false||subjectivenull|null|Attribute|false|false||subjectivenull|Subjective observation (qualifier value)|Modifier|false|false||subjectivenull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Acute deep venous thrombosis|Disorder|false|false||acute DVTnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Plain chest X-ray|Procedure|false|false||CXRnull|Language Ability - Sign|Finding|true|false||sign
null|Physical findings|Finding|true|false||signnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Improvement|Finding|false|false||improvementnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Supplement|Finding|true|false||supplementalnull|Requirement|Finding|false|false||requirementnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|exacerbation acute|Finding|false|false||acute exacerbationnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Exacerbation|Finding|false|false||exacerbationnull|Chronic diastolic heart failure|Disorder|false|false||chronic diastolic heart failurenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Heart Failure, Diastolic|Disorder|false|false||diastolic heart failurenull|Diastole|Attribute|false|false||diastolicnull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Dry body weight (observable entity)|Subject|false|false||Dry weightnull|dry weight (physical finding)|LabModifier|false|false||Dry weightnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Precipitating Factors|Attribute|false|false||triggernull|Triggered by|Modifier|false|false||triggernull|Allergy Clinical Status - Suspect|Finding|false|false||suspect
null|Suspected (qualifier value)|Finding|false|false||suspectnull|Diet|Drug|false|false||dietarynull|Uncontrolled|Modifier|false|false||uncontrollednull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|ACSS2 protein, human|Drug|true|false||ACS
null|ACSS2 protein, human|Drug|true|false||ACSnull|Acrocallosal Syndrome|Disorder|true|false||ACS
null|Acute Chest Syndrome|Disorder|true|false||ACSnull|ACS - Activity Card Sort|Finding|true|false||ACS
null|American Community Survey|Finding|true|false||ACS
null|ACCS gene|Finding|true|false||ACS
null|CO-methylating acetyl-CoA synthase activity|Finding|true|false||ACS
null|PLA2G15 gene|Finding|true|false||ACS
null|ACSS2 wt Allele|Finding|true|false||ACS
null|ACSS2 gene|Finding|true|false||ACS
null|acetate-CoA ligase activity|Finding|true|false||ACSnull|anterior calcarine sulcus (human only)|Anatomy|false|false||ACSnull|Alternate Care Site|Device|true|false||ACSnull|American College of Surgeons|Entity|true|false||ACS
null|American Cancer Society|Entity|true|false||ACS
null|Alternate Care Site|Entity|true|false||ACSnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Transthoracic echocardiography|Procedure|true|false||TTEnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||LV systolic dysfunctionnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|null|Time|false|false||priornull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false||infarctionnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Clavien-Dindo Grade II|Finding|false|false||Grade II
null|G2 stage (tumor staging)|Finding|false|false||Grade II
null|Disease Grade 2|Finding|false|false||Grade II
null|Grade two rank|Finding|false|false||Grade IInull|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Diastolic dysfunction|Finding|false|false||diastolic dysfunctionnull|Diastole|Attribute|false|false||diastolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Similarity|Modifier|false|false||similarnull|null|Time|false|false||priornull|Transthoracic echocardiography|Procedure|false|false||TTEnull|doubt|Finding|false|false||Doubtnull|Peptide Nucleic Acids|Drug|false|false||PNAnull|Plain chest X-ray|Procedure|false|false||CXRnull|Lacking|Modifier|false|false||lacknull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|doubt|Finding|false|false||doubtnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Wells syndrome|Disorder|false|false||Wellsnull|Water Wells|Device|false|false||Wellsnull|Score|Finding|false|false||scorenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Diuresis|Finding|false|false||diuresisnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Rapid|Modifier|false|false||rapidnull|Improvement|Finding|false|false||improvementnull|subjective (symptom)|Finding|false|false||subjectivenull|null|Attribute|false|false||subjectivenull|Subjective observation (qualifier value)|Modifier|false|false||subjectivenull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Early|Time|false|false||earliernull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Observation parameter|Finding|false|false||parametersnull|Clinical Trials|Procedure|false|false||trialnull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Hyperkalemia|Finding|false|false||hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||hyperkalemianull|Increased frequency of micturition|Finding|false|false||Urinary frequencynull|Urinary tract|Anatomy|false|false||Urinarynull|urinary|Modifier|false|false||Urinarynull|Frequency|Finding|false|false||frequency
null|How Often|Finding|false|false||frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Urge Incontinence|Finding|false|false||urge incontinencenull|Incontinence|Disorder|false|false||incontinencenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Diuresis|Finding|false|false||diuresisnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Colonization|Finding|false|false||colonizationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Patient Condition Code - Stable|Finding|false|false||STABLEnull|Stable status|Modifier|false|false||STABLEnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Recent|Time|false|false||recentnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|true|false||bleedingnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Multifactorial|Finding|false|false||multifactorialnull|Anemia of chronic disease|Disorder|false|false||anemia of chronic diseasenull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Chronic disease|Disorder|false|false||chronic diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Disease|Disorder|false|false||diseasenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Production Processing ID|Finding|false|false||productionnull|production|Event|false|false||productionnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|blood anion gap (lab test)|Procedure|false|false||anion gap
null|Anion gap measurement|Procedure|false|false||anion gapnull|Anion Gap|Attribute|false|false||anion gapnull|Anion gap result|Lab|false|false||anion gapnull|Anions|Drug|false|false||anionnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||gap
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||gap
null|GTPase-Activating Proteins|Drug|false|false||gap
null|GTPase-Activating Proteins|Drug|false|false||gapnull|RASA1 wt Allele|Finding|false|false||gap
null|RASA1 gene|Finding|false|false||gapnull|Gap (space)|Modifier|false|false||gapnull|Metabolic acidosis|Finding|false|false||metabolic acidosisnull|Metabolic Process, Cellular|Finding|false|false||metabolic
null|Metabolic|Finding|false|false||metabolicnull|Multisection metabolic|Procedure|false|false||metabolicnull|Acidosis|Finding|false|false||acidosisnull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Recent|Time|false|false||recentnull|rectal discharge diarrhea (physical finding)|Finding|true|false||diarrhea
null|Diarrhea|Finding|true|false||diarrheanull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Renal tubular acidosis|Disorder|false|false||RTAnull|HHV8 ORF50 Gene|Finding|false|false||RTA
null|MRGPRF gene|Finding|false|false||RTA
null|RBFOX2 gene|Finding|false|false||RTAnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Stage level 4|Finding|false|false||Stage IVnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Chronic Kidney Diseases|Disorder|false|false||Chronic Kidney Diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false||Kidney Diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||Kidney
null|Benign neoplasm of kidney|Disorder|false|false||Kidneynull|Kidney problem|Finding|false|false||Kidneynull|examination of kidney|Procedure|false|false||Kidney
null|Procedures on Kidney|Procedure|false|false||Kidneynull|Kidney|Anatomy|false|false||Kidney
null|Both kidneys|Anatomy|false|false||Kidneynull|Disease|Disorder|false|false||Diseasenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Hypertensive disease|Disorder|false|false||HTNnull|Current (present time)|Time|false|false||currentlynull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Phos <Photinae>|Entity|false|false||Phosnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Calcitriol Drug Class|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|Calcitriol Drug Class|Drug|false|false||calcitriolnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||LV systolic dysfunctionnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Old myocardial infarction|Finding|false|false||prior myocardial infarctionnull|null|Time|false|false||priornull|Myocardial Infarction|Disorder|false|false||myocardial infarctionnull|null|Attribute|false|false||myocardial infarctionnull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false||infarctionnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Similarity|Modifier|false|false||similarnull|null|Time|false|false||priornull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Observation parameter|Finding|false|false||parametersnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Once a day, at bedtime|Time|false|false||qHSnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type II Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type II Diabetesnull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Last|Modifier|false|false||lastnull|Glycosylated hemoglobin A|Drug|false|false||HbA1C
null|Glycosylated hemoglobin A|Drug|false|false||HbA1Cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1Cnull|Excellent - LanguageAbilityProficiency|Modifier|false|false||excellent
null|Excellent - Specimen Quality|Modifier|false|false||excellent
null|Excellent (qualifier value)|Modifier|false|false||excellentnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Recent|Time|false|false||recentlynull|Prediabetes syndrome|Disorder|false|false||pre-diabeticnull|Concept model range (foundation metadata concept)|Finding|false|false||rangenull|Sample Range|LabModifier|false|false||range
null|Range|LabModifier|false|false||rangenull|Continuous|Finding|false|false||Continuenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|Blood Glucose|Drug|false|false||blood sugarnull|Blood glucose measurement|Procedure|false|false||blood sugarnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|raw sugar|Drug|false|false||sugar
null|raw sugar|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Carbohydrates|Drug|false|false||sugarnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Blood Glucose|Drug|false|false||blood sugarnull|Blood glucose measurement|Procedure|false|false||blood sugarnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|raw sugar|Drug|false|false||sugar
null|raw sugar|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Carbohydrates|Drug|false|false||sugarnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Insomnia homeopathic medication|Drug|false|false||Insomnianull|Sleeplessness|Finding|false|false||Insomnianull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|Gout|Disorder|false|false||Goutnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|allopurinol|Drug|false|false||allopurinol
null|allopurinol|Drug|false|false||allopurinolnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Diuretic [APC]|Drug|false|false||diuretic
null|Diuretics|Drug|false|false||diureticnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Daily|Time|false|false||dailynull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|EPO protein, human|Drug|false|false||epo
null|epoetin alfa|Drug|false|false||epo
null|epoetin alfa|Drug|false|false||epo
null|Erythropoietin|Drug|false|false||epo
null|Erythropoietin|Drug|false|false||epo
null|Erythropoietin|Drug|false|false||epo
null|EPO protein, human|Drug|false|false||eponull|EPO gene|Finding|false|false||epo
null|TIMP1 wt Allele|Finding|false|false||epo
null|EPX gene|Finding|false|false||epo
null|TIMP1 gene|Finding|false|false||epo
null|Exclusive Provider Organization Plan|Finding|false|false||eponull|Esperanto Language|Entity|false|false||eponull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Agreement|Finding|false|false||accordnull|Amorphous Calcium Carbonate|Drug|false|false||ACC
null|Acetyl-CoA Carboxylase 1|Drug|false|false||ACC
null|Acetyl-CoA Carboxylase 1|Drug|false|false||ACCnull|Agenesis of corpus callosum|Disorder|false|false||ACC
null|Aplasia Cutis Congenita|Disorder|false|false||ACC
null|Adrenocortical carcinoma|Disorder|false|false||ACCnull|ACACA wt Allele|Finding|false|false||ACC
null|ACACA gene|Finding|false|false||ACCnull|Gray matter of anterior cingulate gyrus|Anatomy|false|false||ACC
null|Structure of forceps minor|Anatomy|false|false||ACCnull|acetohydroxamic acid|Drug|false|false||AHA
null|acetohydroxamic acid|Drug|false|false||AHAnull|Factor 8 deficiency, acquired|Disorder|false|false||AHA
null|Autoimmune hemolytic anemia|Disorder|false|false||AHAnull|American Hospital Association|Entity|false|false||AHAnull|Guidelines|Finding|false|false||guidelines
null|Guideline (Publication Type)|Finding|false|false||guidelines
null|guiding characteristics|Finding|false|false||guidelinesnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Additional|Finding|false|false||additionalnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Limited (extensiveness)|Finding|false|false||limitsnull|Use of|Finding|false|false||use ofnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|clonidine|Drug|false|false||clonidine
null|clonidine|Drug|false|false||clonidinenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Transthoracic echocardiography|Procedure|false|false||TTEnull|null|Time|false|false||priornull|Hypokinesia|Finding|false|false||hypokinesisnull|Multiplexed Ion Beam Imaging|Procedure|false|false||MIBInull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Pharmacological stress|Phenomenon|false|false||pharmacological stressnull|pharmacological|Finding|false|false||pharmacologicalnull|Pharmacology|Title|false|false||pharmacologicalnull|Exercise stress test|Procedure|false|false||stress test
null|Stress Test|Procedure|false|false||stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|Urinary Retention|Finding|false|false||urinary retentionnull|Bladder retention of urine|Attribute|false|false||urinary retentionnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Retention of content|Finding|false|false||retention
null|cellular entity retention|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Incontinence|Disorder|false|false||incontinencenull|Diuresis|Finding|false|false||diuresisnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Outpatient visits|Procedure|false|false||outpatient visitsnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Visit|Finding|false|false||visitsnull|Patient Visit|Procedure|false|false||visitsnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|Full|Modifier|false|false||Fullnull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|husband|Subject|false|false||husbandnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Calcitriol Drug Class|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|Calcitriol Drug Class|Drug|false|false||Calcitriolnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Calcitriol Drug Class|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|calcitriol|Drug|false|false||Calcitriol
null|Calcitriol Drug Class|Drug|false|false||Calcitriolnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|sliding scale|Procedure|false|false||Sliding Scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||Scale
null|Base Number|Finding|false|false||Scale
null|Scale - rank|Finding|false|false||Scalenull|Integumentary scale|Anatomy|false|false||Scalenull|Weight measurement scales|Device|false|false||Scalenull|Scaling|Event|false|false||Scalenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Acute on chronic diastolic heart failure|Disorder|false|false||Acute on chronic diastolic congestive heart failurenull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic diastolic heart failure|Disorder|false|false||chronic diastolic congestive heart failurenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|diastolic congestive heart failure|Disorder|false|false||diastolic congestive heart failurenull|Diastole|Attribute|false|false||diastolicnull|Congestive heart failure|Disorder|false|false||congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis|Procedure|false|false||DIAGNOSESnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|null|Time|false|false||priornull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|chronic kidney disease stage|Finding|false|false||Chronic Kidney Disease stagenull|Chronic Kidney Diseases|Disorder|false|false||Chronic Kidney Diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false||Kidney Diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||Kidney
null|Benign neoplasm of kidney|Disorder|false|false||Kidneynull|Kidney problem|Finding|false|false||Kidneynull|examination of kidney|Procedure|false|false||Kidney
null|Procedures on Kidney|Procedure|false|false||Kidneynull|Kidney|Anatomy|false|false||Kidney
null|Both kidneys|Anatomy|false|false||Kidneynull|null|Attribute|false|false||Disease stage
null|disease stage|Attribute|false|false||Disease stagenull|Disease|Disorder|false|false||Diseasenull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Coronary Artery Disease|Disorder|false|false||Coronary Artery Disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary Artery Diseasenull|Coronary artery|Anatomy|false|false||Coronary Arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||Artery Diseasenull|Arterial system|Anatomy|false|false||Artery
null|Arteries|Anatomy|false|false||Arterynull|Disease|Disorder|false|false||Diseasenull|Drug-Eluting Stents|Device|false|false||drug eluting stentnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|null|Device|false|false||stentnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes Mellitus Type 2null|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Type 2|Finding|false|false||Type 2null|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Disease Controlled|Finding|false|false||controlled
null|Control function|Finding|false|false||controlled
null|Controlled mark|Finding|false|false||controllednull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Weight Gain|Finding|false|false||weight gain
null|Gaining Weight question|Finding|false|false||weight gainnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Gain|LabModifier|false|false||gainnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Exacerbation|Finding|false|false||exacerbationnull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Salty|Modifier|false|false||saltynull|Food|Drug|false|false||foodsnull|Holidays|Event|false|false||holidaynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Diuretics|Drug|false|false||diureticsnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Pneumonia|Disorder|false|false||pneumonianull|Plain chest X-ray|Procedure|false|false||chest x-raynull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||x-ray
null|roentgenographic|Finding|false|false||x-raynull|Plain x-ray|Procedure|false|false||x-ray
null|Diagnostic radiologic examination|Procedure|false|false||x-ray
null|Radiographic imaging procedure|Procedure|false|false||x-raynull|Roentgen Rays|Phenomenon|false|false||x-raynull|Language Ability - Sign|Finding|true|false||sign
null|Physical findings|Finding|true|false||signnull|Pneumonia|Disorder|false|false||pneumonianull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Blood Clot|Finding|false|false||clotsnull|Leg|Anatomy|false|false||legsnull|null|Attribute|false|false||legsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Continuous|Finding|false|false||continuenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|salt intake|Subject|false|false||salt intakenull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|gram|LabModifier|false|false||gramsnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Physicians|Subject|false|false||doctorsnull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|Track (course)|Device|false|false||tracknull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|Continuous|Finding|false|false||continuenull|Every morning|Time|false|false||every morningnull|Morning|Time|false|false||morningnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Blood Glucose|Drug|false|false||blood sugarnull|Blood glucose measurement|Procedure|false|false||blood sugarnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|raw sugar|Drug|false|false||sugar
null|raw sugar|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Sugars|Drug|false|false||sugar
null|Carbohydrates|Drug|false|false||sugarnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Hospitalization|Procedure|false|false||Inpatient Carenull|Referral category - Inpatient|Finding|false|false||Inpatient
null|Patient Class - Inpatient|Finding|false|false||Inpatientnull|inpatient encounter|Procedure|false|false||Inpatientnull|inpatient|Subject|false|false||Inpatientnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions