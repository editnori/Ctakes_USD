 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|170,179|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|170,179|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|170,179|false|false|false|C0020517|Hypersensitivity|Allergies
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|182,193|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|182,193|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|182,193|false|false|false|C0030842|penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|182,193|false|false|false|||Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|182,193|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|196,204|false|false|false|C0699512|Dilantin|Dilantin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|196,204|false|false|false|C0699512|Dilantin|Dilantin
Drug|Organic Chemical|SIMPLE_SEGMENT|215,221|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|215,221|false|false|false|C0206046|Zofran|Zofran
Drug|Inorganic Chemical|SIMPLE_SEGMENT|226,239|false|false|false|C1512523|hydrochloride|hydrochloride
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|226,239|false|false|false|C1512523|hydrochloride|hydrochloride
Event|Event|SIMPLE_SEGMENT|243,252|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|243,252|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|261,276|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|267,276|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|267,276|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|267,276|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Functional Concept|SIMPLE_SEGMENT|278,283|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|278,287|false|false|false|C0524470|Right hip region structure|Right hip
Finding|Sign or Symptom|SIMPLE_SEGMENT|278,292|false|false|false|C2202100|Pain of right hip joint|Right hip pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|284,287|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|284,287|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|284,287|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|284,287|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|284,292|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|284,292|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|288,292|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|288,292|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|288,292|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|288,292|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|SIMPLE_SEGMENT|296,301|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|302,310|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|302,310|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|314,332|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|323,332|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|323,332|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|323,332|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|323,332|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|323,332|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|342,349|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|342,349|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|342,349|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|342,349|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|342,352|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|342,368|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|342,368|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|353,360|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|353,360|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|353,368|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|361,368|true|false|false|C0221423|Illness (finding)|Illness
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|399,402|true|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|399,402|true|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|399,402|true|false|false|||CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|404,408|true|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|404,408|true|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|404,408|true|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|SIMPLE_SEGMENT|417,432|true|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|417,432|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|417,432|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|417,432|true|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Finding|SIMPLE_SEGMENT|434,440|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|434,440|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|450,459|true|false|false|C0002395|Alzheimer's Disease|Alzheimer
Event|Event|SIMPLE_SEGMENT|450,459|true|false|false|||Alzheimer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|450,470|true|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|462,470|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|462,470|false|false|false|||dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|473,485|false|false|false|C0029456|Osteoporosis|osteoporosis
Event|Event|SIMPLE_SEGMENT|473,485|false|false|false|||osteoporosis
Finding|Finding|SIMPLE_SEGMENT|473,485|false|false|false|C2911643|Encounter due to family history of osteoporosis|osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|487,490|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|487,490|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|496,504|false|false|false|||presents
Procedure|Health Care Activity|SIMPLE_SEGMENT|510,525|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|SIMPLE_SEGMENT|519,525|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|519,525|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|SIMPLE_SEGMENT|526,534|false|false|false|C4695111|ADMIN.FACILITY|facility
Anatomy|Body Location or Region|SIMPLE_SEGMENT|541,546|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|543,546|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|543,546|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|543,546|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|543,546|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|543,551|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|543,551|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|547,551|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|547,551|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|547,551|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|547,551|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|558,565|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|558,569|false|false|false|C0332310|Has patient|patient has
Finding|Finding|SIMPLE_SEGMENT|570,576|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|570,576|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|570,585|false|false|false|C3494652|Severe dementia|severe dementia
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|577,585|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|577,585|false|false|false|||dementia
Finding|Mental Process|SIMPLE_SEGMENT|592,609|false|false|false|C0025265|Memory, Short-Term|short term memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|592,614|false|false|false|C0701811|Poor short-term memory|short term memory loss
Finding|Idea or Concept|SIMPLE_SEGMENT|598,602|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|598,602|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Finding|SIMPLE_SEGMENT|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|603,609|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|603,614|false|false|false|C0002622|Amnesia|memory loss
Finding|Sign or Symptom|SIMPLE_SEGMENT|603,614|false|false|false|C0751295|Memory Loss|memory loss
Event|Event|SIMPLE_SEGMENT|610,614|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|610,614|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|SIMPLE_SEGMENT|622,628|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|622,628|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|632,639|false|false|false|||provide
Event|Event|SIMPLE_SEGMENT|640,647|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|640,647|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|649,653|false|false|false|||Much
Finding|Finding|SIMPLE_SEGMENT|649,653|false|false|false|C4281574|Much|Much
Event|Event|SIMPLE_SEGMENT|661,668|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|661,668|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|672,680|false|false|false|||obtained
Finding|Classification|SIMPLE_SEGMENT|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|696,702|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Classification|SIMPLE_SEGMENT|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|742,748|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|766,771|false|false|false|||close
Finding|Finding|SIMPLE_SEGMENT|766,771|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|766,771|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|SIMPLE_SEGMENT|783,791|false|false|false|||involved
Event|Activity|SIMPLE_SEGMENT|811,815|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|811,815|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|811,815|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|811,815|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|827,833|false|false|false|||called
Procedure|Health Care Activity|SIMPLE_SEGMENT|843,858|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|SIMPLE_SEGMENT|852,858|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|852,858|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|SIMPLE_SEGMENT|859,867|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Body Substance|SIMPLE_SEGMENT|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|891,898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|910,915|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|910,919|false|false|false|C0524470|Right hip region structure|right hip
Finding|Sign or Symptom|SIMPLE_SEGMENT|910,924|false|false|false|C2202100|Pain of right hip joint|right hip pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|916,919|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|916,919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|916,919|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|916,919|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|916,924|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|916,924|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|920,924|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|920,924|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|920,924|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|920,924|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|932,940|false|false|false|||occurred
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|954,960|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|954,960|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|954,960|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|965,973|true|false|false|||reported
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|974,979|true|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|974,979|true|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|974,979|true|false|false|C0085639|Falls|falls
Event|Event|SIMPLE_SEGMENT|994,1005|true|false|false|||complaining
Event|Event|SIMPLE_SEGMENT|1015,1023|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1015,1023|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|1015,1023|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|1033,1040|false|false|false|||brought
Event|Event|SIMPLE_SEGMENT|1054,1064|false|false|false|||Discussing
Finding|Body Substance|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1087,1092|false|false|false|||moved
Procedure|Health Care Activity|SIMPLE_SEGMENT|1102,1117|false|false|false|C1456630|Assisted Living|Assisted living
Event|Event|SIMPLE_SEGMENT|1111,1117|false|false|false|||living
Finding|Conceptual Entity|SIMPLE_SEGMENT|1111,1117|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|1111,1117|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Event|Event|SIMPLE_SEGMENT|1119,1127|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|1119,1127|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|SIMPLE_SEGMENT|1148,1157|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|1148,1157|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1166,1174|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|1166,1174|false|false|false|||dementia
Event|Event|SIMPLE_SEGMENT|1197,1204|false|false|false|||bowling
Event|Event|SIMPLE_SEGMENT|1221,1227|false|false|false|||social
Finding|Functional Concept|SIMPLE_SEGMENT|1221,1227|false|false|false|C0728831|Social|social
Event|Event|SIMPLE_SEGMENT|1249,1258|false|false|false|||developed
Finding|Intellectual Product|SIMPLE_SEGMENT|1259,1264|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|1265,1268|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1265,1268|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|1274,1284|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1274,1284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|1274,1284|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|SIMPLE_SEGMENT|1296,1305|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1296,1305|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|1327,1332|false|false|false|||noted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1343,1347|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1343,1347|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Intellectual Product|SIMPLE_SEGMENT|1359,1363|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|SIMPLE_SEGMENT|1369,1377|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|1378,1382|false|false|false|||stay
Event|Event|SIMPLE_SEGMENT|1383,1394|false|false|false|||complicated
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1402,1405|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|1402,1405|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|1406,1412|false|false|false|||course
Finding|Functional Concept|SIMPLE_SEGMENT|1420,1428|false|false|false|C0700624|Allergic|allergic
Finding|Pathologic Function|SIMPLE_SEGMENT|1420,1437|false|false|false|C0020517;C1527304|Allergic Reaction;Hypersensitivity|allergic reaction
Event|Event|SIMPLE_SEGMENT|1429,1437|false|false|false|||reaction
Finding|Functional Concept|SIMPLE_SEGMENT|1429,1437|false|false|false|C0443286|Reaction|reaction
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1443,1453|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|1443,1453|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|1443,1453|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Classification|SIMPLE_SEGMENT|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1455,1461|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|1463,1469|false|false|false|||thinks
Drug|Organic Chemical|SIMPLE_SEGMENT|1470,1476|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1470,1476|false|false|false|C0206046|Zofran|Zofran
Event|Event|SIMPLE_SEGMENT|1485,1494|false|false|false|||returning
Event|Event|SIMPLE_SEGMENT|1505,1520|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|1505,1520|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1548,1556|true|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1548,1556|true|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1548,1556|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|1565,1577|true|false|false|||deteriorated
Event|Event|SIMPLE_SEGMENT|1594,1598|false|false|false|||much
Finding|Finding|SIMPLE_SEGMENT|1594,1598|false|false|false|C4281574|Much|much
Finding|Finding|SIMPLE_SEGMENT|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1606,1610|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|SIMPLE_SEGMENT|1611,1621|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Finding|Finding|SIMPLE_SEGMENT|1611,1627|false|false|false|C0558195|Wheelchair bound|wheelchair bound
Event|Activity|SIMPLE_SEGMENT|1622,1627|false|false|false|C1145667|Binding action|bound
Event|Event|SIMPLE_SEGMENT|1622,1627|false|false|false|||bound
Finding|Conceptual Entity|SIMPLE_SEGMENT|1622,1627|false|false|false|C2349209;C2825311|Bound (value);XML Bound|bound
Event|Event|SIMPLE_SEGMENT|1634,1648|false|false|false|||deconditioning
Event|Event|SIMPLE_SEGMENT|1659,1668|false|false|false|||worsening
Finding|Finding|SIMPLE_SEGMENT|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|1669,1675|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|1669,1684|false|false|false|C0025260|Memory|memory function
Event|Event|SIMPLE_SEGMENT|1676,1684|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|1676,1684|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|SIMPLE_SEGMENT|1695,1701|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1695,1701|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|1708,1712|false|false|false|||term
Finding|Idea or Concept|SIMPLE_SEGMENT|1708,1712|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|1708,1712|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Finding|SIMPLE_SEGMENT|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|1714,1720|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1714,1725|false|false|false|C0002622|Amnesia|memory loss
Finding|Sign or Symptom|SIMPLE_SEGMENT|1714,1725|false|false|false|C0751295|Memory Loss|memory loss
Event|Event|SIMPLE_SEGMENT|1721,1725|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1721,1725|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Sign or Symptom|SIMPLE_SEGMENT|1727,1745|false|false|false|C0232462|Decrease in appetite|Decreased appetite
Event|Event|SIMPLE_SEGMENT|1737,1745|false|false|false|||appetite
Finding|Organism Function|SIMPLE_SEGMENT|1737,1745|false|false|false|C0003618|Desire for food|appetite
Event|Event|SIMPLE_SEGMENT|1753,1759|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|1753,1759|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|1753,1759|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|1779,1783|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|1809,1812|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1809,1812|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|SIMPLE_SEGMENT|1809,1822|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1809,1822|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1813,1822|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|1813,1822|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|1813,1822|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|1813,1822|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1813,1822|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1826,1829|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1826,1829|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|1849,1852|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1849,1852|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|SIMPLE_SEGMENT|1877,1885|false|false|false|||evaluate
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1891,1899|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|1900,1908|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|1900,1908|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Idea or Concept|SIMPLE_SEGMENT|1924,1931|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1932,1938|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1978,1982|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1978,1982|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1978,1982|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1987,1998|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|1987,1998|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2005,2010|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2007,2010|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2007,2010|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|2007,2010|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2007,2010|false|false|false|C1292890|Procedure on hip|hip
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2011,2014|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|2011,2014|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|2011,2014|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|2011,2014|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2015,2033|false|false|false|C0223865|Structure of greater trochanter of femur|greater trochanter
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2023,2033|false|false|false|C0162370|Trochanter|trochanter
Finding|Finding|SIMPLE_SEGMENT|2035,2038|false|false|false|C5848551|Neg - answer|neg
Finding|Social Behavior|SIMPLE_SEGMENT|2039,2047|false|false|false|C0019421|Heterosexuality|straight
Finding|Finding|SIMPLE_SEGMENT|2039,2057|false|true|false|C0422926|Straight leg raise test response|straight leg raise
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2048,2051|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|2052,2057|false|false|false|||raise
Drug|Food|SIMPLE_SEGMENT|2064,2070|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2064,2070|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2064,2070|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2064,2070|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|2074,2077|false|false|false|||LLE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2081,2086|false|true|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2081,2086|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2081,2086|false|true|false|C0013604|Edema|edema
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2088,2095|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|2088,2095|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|2088,2095|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2096,2104|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Event|Event|SIMPLE_SEGMENT|2096,2104|false|false|false|||duration
Event|Event|SIMPLE_SEGMENT|2105,2109|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2105,2109|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|2115,2126|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|2115,2126|false|false|false|C0750502|Significant|significant
Anatomy|Cell Component|SIMPLE_SEGMENT|2148,2151|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|2148,2151|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2148,2151|false|false|false|C0009555|Complete Blood Count|CBC
Anatomy|Cell|SIMPLE_SEGMENT|2176,2179|false|false|false|C0023516|Leukocytes|WBC
Finding|Finding|SIMPLE_SEGMENT|2184,2192|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|2184,2192|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|SIMPLE_SEGMENT|2193,2198|false|false|false|||leuks
Finding|Classification|SIMPLE_SEGMENT|2200,2208|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2200,2208|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2200,2208|false|false|false|C5237010|Expression Negative|negative
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2209,2217|false|false|false|C0028137|Nitrites|nitrites
Event|Event|SIMPLE_SEGMENT|2209,2217|false|false|false|||nitrites
Event|Event|SIMPLE_SEGMENT|2220,2227|false|false|false|||Studies
Procedure|Research Activity|SIMPLE_SEGMENT|2220,2227|false|false|false|C0947630|Scientific Study|Studies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2230,2235|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|SIMPLE_SEGMENT|2230,2235|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2230,2245|false|false|false|C0023216|Lower Extremity|Lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2236,2245|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|2246,2256|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|2246,2256|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2246,2256|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2246,2256|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2261,2265|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2261,2270|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2261,2281|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2266,2270|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|2266,2281|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|2271,2281|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2271,2281|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|2289,2293|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|2295,2301|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|2295,2301|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2295,2314|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2302,2309|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2302,2314|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2310,2314|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|2315,2324|false|false|false|||extending
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2343,2352|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2343,2357|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2353,2357|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|SIMPLE_SEGMENT|2360,2364|true|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2360,2369|true|false|false|C0489800|Posterior part of left leg|Left calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2365,2369|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2365,2369|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2370,2375|true|false|false|C0042449|Veins|veins
Event|Event|SIMPLE_SEGMENT|2370,2375|true|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2370,2375|true|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|2393,2403|true|false|false|||identified
Finding|Finding|SIMPLE_SEGMENT|2408,2416|true|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|2423,2431|true|false|false|||occluded
Finding|Finding|SIMPLE_SEGMENT|2423,2431|true|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|2423,2431|true|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2439,2442|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2439,2442|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2439,2442|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|2439,2442|true|false|false|||DVT
Finding|Functional Concept|SIMPLE_SEGMENT|2450,2455|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2450,2471|true|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2456,2461|true|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|2456,2461|true|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2456,2471|true|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2462,2471|true|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|2474,2477|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2474,2477|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Tissue|SIMPLE_SEGMENT|2488,2495|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2488,2495|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|2488,2505|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|2496,2505|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|2496,2505|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|2507,2512|false|false|false|||large
Finding|Gene or Genome|SIMPLE_SEGMENT|2507,2512|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|2520,2525|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|2520,2525|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|2544,2548|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|2544,2548|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2568,2581|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|2568,2581|true|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|2582,2592|true|false|false|||identified
Event|Event|SIMPLE_SEGMENT|2594,2602|true|false|false|||although
Event|Event|SIMPLE_SEGMENT|2604,2614|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|2604,2614|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2604,2614|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|2618,2625|false|false|false|||limited
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2626,2635|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|2626,2635|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|2626,2635|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|2645,2654|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|2645,2654|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|2666,2671|false|false|false|||given
Event|Event|SIMPLE_SEGMENT|2675,2678|false|false|false|||mEq
Drug|Organic Chemical|SIMPLE_SEGMENT|2693,2703|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2693,2703|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|2693,2710|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2693,2710|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2704,2710|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|2704,2710|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|2704,2710|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2704,2710|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|2716,2722|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|2726,2734|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|2726,2734|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|2726,2734|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|2726,2734|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2768,2773|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2768,2773|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|2768,2773|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|2768,2773|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2775,2782|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|SIMPLE_SEGMENT|2775,2782|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|2775,2782|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|2794,2799|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|2808,2815|false|false|false|||resting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2831,2834|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2831,2834|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|2836,2843|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2836,2843|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2848,2856|false|false|false|||obtained
Finding|Idea or Concept|SIMPLE_SEGMENT|2860,2865|false|false|false|C1552828|Table Frame - above|above
Finding|Classification|SIMPLE_SEGMENT|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2871,2877|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|2891,2897|false|false|false|||sleeps
Finding|Finding|SIMPLE_SEGMENT|2914,2921|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|2917,2921|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|2917,2921|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2917,2921|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2917,2921|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|2930,2933|false|false|false|||DOE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2930,2933|false|false|false|C0231807|Dyspnea on exertion|DOE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2953,2958|true|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|2953,2967|true|false|false|C0011135|Defecation|bowel movement
Event|Event|SIMPLE_SEGMENT|2959,2967|true|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2959,2967|true|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|2982,2988|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|2982,2988|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|2982,2988|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|2982,2991|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2982,2999|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2982,2999|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Event|Event|SIMPLE_SEGMENT|2992,2999|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2992,2999|false|false|false|C0449913|System|systems
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3011,3014|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|3011,3014|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|3011,3014|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|3011,3014|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|SIMPLE_SEGMENT|3021,3027|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|3028,3033|true|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|3028,3033|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|3028,3033|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|3035,3041|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|3035,3041|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|3043,3055|true|false|false|C0028081|Night sweats|night sweats
Event|Event|SIMPLE_SEGMENT|3049,3055|true|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|3049,3055|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|3049,3055|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|3057,3063|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|3064,3072|true|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|3064,3072|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3074,3079|true|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3074,3079|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|3074,3079|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3074,3079|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|3081,3091|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3081,3091|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3081,3091|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|3093,3103|true|false|false|||rhinorrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3093,3103|true|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|SIMPLE_SEGMENT|3107,3117|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|3107,3117|false|false|false|C0700148|Congestion|congestion
Event|Event|SIMPLE_SEGMENT|3119,3125|false|false|false|||Denies
Drug|Organic Chemical|SIMPLE_SEGMENT|3126,3131|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3126,3131|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|3126,3131|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|3126,3131|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|3133,3139|false|false|false|||Denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3141,3147|true|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|3141,3147|true|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3141,3147|true|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|3149,3157|true|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|3149,3157|true|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|3159,3167|true|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|3159,3167|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3159,3167|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|3169,3181|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3169,3181|false|false|false|C0009806|Constipation|constipation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3185,3194|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|3185,3199|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3195,3199|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3195,3199|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3195,3199|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3195,3199|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3205,3212|true|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|3205,3212|true|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|3214,3220|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|3221,3232|true|false|false|||arthralgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|3221,3232|true|false|false|C0003862|Arthralgia|arthralgias
Event|Event|SIMPLE_SEGMENT|3236,3244|true|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|3236,3244|true|false|false|C0231528|Myalgia|myalgias
Finding|Finding|SIMPLE_SEGMENT|3251,3271|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|3256,3263|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|3256,3263|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3256,3263|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3256,3263|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3256,3263|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3256,3271|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3264,3271|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3264,3271|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3264,3271|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3273,3285|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|3273,3285|false|false|false|||Hypertension
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3286,3294|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|SIMPLE_SEGMENT|3286,3294|false|false|false|||Dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3295,3307|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|3295,3307|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|3295,3307|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|3308,3317|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Finding|Mental Process|SIMPLE_SEGMENT|3308,3317|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3308,3323|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3308,3332|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3318,3323|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3324,3332|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|3324,3332|false|false|false|||syndrome
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3333,3345|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3333,3345|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Event|Event|SIMPLE_SEGMENT|3333,3345|false|false|false|||Macrocytosis
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3333,3345|false|false|false|C0684332|Macrocytosis (finding)|Macrocytosis
Event|Event|SIMPLE_SEGMENT|3357,3365|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|3357,3365|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|3357,3365|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|3366,3370|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3366,3374|false|false|false|C0229299|Left ear structure|Left ear
Finding|Sign or Symptom|SIMPLE_SEGMENT|3366,3374|false|false|false|C2127178|left ear symptoms (symptom)|Left ear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3371,3374|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3371,3374|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|SIMPLE_SEGMENT|3371,3374|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|SIMPLE_SEGMENT|3371,3374|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Finding|SIMPLE_SEGMENT|3375,3382|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|3375,3382|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3375,3387|false|false|false|C1384666|hearing impairment|hearing loss
Finding|Finding|SIMPLE_SEGMENT|3375,3387|false|false|false|C0011053;C0018772;C2029884;C3887873|Deafness;Hearing Loss;Partial Hearing Loss;hearing loss by exam|hearing loss
Event|Event|SIMPLE_SEGMENT|3383,3387|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|3383,3387|false|false|false|C5890125|Loss (adaptation)|loss
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3388,3394|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|3388,3394|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3388,3394|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|3400,3412|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|3400,3412|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3400,3412|false|false|false|C0020699|Hysterectomy|hysterectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3413,3419|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|3413,3419|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3413,3419|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|3425,3437|false|false|false|||appendectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3425,3437|false|false|false|C0003611;C0003612|Appendectomy;Appendectomy; for ruptured appendix with abscess or generalized peritonitis|appendectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3438,3444|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3438,3444|false|false|false|C1546481|What subject filter - Status|Status
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3450,3457|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3450,3462|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3450,3470|false|false|false|C0195488|Removal of ovarian cyst|ovarian cyst removal
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3458,3462|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|3458,3462|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|3458,3462|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|3458,3462|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3458,3470|false|false|false|C0742962|Cyst removal|cyst removal
Event|Activity|SIMPLE_SEGMENT|3463,3470|false|false|false|C1883720|Removing (action)|removal
Event|Event|SIMPLE_SEGMENT|3463,3470|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3463,3470|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3471,3479|false|false|false|C0086543|Cataract|Cataract
Finding|Finding|SIMPLE_SEGMENT|3471,3479|false|false|false|C1690964|cataract on exam (physical finding)|Cataract
Finding|Finding|SIMPLE_SEGMENT|3471,3487|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Finding|Intellectual Product|SIMPLE_SEGMENT|3471,3487|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3471,3487|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|Cataract surgery
Event|Event|SIMPLE_SEGMENT|3480,3487|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|3480,3487|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3480,3487|false|false|false|C0543467|Operative Surgical Procedures|surgery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3488,3496|false|false|false|C0017601|Glaucoma|Glaucoma
Event|Event|SIMPLE_SEGMENT|3488,3496|false|false|false|||Glaucoma
Finding|Functional Concept|SIMPLE_SEGMENT|3499,3505|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3499,3513|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|3506,3513|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3506,3513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3506,3513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3506,3513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3519,3525|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3519,3525|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3519,3525|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3519,3525|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3519,3533|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3526,3533|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3526,3533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3526,3533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3526,3533|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|3539,3547|true|false|false|||relevant
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3555,3562|true|false|false|C1705970|Electrical Current|current
Event|Event|SIMPLE_SEGMENT|3563,3572|true|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3563,3572|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|3576,3584|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3576,3584|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3576,3584|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3576,3584|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3576,3589|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3576,3589|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3585,3589|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3585,3589|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3585,3589|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3591,3600|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3601,3605|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3601,3605|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3601,3605|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|SIMPLE_SEGMENT|3622,3627|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3622,3633|false|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|3622,3633|false|false|false|C0150404|Taking vital signs|Vital Signs
Event|Event|SIMPLE_SEGMENT|3628,3633|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|3628,3633|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|3628,3633|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Event|Event|SIMPLE_SEGMENT|3668,3675|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3668,3675|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3668,3675|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|3677,3681|false|false|false|||AOx1
Finding|Gene or Genome|SIMPLE_SEGMENT|3677,3681|false|false|false|C1412433|AOX1 gene|AOx1
Event|Event|SIMPLE_SEGMENT|3683,3691|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|3683,3691|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|3693,3700|false|false|false|||smiling
Finding|Social Behavior|SIMPLE_SEGMENT|3693,3700|false|false|false|C0037363|Smiling|smiling
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3705,3713|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|3705,3713|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|3705,3713|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|SIMPLE_SEGMENT|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3718,3724|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3751,3757|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3751,3757|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3751,3757|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3751,3757|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3758,3767|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3758,3767|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3769,3772|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3769,3772|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3774,3784|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|3785,3790|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3785,3790|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|3792,3796|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|3798,3803|true|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3798,3803|true|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3806,3810|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3806,3810|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|3806,3810|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|SIMPLE_SEGMENT|3806,3817|true|false|false|C2230237|Supple neck|neck supple
Event|Event|SIMPLE_SEGMENT|3811,3817|true|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3811,3817|true|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|3819,3822|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3819,3822|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|3827,3835|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3840,3843|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3840,3843|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3840,3843|true|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3840,3843|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Activity|SIMPLE_SEGMENT|3858,3862|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|3858,3862|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3858,3862|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|3867,3873|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|3867,3873|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3867,3873|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3891,3895|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3891,3895|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3900,3908|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3900,3908|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|3910,3916|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3910,3916|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3921,3926|false|false|false|C0024109|Lung|Lungs
Finding|Finding|SIMPLE_SEGMENT|3928,3936|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|3928,3936|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Organism Function|SIMPLE_SEGMENT|3937,3948|false|false|false|C0004048|Inspiration (function)|inspiratory
Event|Event|SIMPLE_SEGMENT|3949,3955|false|false|false|||effort
Finding|Organism Function|SIMPLE_SEGMENT|3949,3955|false|false|false|C0015264|Exertion|effort
Event|Event|SIMPLE_SEGMENT|3957,3966|false|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|3957,3980|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|SIMPLE_SEGMENT|3967,3973|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3967,3980|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|3974,3980|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3974,3980|false|false|false|C0037709||sounds
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|3997,4002|true|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|4011,4018|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|4011,4018|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|4020,4025|true|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|4020,4025|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|4027,4034|true|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|4027,4034|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4037,4044|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4037,4044|true|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|4037,4044|true|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|4037,4044|true|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4046,4050|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|4046,4050|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4079,4084|true|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|4079,4091|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|4085,4091|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4085,4091|true|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|4092,4099|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4092,4099|true|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|4105,4117|true|false|false|||organomegaly
Finding|Finding|SIMPLE_SEGMENT|4105,4117|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|SIMPLE_SEGMENT|4122,4129|true|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|4133,4141|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|4133,4141|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4159,4162|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|4159,4162|true|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|4159,4162|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|4164,4168|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|4164,4168|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4164,4168|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|4170,4174|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4175,4183|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|4188,4194|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4188,4194|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4188,4194|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4188,4194|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4200,4205|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4200,4205|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4200,4215|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4206,4215|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|4217,4225|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|4217,4225|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|4217,4225|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|SIMPLE_SEGMENT|4231,4235|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4231,4239|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4236,4239|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|4240,4252|false|false|false|||erythematous
Finding|Functional Concept|SIMPLE_SEGMENT|4240,4252|false|false|false|C0332476|erythematous|erythematous
Event|Event|SIMPLE_SEGMENT|4257,4263|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|4267,4276|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4267,4276|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|SIMPLE_SEGMENT|4282,4289|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|4282,4295|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4290,4295|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4290,4295|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4290,4295|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|4304,4309|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4304,4325|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4310,4315|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4310,4315|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4310,4325|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4316,4325|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|4335,4342|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|4335,4342|false|true|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|4335,4342|false|true|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4344,4350|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4344,4357|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4344,4357|false|false|false|C4551518|Venous stasis|venous stasis
Event|Event|SIMPLE_SEGMENT|4351,4357|false|false|false|||stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|4351,4357|false|false|false|C0333138|Stasis|stasis
Event|Event|SIMPLE_SEGMENT|4358,4365|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|4358,4365|false|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|4367,4383|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|4370,4377|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|4370,4383|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4378,4383|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4378,4383|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|4405,4409|false|false|false|||AOx1
Finding|Gene or Genome|SIMPLE_SEGMENT|4405,4409|false|false|false|C1412433|AOX1 gene|AOx1
Event|Event|SIMPLE_SEGMENT|4411,4419|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|4411,4419|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4434,4439|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4434,4439|false|false|false|C2003888|Lower (action)|lower
Event|Event|SIMPLE_SEGMENT|4440,4452|false|false|false|||exteremities
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4459,4465|false|false|false|C0015450|Face|facial
Event|Event|SIMPLE_SEGMENT|4466,4475|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|4466,4475|false|false|false|C0026649|Movement|movements
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Immunologic Factor|SIMPLE_SEGMENT|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4479,4483|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Event|Event|SIMPLE_SEGMENT|4485,4494|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|4485,4494|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4485,4494|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|4485,4494|false|false|false|C2229507|sensory exam|sensation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Immunologic Factor|SIMPLE_SEGMENT|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4506,4510|false|false|false|C0618927;C5239612|Tact;bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|tact
Event|Event|SIMPLE_SEGMENT|4512,4516|false|false|false|||gait
Finding|Finding|SIMPLE_SEGMENT|4512,4516|false|false|false|C0016928|Gait|gait
Event|Event|SIMPLE_SEGMENT|4518,4526|false|false|false|||deferred
Finding|Body Substance|SIMPLE_SEGMENT|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4532,4541|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4532,4541|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4542,4546|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4542,4546|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4542,4546|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|4603,4610|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|4603,4610|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|4603,4610|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|4612,4616|false|false|false|||AOx1
Finding|Gene or Genome|SIMPLE_SEGMENT|4612,4616|false|false|false|C1412433|AOX1 gene|AOx1
Event|Event|SIMPLE_SEGMENT|4618,4626|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|4618,4626|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|4628,4635|false|false|false|||smiling
Finding|Social Behavior|SIMPLE_SEGMENT|4628,4635|false|false|false|C0037363|Smiling|smiling
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4640,4648|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|4640,4648|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|4640,4648|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|SIMPLE_SEGMENT|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|4653,4659|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4686,4692|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4686,4692|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|4686,4692|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|4686,4692|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|4693,4702|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|4693,4702|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4704,4707|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4704,4707|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|SIMPLE_SEGMENT|4726,4735|false|false|false|||irregular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4753,4757|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4753,4757|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|4762,4770|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4762,4770|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|4772,4778|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|4772,4778|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4783,4788|false|false|false|C0024109|Lung|Lungs
Finding|Finding|SIMPLE_SEGMENT|4790,4798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|4790,4798|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Organism Function|SIMPLE_SEGMENT|4799,4810|false|false|false|C0004048|Inspiration (function)|inspiratory
Event|Event|SIMPLE_SEGMENT|4811,4817|false|false|false|||effort
Finding|Organism Function|SIMPLE_SEGMENT|4811,4817|false|false|false|C0015264|Exertion|effort
Event|Event|SIMPLE_SEGMENT|4819,4828|false|false|false|||decreased
Finding|Finding|SIMPLE_SEGMENT|4819,4842|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|SIMPLE_SEGMENT|4829,4835|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4829,4842|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|4836,4842|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4836,4842|false|false|false|C0037709||sounds
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|4854,4859|false|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|4854,4859|false|false|false|||bases
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4861,4864|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|4861,4864|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|4861,4864|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|4866,4870|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|4866,4870|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4866,4870|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|4872,4876|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4877,4885|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|4890,4896|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4890,4896|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4890,4896|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4890,4896|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4902,4907|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4902,4907|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4902,4917|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4908,4917|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|4919,4927|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|4919,4927|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|4919,4927|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|SIMPLE_SEGMENT|4933,4937|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4933,4941|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4938,4941|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|4942,4954|false|false|false|||erythematous
Finding|Functional Concept|SIMPLE_SEGMENT|4942,4954|false|false|false|C0332476|erythematous|erythematous
Event|Event|SIMPLE_SEGMENT|4967,4973|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|4978,4987|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4978,4987|false|false|false|C0030247|Palpation|palpation
Finding|Finding|SIMPLE_SEGMENT|4989,5005|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|4992,4999|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|4992,5005|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5000,5005|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5000,5005|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|SIMPLE_SEGMENT|5014,5019|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5014,5035|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5020,5025|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5020,5025|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5020,5035|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5026,5035|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|SIMPLE_SEGMENT|5046,5053|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5046,5053|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5054,5060|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5054,5067|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|5054,5067|false|false|false|C4551518|Venous stasis|venous stasis
Event|Event|SIMPLE_SEGMENT|5061,5067|false|false|false|||stasis
Finding|Pathologic Function|SIMPLE_SEGMENT|5061,5067|false|false|false|C0333138|Stasis|stasis
Event|Event|SIMPLE_SEGMENT|5068,5075|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5068,5075|false|false|false|C0392747|Changing|changes
Finding|Finding|SIMPLE_SEGMENT|5077,5093|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|5080,5087|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|5080,5093|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5088,5093|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5088,5093|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|SIMPLE_SEGMENT|5116,5120|false|false|false|C1412433|AOX1 gene|AOx1
Procedure|Health Care Activity|SIMPLE_SEGMENT|5145,5154|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|5155,5159|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5155,5159|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Body Substance|SIMPLE_SEGMENT|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5187,5192|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5187,5197|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|SIMPLE_SEGMENT|5194,5197|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5194,5197|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5194,5197|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|5200,5203|true|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|SIMPLE_SEGMENT|5208,5216|true|false|false|C1510439|bacteria aspects|BACTERIA
Drug|Food|SIMPLE_SEGMENT|5222,5227|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|5222,5227|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5222,5227|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5222,5227|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|5222,5227|true|false|false|||YEAST
Event|Event|SIMPLE_SEGMENT|5228,5232|true|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5234,5237|true|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5234,5237|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5234,5237|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|SIMPLE_SEGMENT|5234,5237|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|SIMPLE_SEGMENT|5234,5237|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5234,5237|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|SIMPLE_SEGMENT|5234,5237|true|false|false|||EPI
Finding|Gene or Genome|SIMPLE_SEGMENT|5234,5237|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|SIMPLE_SEGMENT|5234,5237|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5234,5237|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Finding|SIMPLE_SEGMENT|5241,5246|true|false|false|C0558141|Transsexual (finding)|TRANS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5247,5250|true|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5247,5250|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5247,5250|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|SIMPLE_SEGMENT|5247,5250|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|SIMPLE_SEGMENT|5247,5250|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5247,5250|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|SIMPLE_SEGMENT|5247,5250|true|false|false|||EPI
Finding|Gene or Genome|SIMPLE_SEGMENT|5247,5250|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|SIMPLE_SEGMENT|5247,5250|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5247,5250|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|SIMPLE_SEGMENT|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5266,5271|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5266,5278|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5273,5278|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5273,5278|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5273,5278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|5279,5282|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5279,5282|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5283,5290|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|SIMPLE_SEGMENT|5291,5294|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5295,5302|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5295,5302|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|SIMPLE_SEGMENT|5295,5302|false|false|false|||PROTEIN
Finding|Conceptual Entity|SIMPLE_SEGMENT|5295,5302|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5295,5302|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|SIMPLE_SEGMENT|5303,5306|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5303,5306|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5308,5315|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|5308,5315|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5308,5315|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5308,5315|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|SIMPLE_SEGMENT|5316,5319|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5316,5319|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|5320,5326|false|false|false|C0022634|Ketones|KETONE
Event|Event|SIMPLE_SEGMENT|5327,5330|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5327,5330|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5331,5340|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5331,5340|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|SIMPLE_SEGMENT|5341,5344|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5341,5344|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5355,5358|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5355,5358|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5372,5375|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|SIMPLE_SEGMENT|5372,5375|false|false|false|||MOD
Event|Event|SIMPLE_SEGMENT|5390,5393|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5390,5393|false|false|false|C0201617|Primed lymphocyte test|PLT
Event|Event|SIMPLE_SEGMENT|5418,5423|false|false|false|||NEUTS
Finding|Body Substance|SIMPLE_SEGMENT|5430,5436|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|5443,5448|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5453,5456|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|5453,5456|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|5453,5456|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Anatomy|Cell|SIMPLE_SEGMENT|5563,5566|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5573,5576|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5573,5576|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5573,5576|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5583,5586|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5583,5586|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|5583,5586|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|5583,5586|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5583,5586|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|5592,5595|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5592,5595|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5592,5595|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|5602,5605|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5602,5605|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5602,5605|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5602,5605|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5602,5605|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5611,5614|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5611,5614|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5611,5614|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5611,5614|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5611,5614|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5611,5614|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5621,5625|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5621,5625|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|5667,5674|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|5667,5674|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|5667,5674|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5667,5674|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5680,5689|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5680,5689|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5694,5703|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5694,5703|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5736,5742|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|5736,5742|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5763,5770|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|5763,5770|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5763,5770|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5763,5770|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5776,5780|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|5776,5780|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5776,5780|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|5776,5780|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5776,5780|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5797,5803|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|5797,5803|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|5797,5803|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5797,5803|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5809,5818|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|5809,5818|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|5809,5818|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5809,5818|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5824,5832|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|5824,5832|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|5824,5832|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5824,5832|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5843,5846|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5843,5846|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|5843,5846|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|5843,5846|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|5843,5846|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5851,5856|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5851,5860|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5851,5860|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5851,5860|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5857,5860|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5857,5860|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|5857,5860|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|5857,5860|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Event|Event|SIMPLE_SEGMENT|5865,5872|false|false|false|||STUDIES
Procedure|Research Activity|SIMPLE_SEGMENT|5865,5872|false|false|false|C0947630|Scientific Study|STUDIES
Event|Event|SIMPLE_SEGMENT|5882,5885|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5882,5885|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Tissue|SIMPLE_SEGMENT|5897,5904|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5897,5904|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|5897,5914|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|5905,5914|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|5905,5914|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|5916,5921|false|false|false|||large
Finding|Gene or Genome|SIMPLE_SEGMENT|5916,5921|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|5929,5934|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|5929,5934|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|5953,5957|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|5953,5957|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5979,5992|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|5979,5992|true|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|5993,6003|true|false|false|||identified
Event|Event|SIMPLE_SEGMENT|6014,6024|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|6014,6024|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6014,6024|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Functional Concept|SIMPLE_SEGMENT|6029,6036|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|SIMPLE_SEGMENT|6029,6036|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6038,6047|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|6038,6047|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6038,6047|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|6057,6066|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|6057,6066|false|false|false|C0013687|effusion|effusions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6070,6076|true|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6070,6076|true|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6070,6076|true|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|SIMPLE_SEGMENT|6070,6076|true|false|false|C0812455|Pelvis problem|Pelvis
Event|Event|SIMPLE_SEGMENT|6077,6081|true|false|false|||Xray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6077,6081|true|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6077,6081|true|false|false|C0043299|Diagnostic radiologic examination|Xray
Finding|Intellectual Product|SIMPLE_SEGMENT|6095,6100|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6101,6109|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|6101,6109|true|false|false|||fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6113,6124|true|false|false|C0012691|Dislocations|dislocation
Event|Event|SIMPLE_SEGMENT|6113,6124|true|false|false|||dislocation
Event|Event|SIMPLE_SEGMENT|6136,6141|true|false|false|||lytic
Finding|Pathologic Function|SIMPLE_SEGMENT|6136,6141|true|false|false|C0024348|Lysis|lytic
Event|Event|SIMPLE_SEGMENT|6146,6155|true|false|false|||sclerotic
Finding|Functional Concept|SIMPLE_SEGMENT|6146,6155|true|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Finding|Pathologic Function|SIMPLE_SEGMENT|6146,6155|true|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6157,6164|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|6157,6164|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|SIMPLE_SEGMENT|6165,6171|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|6165,6171|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|6165,6171|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|6175,6179|false|false|false|||seen
Finding|Idea or Concept|SIMPLE_SEGMENT|6205,6212|true|false|false|C0376327|International Aspects|foreign
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6205,6217|true|false|false|C0016542|Foreign Bodies|foreign body
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6213,6217|true|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6213,6217|true|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|6213,6217|true|false|false|C1551342|Document Body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6221,6229|false|false|false|C0005847|Blood Vessel|Vascular
Event|Event|SIMPLE_SEGMENT|6231,6245|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|6231,6245|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6231,6245|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Event|Event|SIMPLE_SEGMENT|6250,6255|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6273,6278|false|false|false|C0021853|Intestines|bowel
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|SIMPLE_SEGMENT|6279,6282|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Event|Event|SIMPLE_SEGMENT|6279,6282|false|false|false|||gas
Finding|Gene or Genome|SIMPLE_SEGMENT|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|SIMPLE_SEGMENT|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|SIMPLE_SEGMENT|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|SIMPLE_SEGMENT|6279,6282|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Event|Event|SIMPLE_SEGMENT|6295,6309|false|false|false|||nonobstructive
Event|Event|SIMPLE_SEGMENT|6315,6325|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6315,6325|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6315,6325|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6331,6336|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6337,6345|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|6337,6345|true|false|false|||fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6349,6360|true|false|false|C0012691|Dislocations|dislocation
Event|Event|SIMPLE_SEGMENT|6349,6360|true|false|false|||dislocation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6364,6369|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|SIMPLE_SEGMENT|6364,6369|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6364,6379|false|false|false|C0023216|Lower Extremity|Lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6370,6379|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|6380,6390|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|6380,6390|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6380,6390|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6380,6390|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6395,6399|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6395,6404|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6395,6415|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6400,6404|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|6400,6415|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|6405,6415|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6405,6415|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|6423,6427|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|6428,6434|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|6428,6434|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6428,6447|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6435,6442|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6435,6447|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6443,6447|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|6449,6458|false|false|false|||extending
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6478,6487|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6478,6492|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6488,6492|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|SIMPLE_SEGMENT|6495,6499|true|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6495,6504|true|false|false|C0489800|Posterior part of left leg|Left calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6500,6504|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6500,6504|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6505,6510|true|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6505,6510|true|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|6529,6539|true|false|false|||identified
Finding|Finding|SIMPLE_SEGMENT|6542,6550|true|false|false|C0332149|Possible|possibly
Event|Event|SIMPLE_SEGMENT|6556,6564|false|false|false|||occluded
Finding|Finding|SIMPLE_SEGMENT|6556,6564|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6556,6564|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|6574,6579|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6580,6583|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6580,6583|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6580,6583|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|6580,6583|true|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|6592,6596|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6592,6596|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|SIMPLE_SEGMENT|6604,6613|false|false|false|||DISCHARGE
Finding|Body Substance|SIMPLE_SEGMENT|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|6604,6613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|6604,6613|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6659,6664|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6659,6664|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6659,6664|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|6665,6668|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|6675,6678|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6675,6678|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6675,6678|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6685,6688|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6685,6688|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|6685,6688|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6685,6688|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6694,6697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6694,6697|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|6704,6707|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|6704,6707|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6704,6707|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6704,6707|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6704,6707|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|6713,6716|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6713,6716|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|6713,6716|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|6713,6716|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|6713,6716|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6713,6716|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6723,6727|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6755,6758|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6775,6780|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6775,6780|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6775,6780|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|6775,6788|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6775,6788|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6775,6788|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6781,6788|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|6781,6788|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6781,6788|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|6781,6788|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6781,6788|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6781,6788|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6834,6838|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6834,6838|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6834,6838|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6864,6869|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6864,6869|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6864,6869|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6864,6877|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6870,6877|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|6870,6877|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|6870,6877|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|6870,6877|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6870,6877|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|6883,6890|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|6883,6890|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6883,6890|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6883,6890|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Intellectual Product|SIMPLE_SEGMENT|6916,6921|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|6922,6930|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6922,6937|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|6922,6937|false|false|false|C0489547|Hospital course|Hospital Course
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6968,6971|true|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6968,6971|true|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|6968,6971|true|false|false|||CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6973,6977|true|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|6973,6977|true|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6973,6977|true|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|SIMPLE_SEGMENT|6986,7001|true|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|6986,7001|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|6986,7001|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6986,7001|true|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Finding|SIMPLE_SEGMENT|7003,7009|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7003,7009|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7019,7028|true|false|false|C0002395|Alzheimer's Disease|Alzheimer
Event|Event|SIMPLE_SEGMENT|7019,7028|true|false|false|||Alzheimer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7019,7039|true|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7031,7039|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|7031,7039|false|false|false|||dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7042,7054|false|false|false|C0029456|Osteoporosis|osteoporosis
Event|Event|SIMPLE_SEGMENT|7042,7054|false|false|false|||osteoporosis
Finding|Finding|SIMPLE_SEGMENT|7042,7054|false|false|false|C2911643|Encounter due to family history of osteoporosis|osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7056,7059|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|7056,7059|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|7065,7073|false|false|false|||presents
Procedure|Health Care Activity|SIMPLE_SEGMENT|7079,7094|false|false|false|C1456630|Assisted Living|assisted living
Finding|Conceptual Entity|SIMPLE_SEGMENT|7088,7094|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|7088,7094|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|SIMPLE_SEGMENT|7095,7103|false|false|false|C4695111|ADMIN.FACILITY|facility
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7110,7115|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7112,7115|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7112,7115|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|7112,7115|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7112,7115|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7112,7120|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7112,7120|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7116,7120|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7116,7120|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7116,7120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7116,7120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7122,7127|false|false|false|||found
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7136,7139|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7136,7139|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7136,7139|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Functional Concept|SIMPLE_SEGMENT|7140,7144|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|7145,7151|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|7145,7151|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7145,7164|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7152,7159|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7152,7164|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7160,7164|false|false|false|C0042449|Veins|vein
Finding|Intellectual Product|SIMPLE_SEGMENT|7171,7177|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|7171,7186|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|7178,7186|false|false|false|||overload
Event|Activity|SIMPLE_SEGMENT|7197,7204|false|false|false|C0556656|Meetings|meeting
Event|Event|SIMPLE_SEGMENT|7197,7204|false|false|false|||meeting
Finding|Body Substance|SIMPLE_SEGMENT|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7210,7217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|7222,7232|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|7226,7232|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|7226,7232|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|7235,7243|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|7235,7243|false|false|false|C0679006|Decision|decision
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7256,7266|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|SIMPLE_SEGMENT|7256,7266|false|false|false|C2700061|Transition (action)|transition
Procedure|Health Care Activity|SIMPLE_SEGMENT|7256,7271|false|false|false|C4019071|Transitional Care|transition care
Event|Activity|SIMPLE_SEGMENT|7267,7271|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|7267,7271|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|7267,7271|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7267,7271|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Organic Chemical|SIMPLE_SEGMENT|7275,7282|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7275,7282|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Finding|Mental Process|SIMPLE_SEGMENT|7275,7282|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|7283,7291|false|false|false|||directed
Event|Event|SIMPLE_SEGMENT|7293,7301|false|false|false|||measures
Procedure|Health Care Activity|SIMPLE_SEGMENT|7321,7328|false|false|false|C0085555|Hospice Care|hospice
Event|Occupational Activity|SIMPLE_SEGMENT|7321,7337|false|false|false|C5423046|Purchased Services, Clinical and Biomedical, Home Healthcare, Hospice|hospice services
Event|Event|SIMPLE_SEGMENT|7329,7337|false|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|7329,7337|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|7329,7337|false|false|false|C1704289|Clinical Service|services
Event|Event|SIMPLE_SEGMENT|7341,7350|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7341,7350|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7341,7350|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7385,7388|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Event|SIMPLE_SEGMENT|7385,7388|false|false|false|||CMO
Finding|Classification|SIMPLE_SEGMENT|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|7405,7411|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Activity|SIMPLE_SEGMENT|7412,7419|false|false|false|C0556656|Meetings|meeting
Event|Event|SIMPLE_SEGMENT|7412,7419|false|false|false|||meeting
Event|Event|SIMPLE_SEGMENT|7431,7439|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|7431,7439|false|false|false|C0679006|Decision|decision
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7453,7463|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|SIMPLE_SEGMENT|7453,7463|false|false|false|C2700061|Transition (action)|transition
Procedure|Health Care Activity|SIMPLE_SEGMENT|7453,7468|false|false|false|C4019071|Transitional Care|transition care
Event|Activity|SIMPLE_SEGMENT|7464,7468|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|7464,7468|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|7464,7468|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7464,7468|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7472,7475|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Event|SIMPLE_SEGMENT|7472,7475|false|false|false|||CMO
Event|Event|SIMPLE_SEGMENT|7495,7502|false|false|false|||hospice
Procedure|Health Care Activity|SIMPLE_SEGMENT|7495,7502|false|false|false|C0085555|Hospice Care|hospice
Event|Event|SIMPLE_SEGMENT|7504,7512|false|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|7504,7512|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|7504,7512|false|false|false|C1704289|Clinical Service|services
Event|Event|SIMPLE_SEGMENT|7516,7525|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7516,7525|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7516,7525|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7527,7533|true|false|false|||Family
Finding|Classification|SIMPLE_SEGMENT|7527,7533|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|7527,7533|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|7527,7533|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|7527,7533|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Event|Event|SIMPLE_SEGMENT|7542,7546|true|false|false|||want
Event|Event|SIMPLE_SEGMENT|7557,7563|true|false|false|||active
Event|Event|SIMPLE_SEGMENT|7565,7575|true|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7565,7575|true|false|false|C0087111|Therapeutic procedure|treatments
Drug|Organic Chemical|SIMPLE_SEGMENT|7584,7589|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7584,7589|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|7603,7607|false|false|false|||make
Event|Event|SIMPLE_SEGMENT|7612,7625|false|false|false|||uncomfortable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7633,7645|false|false|false|C0021167|Incontinence|incontinence
Event|Event|SIMPLE_SEGMENT|7633,7645|false|false|false|||incontinence
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Drug|Immunologic Factor|SIMPLE_SEGMENT|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7649,7654|false|false|false|C1456647|Childhood Vaccines|shots
Event|Event|SIMPLE_SEGMENT|7649,7654|false|false|false|||shots
Drug|Organic Chemical|SIMPLE_SEGMENT|7663,7670|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7663,7670|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|7663,7670|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|7675,7684|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|7675,7684|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7675,7684|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7689,7692|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7689,7692|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7689,7692|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|7689,7692|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|7694,7698|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|7694,7698|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|7694,7698|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7694,7698|false|false|false|C1553498|home health encounter|Home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7699,7710|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7699,7710|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7699,7710|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7699,7710|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|7711,7721|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7711,7721|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|7711,7721|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|7723,7732|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7723,7732|false|false|false|C0527316|donepezil|donepezil
Event|Event|SIMPLE_SEGMENT|7723,7732|false|false|false|||donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7723,7746|false|false|false|C3652776|donepezil / memantine|donepezil and Memantine
Drug|Organic Chemical|SIMPLE_SEGMENT|7737,7746|false|false|false|C0025242|memantine|Memantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7737,7746|false|false|false|C0025242|memantine|Memantine
Event|Event|SIMPLE_SEGMENT|7737,7746|false|false|false|||Memantine
Event|Event|SIMPLE_SEGMENT|7753,7762|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|7767,7774|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7767,7774|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|7767,7774|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|7767,7774|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|7784,7794|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|7810,7818|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|7810,7818|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Idea or Concept|SIMPLE_SEGMENT|7828,7836|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|7837,7843|false|false|false|||ISSUES
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7870,7873|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7870,7873|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7870,7873|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|7870,7873|false|false|false|||DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7875,7879|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7875,7884|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7875,7895|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7880,7884|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|7880,7895|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|7885,7895|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|7885,7895|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|7903,7907|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|SIMPLE_SEGMENT|7908,7914|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|7908,7914|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7908,7927|false|false|false|C1275667|Common femoral vein|common femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7915,7922|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7915,7927|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7923,7927|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|7929,7938|false|false|false|||extending
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7957,7966|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7957,7971|false|false|false|C0032652|Structure of popliteal vein|popliteal vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7967,7971|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|7972,7981|false|false|false|||diagnosed
Event|Event|SIMPLE_SEGMENT|7986,7996|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|7986,7996|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7986,7996|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7986,7996|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|8000,8009|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8000,8009|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|8020,8026|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|8020,8026|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|8027,8035|false|false|false|||acquired
Finding|Mental Process|SIMPLE_SEGMENT|8043,8050|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|8055,8065|false|false|false|||immobility
Finding|Finding|SIMPLE_SEGMENT|8055,8065|false|false|false|C0231441|Immobile|immobility
Finding|Body Substance|SIMPLE_SEGMENT|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8074,8081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|8091,8101|false|false|false|||restricted
Event|Event|SIMPLE_SEGMENT|8110,8120|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|8110,8120|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Procedure|Health Care Activity|SIMPLE_SEGMENT|8128,8143|false|false|false|C1456630|Assisted Living|assisted living
Event|Event|SIMPLE_SEGMENT|8137,8143|false|false|false|||living
Finding|Conceptual Entity|SIMPLE_SEGMENT|8137,8143|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|SIMPLE_SEGMENT|8137,8143|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Idea or Concept|SIMPLE_SEGMENT|8163,8168|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|8163,8168|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|SIMPLE_SEGMENT|8169,8172|false|false|false|||due
Finding|Functional Concept|SIMPLE_SEGMENT|8169,8172|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|SIMPLE_SEGMENT|8169,8172|false|false|false|C0678226;C3146286|Due;Due to|due
Event|Event|SIMPLE_SEGMENT|8177,8191|false|false|false|||deconditioning
Event|Event|SIMPLE_SEGMENT|8211,8218|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|8222,8229|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8222,8229|false|false|false|C0728963|Lovenox|Lovenox
Event|Event|SIMPLE_SEGMENT|8235,8244|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|8235,8244|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|8235,8244|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|8235,8244|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8235,8244|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|8258,8270|false|false|false|||discontinued
Finding|Mental Process|SIMPLE_SEGMENT|8278,8285|false|false|false|C0542559|contextual factors|setting
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|8289,8299|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|SIMPLE_SEGMENT|8289,8299|false|false|false|C2700061|Transition (action)|transition
Event|Event|SIMPLE_SEGMENT|8289,8299|false|false|false|||transition
Event|Activity|SIMPLE_SEGMENT|8304,8308|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8304,8308|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8304,8308|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8304,8308|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8312,8315|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Event|SIMPLE_SEGMENT|8312,8315|false|false|false|||CMO
Finding|Idea or Concept|SIMPLE_SEGMENT|8319,8324|false|false|false|C1552828|Table Frame - above|above
Finding|Intellectual Product|SIMPLE_SEGMENT|8330,8335|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8336,8339|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8336,8339|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|8336,8339|false|false|false|||CHF
Finding|Body Substance|SIMPLE_SEGMENT|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8341,8348|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8353,8359|false|false|false|||volume
Finding|Intellectual Product|SIMPLE_SEGMENT|8353,8359|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|8360,8370|false|false|false|||overloaded
Event|Event|SIMPLE_SEGMENT|8374,8386|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|8374,8386|false|false|false|C0449450|Presentation|presentation
Anatomy|Tissue|SIMPLE_SEGMENT|8393,8400|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8393,8400|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|8393,8410|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|8401,8410|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|8401,8410|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|8420,8428|false|false|false|||diuresed
Drug|Organic Chemical|SIMPLE_SEGMENT|8437,8442|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8437,8442|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|8437,8442|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|8444,8448|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8444,8448|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8444,8448|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8444,8448|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|8450,8460|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8450,8460|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8450,8460|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|8465,8474|false|false|false|||continued
Finding|Finding|SIMPLE_SEGMENT|8480,8489|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Event|Event|SIMPLE_SEGMENT|8490,8494|false|false|false|||dose
Finding|Mental Process|SIMPLE_SEGMENT|8503,8510|false|false|false|C0542559|contextual factors|setting
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|8515,8525|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|SIMPLE_SEGMENT|8515,8525|false|false|false|C2700061|Transition (action)|transition
Event|Event|SIMPLE_SEGMENT|8515,8525|false|false|false|||transition
Event|Activity|SIMPLE_SEGMENT|8529,8533|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8529,8533|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8529,8533|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8529,8533|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8537,8540|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Event|SIMPLE_SEGMENT|8537,8540|false|false|false|||CMO
Drug|Organic Chemical|SIMPLE_SEGMENT|8542,8547|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8542,8547|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|8542,8547|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|8552,8564|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|8575,8584|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8575,8584|false|false|false|C0549178|Continuous|continued
Drug|Organic Chemical|SIMPLE_SEGMENT|8588,8598|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8588,8598|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8588,8598|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8603,8610|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8603,8610|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|8603,8610|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|8603,8610|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|8616,8624|true|false|false|||remained
Finding|Finding|SIMPLE_SEGMENT|8625,8636|true|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8628,8636|true|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8633,8636|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8633,8636|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|8633,8636|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|8633,8636|true|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|8633,8636|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|8633,8636|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|8633,8636|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8646,8657|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|8646,8657|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|8646,8657|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|8646,8657|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|8646,8666|true|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|8658,8666|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|8658,8666|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|8658,8666|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|8683,8692|false|false|false|||presented
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8696,8701|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8696,8701|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|8696,8701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8696,8701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|SIMPLE_SEGMENT|8696,8708|false|false|false|C0232201;C2041122|Sinus rhythm|sinus rhythm
Event|Event|SIMPLE_SEGMENT|8702,8708|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|8702,8708|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|8702,8708|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|SIMPLE_SEGMENT|8710,8714|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|8710,8714|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|8710,8714|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|8715,8725|false|false|false|||controlled
Drug|Organic Chemical|SIMPLE_SEGMENT|8730,8740|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8730,8740|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8730,8740|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8742,8752|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8742,8752|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|8742,8752|false|false|false|||Metoprolol
Event|Event|SIMPLE_SEGMENT|8757,8766|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|8782,8786|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|8792,8799|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8792,8799|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|8792,8799|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|8792,8799|false|false|false|C1331418|Comfort|comfort
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8805,8808|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|Hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8805,8808|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|Hip
Finding|Gene or Genome|SIMPLE_SEGMENT|8805,8808|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|Hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8805,8808|false|false|false|C1292890|Procedure on hip|Hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8805,8813|false|false|false|C1716793||Hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8805,8813|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|Hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8809,8813|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8809,8813|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|8819,8824|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8819,8828|false|false|false|C0524470|Right hip region structure|right hip
Finding|Sign or Symptom|SIMPLE_SEGMENT|8819,8833|false|false|false|C2202100|Pain of right hip joint|right hip pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8825,8828|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8825,8828|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|8825,8828|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8825,8828|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8825,8833|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8825,8833|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8829,8833|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8829,8833|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8829,8833|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8829,8833|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|8843,8852|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|8863,8871|false|false|false|||resolved
Finding|Finding|SIMPLE_SEGMENT|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|8879,8883|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|8887,8896|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8887,8896|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8898,8904|true|false|false|C0030797|Pelvis|Pelvic
Event|Event|SIMPLE_SEGMENT|8905,8909|true|false|false|||xray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8905,8909|true|false|false|C0043309|Roentgen Rays|xray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8905,8909|true|false|false|C0043299|Diagnostic radiologic examination|xray
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8923,8931|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|8923,8931|true|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|8941,8948|false|false|false|||treated
Drug|Organic Chemical|SIMPLE_SEGMENT|8954,8961|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8954,8961|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|SIMPLE_SEGMENT|8954,8961|false|false|false|||Tylenol
Event|Event|SIMPLE_SEGMENT|8962,8971|false|false|false|||scheduled
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8976,8980|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8976,8980|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8976,8980|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8976,8980|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|8982,8989|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|8982,8989|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|8982,8989|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9001,9009|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|SIMPLE_SEGMENT|9001,9009|false|false|false|||Dementia
Finding|Gene or Genome|SIMPLE_SEGMENT|9019,9023|false|false|false|C1412433|AOX1 gene|AOx1
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9031,9039|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|9031,9039|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|9031,9039|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|9044,9050|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|9044,9050|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|9052,9059|false|false|false|||members
Event|Event|SIMPLE_SEGMENT|9069,9078|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|9082,9089|false|false|false|C0527315|Aricept|Aricept
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9082,9089|false|false|false|C0527315|Aricept|Aricept
Drug|Organic Chemical|SIMPLE_SEGMENT|9090,9097|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9090,9097|false|false|false|C1330412|Namenda|Namenda
Finding|Idea or Concept|SIMPLE_SEGMENT|9102,9114|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|9150,9158|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9150,9158|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|SIMPLE_SEGMENT|9162,9170|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|9179,9185|false|false|false|||orders
Finding|Intellectual Product|SIMPLE_SEGMENT|9179,9185|false|false|false|C3244315|orders - HL7PublishingDomain|orders
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9191,9195|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9191,9195|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9191,9195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9191,9195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9196,9203|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|9196,9203|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|9196,9203|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|SIMPLE_SEGMENT|9204,9214|false|false|false|||secretions
Finding|Body Substance|SIMPLE_SEGMENT|9204,9214|false|false|false|C0036537|Bodily secretions|secretions
Event|Event|SIMPLE_SEGMENT|9225,9233|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|9225,9233|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|9225,9233|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|SIMPLE_SEGMENT|9248,9258|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9248,9258|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9248,9268|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9248,9268|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9259,9268|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Event|Event|SIMPLE_SEGMENT|9259,9268|false|false|false|||succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9273,9282|false|false|false|C0025242|memantine|Memantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9273,9282|false|false|false|C0025242|memantine|Memantine
Event|Event|SIMPLE_SEGMENT|9273,9282|false|false|false|||Memantine
Drug|Organic Chemical|SIMPLE_SEGMENT|9287,9296|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9287,9296|false|false|false|C0527316|donepezil|donepezil
Event|Event|SIMPLE_SEGMENT|9287,9296|false|false|false|||donepezil
Event|Event|SIMPLE_SEGMENT|9301,9310|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9301,9310|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9301,9310|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|SIMPLE_SEGMENT|9315,9322|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9315,9322|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|9315,9322|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|9315,9322|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|9324,9336|false|false|false|||Continuation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9346,9357|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9346,9357|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9346,9357|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9346,9357|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9374,9381|false|false|false|||decided
Finding|Idea or Concept|SIMPLE_SEGMENT|9385,9394|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|9385,9394|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|9395,9402|false|false|false|||hospice
Procedure|Health Care Activity|SIMPLE_SEGMENT|9395,9402|false|false|false|C0085555|Hospice Care|hospice
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9413,9417|false|false|false|C4255237||form
Event|Event|SIMPLE_SEGMENT|9413,9417|false|false|false|||form
Finding|Functional Concept|SIMPLE_SEGMENT|9413,9417|false|false|false|C1522492|Formation|form
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9419,9422|true|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|9419,9422|true|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|9419,9422|true|false|false|C0011015|daunorubicin|DNR
Event|Event|SIMPLE_SEGMENT|9419,9422|true|false|false|||DNR
Finding|Finding|SIMPLE_SEGMENT|9419,9422|true|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|9419,9422|true|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Event|SIMPLE_SEGMENT|9435,9449|true|false|false|||re-hospitalize
Event|Event|SIMPLE_SEGMENT|9454,9458|true|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|9454,9458|true|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|9454,9458|true|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9460,9463|false|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|9460,9463|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|9460,9463|false|false|false|C0011015|daunorubicin|DNR
Event|Event|SIMPLE_SEGMENT|9460,9463|false|false|false|||DNR
Finding|Finding|SIMPLE_SEGMENT|9460,9463|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|9460,9463|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9469,9472|false|false|false|C0410422|Chronic multifocal osteomyelitis|CMO
Event|Event|SIMPLE_SEGMENT|9469,9472|false|false|false|||CMO
Event|Activity|SIMPLE_SEGMENT|9476,9483|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|9476,9483|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|9476,9483|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9476,9483|false|false|false|C0392367|Physical contact|CONTACT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9485,9488|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|9485,9488|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|9485,9488|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9518,9527|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|9518,9527|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|9518,9527|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Gene or Genome|SIMPLE_SEGMENT|9533,9536|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9544,9555|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9544,9555|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9544,9555|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9544,9555|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|9544,9568|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|9559,9568|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9559,9568|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9587,9597|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9587,9597|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9587,9602|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|9598,9602|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|9598,9602|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|9606,9614|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|9619,9627|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|9619,9627|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|9619,9627|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|9619,9627|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|9632,9642|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9632,9642|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9632,9652|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9632,9652|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|9643,9652|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|9643,9652|false|false|false|||Succinate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9666,9669|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9666,9669|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9666,9669|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9666,9669|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9666,9669|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|9674,9683|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9674,9683|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|SIMPLE_SEGMENT|9703,9710|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9703,9710|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9730,9739|false|false|false|C0527316|donepezil|Donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9730,9739|false|false|false|C0527316|donepezil|Donepezil
Drug|Organic Chemical|SIMPLE_SEGMENT|9757,9767|false|false|false|C0244404|raloxifene|raloxifene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9757,9767|false|false|false|C0244404|raloxifene|raloxifene
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9774,9778|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9774,9778|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9774,9778|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9774,9778|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|9779,9784|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9789,9802|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|9789,9802|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9805,9808|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9805,9808|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|9822,9829|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9822,9829|false|false|false|C1330412|Namenda|Namenda
Event|Event|SIMPLE_SEGMENT|9822,9829|false|false|false|||Namenda
Drug|Organic Chemical|SIMPLE_SEGMENT|9822,9832|false|false|false|C1330412|Namenda|Namenda XR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9822,9832|false|false|false|C1330412|Namenda|Namenda XR
Drug|Organic Chemical|SIMPLE_SEGMENT|9834,9843|false|false|false|C0025242|memantine|MEMAntine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9834,9843|false|false|false|C0025242|memantine|MEMAntine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9851,9855|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9851,9855|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|9851,9855|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|9851,9855|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|9856,9861|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Vitamin|SIMPLE_SEGMENT|9866,9879|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9866,9879|false|false|false|C0201898|Ascorbic acid measurement|Ascorbic Acid
Event|Event|SIMPLE_SEGMENT|9875,9879|false|false|false|||Acid
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|9900,9907|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|9900,9907|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|9900,9907|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9900,9907|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9900,9917|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9900,9917|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9908,9917|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Event|Event|SIMPLE_SEGMENT|9908,9917|false|false|false|||Carbonate
Drug|Organic Chemical|SIMPLE_SEGMENT|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9940,9947|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9940,9949|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9940,9949|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|9955,9959|false|false|false|||UNIT
Drug|Food|SIMPLE_SEGMENT|9974,9978|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Drug|Organic Chemical|SIMPLE_SEGMENT|9974,9978|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Event|Event|SIMPLE_SEGMENT|9974,9978|false|false|false|||Fish
Finding|Gene or Genome|SIMPLE_SEGMENT|9974,9978|false|false|false|C1822711;C3274826|SH3PXD2A gene;SH3PXD2A wt Allele|Fish
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|9974,9978|false|false|false|C0162789|Fluorescent in Situ Hybridization|Fish
Drug|Organic Chemical|SIMPLE_SEGMENT|9974,9982|false|false|false|C0016157|fish oils|Fish Oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9974,9982|false|false|false|C0016157|fish oils|Fish Oil
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Food|SIMPLE_SEGMENT|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Organic Chemical|SIMPLE_SEGMENT|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9979,9982|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Finding|Intellectual Product|SIMPLE_SEGMENT|9984,9989|false|false|false|C1719844|Omega|Omega
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Drug|Organic Chemical|SIMPLE_SEGMENT|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9984,9991|false|false|false|C0015689|omega-3 fatty acids|Omega 3
Event|Event|SIMPLE_SEGMENT|10014,10023|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10014,10023|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10014,10023|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10014,10035|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10024,10035|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10024,10035|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|10024,10035|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10024,10035|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|10040,10049|false|false|false|C0527316|donepezil|Donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10040,10049|false|false|false|C0527316|donepezil|Donepezil
Drug|Organic Chemical|SIMPLE_SEGMENT|10067,10077|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10067,10077|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|10067,10087|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10067,10087|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10078,10087|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|10078,10087|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|10111,10118|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10111,10118|false|false|false|C1330412|Namenda|Namenda
Drug|Organic Chemical|SIMPLE_SEGMENT|10111,10121|false|false|false|C1330412|Namenda|Namenda XR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10111,10121|false|false|false|C1330412|Namenda|Namenda XR
Drug|Organic Chemical|SIMPLE_SEGMENT|10123,10132|false|false|false|C0025242|memantine|MEMAntine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10123,10132|false|false|false|C0025242|memantine|MEMAntine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10140,10144|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10140,10144|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|10140,10144|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|10140,10144|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|10145,10150|false|false|false|||DAILY
Drug|Organic Chemical|SIMPLE_SEGMENT|10155,10168|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10155,10168|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10155,10168|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10155,10168|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Event|Event|SIMPLE_SEGMENT|10180,10183|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|10188,10202|true|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10188,10202|true|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Finding|Gene or Genome|SIMPLE_SEGMENT|10217,10220|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|10228,10238|false|false|false|||secretions
Finding|Body Substance|SIMPLE_SEGMENT|10228,10238|false|false|false|C0036537|Bodily secretions|secretions
Drug|Organic Chemical|SIMPLE_SEGMENT|10243,10254|false|false|false|C0596004|hyoscyamine|Hyoscyamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10243,10254|false|false|false|C0596004|hyoscyamine|Hyoscyamine
Finding|Gene or Genome|SIMPLE_SEGMENT|10271,10274|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|10282,10292|false|false|false|||secretions
Finding|Body Substance|SIMPLE_SEGMENT|10282,10292|false|false|false|C0036537|Bodily secretions|secretions
Event|Event|SIMPLE_SEGMENT|10298,10307|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10298,10307|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10298,10307|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10298,10319|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10298,10319|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10308,10319|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10308,10319|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10308,10319|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|10321,10329|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10321,10329|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|10321,10334|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|10330,10334|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|10330,10334|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|10330,10334|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|10330,10334|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|10337,10345|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|10337,10345|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|10353,10362|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10353,10362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10353,10362|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10353,10372|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10363,10372|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10363,10372|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10363,10372|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10363,10372|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10363,10372|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10374,10391|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10382,10391|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10382,10391|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10382,10391|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10382,10391|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10382,10391|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10411,10415|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10411,10420|false|false|false|C0226514|Structure of deep vein|Deep Vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10411,10431|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep Vein Thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10416,10420|false|false|false|C0042449|Veins|Vein
Finding|Pathologic Function|SIMPLE_SEGMENT|10416,10431|false|false|false|C0042487|Venous Thrombosis|Vein Thrombosis
Event|Event|SIMPLE_SEGMENT|10421,10431|false|false|false|||Thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|10421,10431|false|false|false|C0040053|Thrombosis|Thrombosis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10436,10445|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|10436,10445|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|10436,10445|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10436,10455|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|SIMPLE_SEGMENT|10436,10455|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10446,10455|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10446,10455|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10446,10455|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10446,10455|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10446,10455|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10478,10502|false|false|false|C0018802|Congestive heart failure|Congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10489,10494|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10489,10494|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|10489,10494|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10489,10502|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|10495,10502|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10495,10502|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10504,10510|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10504,10523|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10504,10523|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10504,10523|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10511,10523|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|10511,10523|false|false|false|||fibrillation
Finding|Sign or Symptom|SIMPLE_SEGMENT|10526,10538|false|false|false|C0009806|Constipation|Constipation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10541,10553|false|false|false|C0162429|Malnutrition|Malnutrition
Event|Event|SIMPLE_SEGMENT|10541,10553|false|false|false|||Malnutrition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10556,10568|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|10556,10568|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10571,10580|false|false|false|C0002395|Alzheimer's Disease|Alzheimer
Event|Event|SIMPLE_SEGMENT|10571,10580|false|false|false|||Alzheimer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10571,10591|false|false|false|C0002395|Alzheimer's Disease|Alzheimer's dementia
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10583,10591|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|10583,10591|false|false|false|||dementia
Event|Event|SIMPLE_SEGMENT|10597,10606|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10597,10606|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10597,10606|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10597,10606|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10597,10606|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10607,10616|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10607,10616|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10607,10616|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10607,10616|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10618,10624|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10618,10631|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10618,10631|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10625,10631|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10625,10631|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10633,10641|false|false|false|C0009676|Confusion|Confused
Event|Event|SIMPLE_SEGMENT|10633,10641|false|false|false|||Confused
Finding|Finding|SIMPLE_SEGMENT|10633,10641|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|10633,10641|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Finding|SIMPLE_SEGMENT|10644,10650|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Finding|Idea or Concept|SIMPLE_SEGMENT|10644,10650|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|always
Event|Event|SIMPLE_SEGMENT|10652,10657|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10652,10674|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10652,10674|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10661,10674|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10661,10674|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10661,10674|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10676,10681|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10676,10681|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10676,10681|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10676,10681|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10676,10681|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10686,10697|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10686,10697|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10699,10707|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10699,10707|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10699,10707|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10708,10714|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10708,10714|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10708,10714|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10723,10726|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|10723,10726|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|10723,10726|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|10732,10742|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|10732,10742|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|10756,10766|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|10756,10766|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|10771,10780|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10771,10780|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10771,10780|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10771,10780|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10771,10780|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10771,10793|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10771,10793|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|10771,10793|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10781,10793|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10781,10793|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10781,10793|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|10795,10799|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|10816,10824|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|10816,10824|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|10816,10824|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|10832,10836|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10832,10836|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10832,10836|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10832,10836|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10832,10839|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|10857,10872|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10857,10872|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|10892,10904|false|false|false|||hospitalized
Finding|Functional Concept|SIMPLE_SEGMENT|10910,10915|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10910,10919|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10916,10919|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10916,10919|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|SIMPLE_SEGMENT|10916,10919|false|false|false|||hip
Finding|Gene or Genome|SIMPLE_SEGMENT|10916,10919|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10916,10919|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10921,10925|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10921,10925|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10921,10925|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10921,10925|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10934,10939|false|false|false|||Xrays
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10934,10939|false|false|false|C0043309|Roentgen Rays|Xrays
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10948,10951|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10948,10951|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|SIMPLE_SEGMENT|10948,10951|false|false|false|||hip
Finding|Gene or Genome|SIMPLE_SEGMENT|10948,10951|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10948,10951|false|false|false|C1292890|Procedure on hip|hip
Event|Event|SIMPLE_SEGMENT|10966,10970|true|false|false|||show
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10975,10984|true|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|10975,10984|true|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|10975,10984|true|false|false|C4554413|Fractured|fractures
Event|Event|SIMPLE_SEGMENT|10995,11000|false|false|false|||found
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11003,11008|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|11003,11008|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|11003,11008|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|11003,11013|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|SIMPLE_SEGMENT|11009,11013|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11009,11013|false|false|false|C0009074|clotrimazole|clot
Event|Event|SIMPLE_SEGMENT|11009,11013|false|false|false|||clot
Finding|Pathologic Function|SIMPLE_SEGMENT|11009,11013|false|false|false|C0302148|Blood Clot|clot
Finding|Functional Concept|SIMPLE_SEGMENT|11022,11026|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11022,11030|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11027,11030|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|SIMPLE_SEGMENT|11035,11042|true|false|false|||noticed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11054,11059|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11054,11059|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|11054,11059|true|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|11054,11059|true|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|11067,11074|true|false|false|||pumping
Event|Event|SIMPLE_SEGMENT|11096,11102|false|false|false|||talked
Event|Event|SIMPLE_SEGMENT|11122,11128|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|11122,11128|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|11134,11140|false|false|false|||shared
Event|Event|SIMPLE_SEGMENT|11162,11168|false|false|false|||wishes
Event|Event|SIMPLE_SEGMENT|11182,11194|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|11203,11207|false|false|false|||type
Finding|Gene or Genome|SIMPLE_SEGMENT|11203,11207|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|11203,11207|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Activity|SIMPLE_SEGMENT|11211,11215|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11211,11215|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11211,11215|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11211,11215|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|11247,11254|false|false|false|||decided
Event|Event|SIMPLE_SEGMENT|11258,11263|false|false|false|||focus
Drug|Organic Chemical|SIMPLE_SEGMENT|11272,11279|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11272,11279|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|SIMPLE_SEGMENT|11272,11279|false|false|false|||comfort
Finding|Mental Process|SIMPLE_SEGMENT|11272,11279|false|false|false|C1331418|Comfort|comfort
Event|Event|SIMPLE_SEGMENT|11313,11323|false|false|false|||discharged
Procedure|Health Care Activity|SIMPLE_SEGMENT|11335,11342|false|false|false|C0085555|Hospice Care|hospice
Finding|Finding|SIMPLE_SEGMENT|11335,11347|false|false|false|C0869461|Encounter for Hospice Care|hospice care
Procedure|Health Care Activity|SIMPLE_SEGMENT|11335,11347|false|false|false|C0085555|Hospice Care|hospice care
Event|Activity|SIMPLE_SEGMENT|11343,11347|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11343,11347|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11343,11347|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11343,11347|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Classification|SIMPLE_SEGMENT|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|11374,11380|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|11401,11410|false|false|false|||Treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|11401,11410|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Finding|Functional Concept|SIMPLE_SEGMENT|11401,11410|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11401,11410|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11401,11410|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11419,11427|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11428,11440|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11428,11440|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11428,11440|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

