CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Cardiothoracic|Modifier|false|false||CARDIOTHORACICnull|Dyes|Drug|false|false||Dyenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Contrast Media|Drug|false|false||Contrast Medianull|Contrast Media|Drug|false|false||Contrastnull|Contrast|Modifier|false|false||Contrastnull|Communications Media|Finding|false|false||Media
null|PAMS Media|Finding|false|false||Medianull|Tunica Media|Anatomy|false|false||Media
null|Media layer|Anatomy|false|false||Medianull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|cilostazol|Drug|false|false||cilostazol
null|cilostazol|Drug|false|false||cilostazolnull|varenicline|Drug|false|false||Varenicline
null|varenicline|Drug|false|false||Vareniclinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Intubation (procedure)|Procedure|false|false||Intubationnull|Mechanical ventilation finding|Finding|false|false||Mechanical Ventilationnull|Mechanical ventilation|Procedure|false|false||Mechanical Ventilationnull|mechanical method|Finding|false|false||Mechanicalnull|Mechanical Treatments|Procedure|false|false||Mechanicalnull|Ventilation, function (observable entity)|Finding|false|false||Ventilation
null|Respiration|Finding|false|false||Ventilationnull|Assisted breathing|Procedure|false|false||Ventilationnull|Environmental air flow|Phenomenon|false|false||Ventilationnull|Tracheal Extubation|Procedure|false|false||Extubatednull|EntityNameUseR2 - temporary|Finding|false|false||Temporary
null|Job Status - Temporary|Finding|false|false||Temporarynull|Transitory|Time|false|false||Temporarynull|PACERR gene|Finding|false|false||Pacer
null|RUBCNL gene|Finding|false|false||Pacernull|null|Procedure|false|false||Placement
null|Implantation procedure|Procedure|false|false||Placement
null|Clinical act of insertion|Procedure|false|false||Placementnull|Placement|Modifier|false|false||Placementnull|EZR wt Allele|Finding|false|false||CVL
null|EZR gene|Finding|false|false||CVLnull|Insertion Mutation|Finding|false|false||Insertion
null|Insert (object)|Finding|false|false||Insertionnull|Clinical act of insertion|Procedure|false|false||Insertion
null|Implantation procedure|Procedure|false|false||Insertionnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Atrial Fibrillation|Disorder|false|false||atrial fibrillationnull|null|Attribute|false|false||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Home with services|Finding|false|false||home with servicesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Recent|Time|false|false||recentnull|Severe (severity modifier)|Finding|false|false||severelynull|Reduced forced expiratory volume in one second|Finding|false|false||reduced FEV1null|Pulmonary Function Test/Forced Expiratory Volume 1|Procedure|false|false||FEV1null|null|Attribute|false|false||FEV1null|Volume expired during 1.0 s of forced expiration|LabModifier|false|false||FEV1null|Moderate Response|Finding|false|false||moderately
null|Moderate|Finding|false|false||moderately
null|Moderate Effect|Finding|false|false||moderatelynull|Moderate (severity modifier)|Modifier|false|false||moderately
null|Moderation|Modifier|false|false||moderatelynull|Reduced forced expiratory volume in one second|Finding|false|false||reduced FEV1null|Forced Expiratory Volume in 1 Second to Forced Vital Capacity Ratio Measurement|Procedure|false|false||FEV1/FVCnull|null|Attribute|false|false||FEV1/FVCnull|Pulmonary Function Test/Forced Expiratory Volume 1|Procedure|false|false||FEV1null|null|Attribute|false|false||FEV1null|Volume expired during 1.0 s of forced expiration|LabModifier|false|false||FEV1null|Forced Vital Capacity|Lab|false|false||FVCnull|Psychological Well Being|Finding|false|false||feeling betternull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Presentation|Finding|false|false||presentationnull|Dyspnea|Finding|false|false||short of breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|Exertion|Finding|false|false||exertionnull|Productive Cough|Finding|false|false||cough productivenull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Brown sputum|Finding|false|false||brown sputumnull|Brown Tendon Sheath Syndrome|Disorder|false|false||brownnull|Brown color|Modifier|false|false||brownnull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Pillow|Device|false|false||pillowsnull|Side|Modifier|false|false||sidenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Concern|Finding|false|false||concernnull|Due to|Finding|false|false||due
null|Due|Finding|false|false||duenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Weight-Bearing state|Subject|false|false||weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Bearing Device|Device|false|false||bearingnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Accidental Falls|Disorder|true|false||fallsnull|Falls|Finding|true|false||fallsnull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Numbness|Finding|true|false||loss of sensationnull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Fecal Incontinence|Disorder|false|false||fecal incontinencenull|Feces|Finding|false|false||fecalnull|Incontinence|Disorder|false|false||incontinencenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Specimen Type - Cannula|Finding|false|false||Cannula
null|null|Finding|false|false||Cannulanull|Body Parts - Cannula|Anatomy|false|false||Cannulanull|Cannula device|Device|false|false||Cannulanull|Calamus <grasshoppers>|Entity|false|false||Cannulanull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Diffuse|Modifier|false|false||diffusenull|Worst|Modifier|false|false||worstnull|Radiolucent Lines|Finding|false|false||RLLnull|Structure of right lower lobe of lung|Anatomy|false|false||RLLnull|Tripod|Device|false|false||tripodingnull|Laboratory test finding|Lab|false|false||Labsnull|Influenza|Disorder|false|false||flunull|ZMYND10 wt Allele|Finding|false|false||flunull|Fluorescence Units|LabModifier|false|false||flunull|Swab Dosage Form|Drug|false|false||swab
null|Swab specimen|Drug|false|false||swabnull|Taking of swab|Procedure|false|false||swabnull|Swab|Device|false|false||swabnull|Swab Dosing Unit|LabModifier|false|false||swabnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Leukocytes|Anatomy|false|false||WBCnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|shift displacement|Finding|false|false||shiftnull|Physical Shift|Phenomenon|false|false||shiftnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Cloudy|Modifier|false|false||cloudynull|Proteins|Drug|false|false||protein
null|Proteins|Drug|false|false||proteinnull|Protein Info|Finding|false|false||proteinnull|Protein measurement|Procedure|false|false||proteinnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Plain chest X-ray|Procedure|false|false||CXRnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Atelectasis|Finding|false|false||atelectasisnull|Physicians|Subject|false|false||physiciansnull|Pneumonia|Disorder|false|false||pneumonianull|Lateral|Modifier|false|false||lateralnull|View|Modifier|false|false||viewnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|DuoNeb|Drug|false|false||duoneb
null|DuoNeb|Drug|false|false||duonebnull|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisone
null|prednisone|Drug|false|false||prednisonenull|Total|Modifier|false|false||totalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Consultation|Procedure|false|false||Consultsnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Slightly better|Modifier|false|false||slightly betternull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Breath|Finding|false|false||breathnull|EPRS1 gene|Finding|false|false||earsnull|null|Anatomy|false|false||ears
null|Ear structure|Anatomy|false|false||earsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Asthma|Disorder|false|false||Asthmanull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Atypical chest pain|Finding|false|false||Atypical Chest Painnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false||Chest Painnull|null|Attribute|false|false||Chest Painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Atrial Fibrillation|Disorder|false|false||Atrial Fibrillationnull|null|Attribute|false|false||Atrial Fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Atrial Fibrillationnull|Heart Atrium|Anatomy|false|false||Atrialnull|Fibrillation|Disorder|false|false||Fibrillationnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|Anxiety Disorders|Disorder|false|false||Anxiety
null|Anxiety|Disorder|false|false||Anxietynull|Anxiety symptoms|Finding|false|false||Anxietynull|Cervical radiculitis|Disorder|false|false||Cervical Radiculitisnull|Neck|Anatomy|false|false||Cervicalnull|Cervical|Modifier|false|false||Cervicalnull|Radiculitis|Disorder|false|false||Radiculitisnull|Cervical spondylosis without myelopathy|Disorder|false|false||Cervical Spondylosis
null|Cervical spondylosis|Disorder|false|false||Cervical Spondylosisnull|Neck|Anatomy|false|false||Cervicalnull|Cervical|Modifier|false|false||Cervicalnull|Spondylosis|Disorder|false|false||Spondylosisnull|Coronary Artery Disease|Disorder|false|false||Coronary Artery Disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary Artery Diseasenull|Coronary artery|Anatomy|false|false||Coronary Arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||Artery Diseasenull|Arterial system|Anatomy|false|false||Artery
null|Arteries|Anatomy|false|false||Arterynull|Disease|Disorder|false|false||Diseasenull|Headache|Finding|false|false||Headachenull|Herpes zoster (disorder)|Disorder|false|false||Herpes Zoster
null|herpesvirus 3, human|Disorder|false|false||Herpes Zosternull|Herpes simplex dermatitis|Disorder|false|false||Herpes
null|null|Disorder|false|false||Herpesnull|Herpes <Hyperinae>|Entity|false|false||Herpesnull|Herpes zoster (disorder)|Disorder|false|false||Zosternull|Gastrointestinal Hemorrhage|Finding|false|false||GI Bleedingnull|Hemorrhage|Finding|false|false||Bleedingnull|Peripheral Vascular Diseases|Disorder|false|false||Peripheral Vascular Diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false||Vascular Diseasenull|Blood Vessel|Anatomy|false|false||Vascularnull|Vascular|Modifier|false|false||Vascularnull|Disease|Disorder|false|false||Diseasenull|Bilateral|Modifier|false|false||bilateralnull|iliac stents|Procedure|false|false||iliac stentsnull|Bone structure of ilium|Anatomy|false|false||iliacnull|null|Device|false|false||stentsnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false||hip replacementnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Asthma|Disorder|false|false||asthmanull|Hypertensive disease|Disorder|false|false||hypertensionnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Malignant tumor of colon|Disorder|false|false||colon cancer
null|Malignant neoplasm of large intestine|Disorder|false|false||colon cancer
null|Colon Carcinoma|Disorder|false|false||colon cancernull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|leukemia|Disorder|false|false||leukemianull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Somewhat|Finding|false|false||somewhatnull|Wheezing|Finding|false|false||wheezenull|HEENT|Anatomy|false|false||HEENTnull|Pallor of skin|Finding|true|false||pallornull|Icterus|Finding|true|false||icterusnull|Icterus <Icteridae>|Entity|true|false||icterusnull|null|LabModifier|false|false||icterusnull|Oropharyngeal lesion|Disorder|true|false||oropharyngeal lesionnull|Disorder of oropharynx|Disorder|false|false||oropharyngealnull|Oropharyngeal Route of Administration|Finding|false|false||oropharyngealnull|Oropharyngeal|Anatomy|false|false||oropharyngealnull|Lesion|Finding|true|false||lesion
null|null|Finding|true|false||lesionnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|true|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|true|false||sinusnull|pathologic fistula|Disorder|true|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Unable|Finding|false|false||unablenull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Pulmonary (intended site)|Finding|false|false||PULMONARYnull|Lung|Anatomy|false|false||PULMONARYnull|null|Attribute|false|false||PULMONARYnull|Pulmonary (qualifier value)|Modifier|false|false||PULMONARYnull|Diffuse|Modifier|false|false||diffusenull|Wheezing|Finding|false|false||wheezesnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Edema of lower extremity|Finding|false|false||lower extremity edemanull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false||extremity edemanull|Limb structure|Anatomy|false|false||extremitynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Shin|Anatomy|false|false||shinsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Style|Modifier|false|false||stylenull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Neurologic (qualifier value)|Modifier|false|false||NEUROLOGICnull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|PURPOSE (pharmacologic preparation)|Drug|false|false||purpose
null|PURPOSE (pharmacologic preparation)|Drug|false|false||purposenull|Purpose|Finding|false|false||purposenull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Continuous|Finding|false|false||continuousnull|Telemetry|Procedure|false|false||telemetrynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|vocal|Finding|false|false||vocalnull|CD96 wt Allele|Finding|false|false||tactile
null|CD96 gene|Finding|false|false||tactilenull|Tactile|Modifier|false|false||tactilenull|Stimulus|Phenomenon|false|false||stimulinull|Pupil|Anatomy|false|false||Pupilsnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Respiratory Sounds|Attribute|true|false||lung soundsnull|Lung diseases|Disorder|true|false||lungnull|Lung Problem|Finding|true|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|null|Device|true|false||soundsnull|null|Phenomenon|true|false||soundsnull|1 Minute|LabModifier|false|false||1 minutenull|Minute of time|Time|false|false||minutenull|Minute Unit of Plane Angle|LabModifier|false|false||minute
null|Minute (diminutive)|LabModifier|false|false||minute
null|Small|LabModifier|false|false||minutenull|Auscultation|Procedure|false|false||auscultationnull|Pronounced Dead|Finding|false|false||pronounced deadnull|Dead (finding)|Finding|false|false||dead
null|Death (finding)|Finding|false|false||dead
null|Cessation of life|Finding|false|false||deadnull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|Autopsy|Procedure|false|false||an autopsynull|null|Finding|false|false||autopsynull|Autopsy - Consent type|Procedure|false|false||autopsy
null|Autopsy|Procedure|false|false||autopsynull|Laboratory test finding|Lab|false|false||LABSnull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Natriuretic Peptides B, human|Drug|false|false||proBNP
null|Natriuretic Peptides B, human|Drug|false|false||proBNPnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false||Base
null|Base|Drug|false|false||Base
null|Dental Base|Drug|false|false||Base
null|base - RoleClass|Drug|false|false||Basenull|Base - General Qualifier|Finding|false|false||Base
null|BPIFA4P gene|Finding|false|false||Base
null|Base - RX Component Type|Finding|false|false||Basenull|Anatomical base|Anatomy|false|false||Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Published Comment|Finding|false|false||Comment
null|Comment|Finding|false|false||Commentnull|Green color|Modifier|false|false||GREENnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Laboratory test finding|Lab|false|false||LABSnull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Selenium and Vitamin E Efficacy Trial|Procedure|false|false||SELECTnull|Choose (action)|Event|false|false||SELECTnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|Comparison|Event|false|false||COMPARISONnull|heart size|Finding|false|false||Heart sizenull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Mildly enlarged|Finding|false|false||mildly enlargednull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Chest>Aorta.thoracic|Anatomy|false|false||thoracic aorta
null|Thoracic aorta|Anatomy|false|false||thoracic aortanull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false||thoracicnull|Chest|Anatomy|false|false||thoracicnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|Hilar|Modifier|false|false||hilarnull|Contour form|Modifier|false|false||contoursnull|null|Modifier|false|false||unremarkablenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Atelectasis|Finding|false|false||atelectasisnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pleural Diseases|Disorder|false|false||Pleuralnull|Pleura|Anatomy|false|false||Pleuralnull|Pleural|Modifier|false|false||Pleuralnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Pneumothorax|Disorder|false|false||pneumothoraxnull|Has focus|Finding|false|false||Focusnull|Focal|Modifier|false|false||Focusnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of hemidiaphragm|Anatomy|false|false||hemidiaphragmnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Excision of large intestine for interposition|Procedure|false|false||colonic interpositionnull|Colon structure (body structure)|Anatomy|false|false||colonicnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false||cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false||cardiopulmonarynull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Ruta graveolens preparation|Drug|false|false||RUE
null|Ruta graveolens preparation|Drug|false|false||RUEnull|Ruta graveolens|Entity|false|false||RUE
null|Ruta|Entity|false|false||RUEnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Deep vein thrombosis of lower limb|Disorder|false|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Middle|Modifier|false|false||midnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of brachial vein|Anatomy|false|false||brachial veinnull|Brachial (qualifier value)|Modifier|false|false||brachialnull|Veins|Anatomy|false|false||veinnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Plain chest X-ray|Procedure|false|false||CXRnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Endotracheal tube|Device|false|false||endotracheal tubenull|endotracheal|Modifier|false|false||endotrachealnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|KAT5 wt Allele|Finding|false|false||tip
null|ITFG1 gene|Finding|false|false||tip
null|METTL8 gene|Finding|false|false||tip
null|TIPRL gene|Finding|false|false||tipnull|TIP regimen|Procedure|false|false||tipnull|Device tip (physical object)|Device|false|false||tipnull|Tip|Modifier|false|false||tipnull|Structure of carina|Anatomy|false|false||carina
null|Keel structure|Anatomy|false|false||carinanull|Nasogastric tube procedures|Procedure|false|false||Nasogastric tubenull|Nasogastric tube|Device|false|false||Nasogastric tubenull|Nasogastric Route of Administration|Finding|false|false||Nasogastricnull|Nasogastric|Anatomy|false|false||Nasogastricnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|KAT5 wt Allele|Finding|false|false||tip
null|ITFG1 gene|Finding|false|false||tip
null|METTL8 gene|Finding|false|false||tip
null|TIPRL gene|Finding|false|false||tipnull|TIP regimen|Procedure|false|false||tipnull|Device tip (physical object)|Device|false|false||tipnull|Tip|Modifier|false|false||tipnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|Film Dosage Form|Drug|false|false||film
null|film - layer|Drug|false|false||filmnull|null|Finding|false|false||filmnull|film (photographic)|Device|false|false||film
null|Film Device|Device|false|false||film
null|Film Container Cap|Device|false|false||filmnull|Film (unit of presentation)|LabModifier|false|false||film
null|Film Dosing Unit|LabModifier|false|false||filmnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|null|Device|false|false||central linenull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|KAT5 wt Allele|Finding|false|false||tip
null|ITFG1 gene|Finding|false|false||tip
null|METTL8 gene|Finding|false|false||tip
null|TIPRL gene|Finding|false|false||tipnull|TIP regimen|Procedure|false|false||tipnull|Device tip (physical object)|Device|false|false||tipnull|Tip|Modifier|false|false||tipnull|Middle|Modifier|false|false||midnull|Slow vital capacity|Finding|false|false||SVCnull|null|Finding|false|false||pacemakernull|Artificial cardiac pacemaker|Device|false|false||pacemaker
null|Pacemakers|Device|false|false||pacemakernull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|lead|Drug|false|false||lead
null|Plumbum metallicum, homeopathic preparation|Drug|false|false||lead
null|Plumbum metallicum, homeopathic preparation|Drug|false|false||lead
null|lead|Drug|false|false||leadnull|Leading|Finding|false|false||leadnull|Lead measurement|Procedure|false|false||lead
null|Long Ensemble Angular-Coherence Doppler Ultrasound|Procedure|false|false||leadnull|Lead Device|Device|false|false||leadnull|Right ventricular structure|Anatomy|false|false||right ventriclenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Heart Ventricle|Anatomy|false|false||ventricle
null|Cerebral Ventricles|Anatomy|false|false||ventricle
null|Ventricle|Anatomy|false|false||ventriclenull|Probable diagnosis|Finding|false|false||probablenull|Probability|LabModifier|false|false||probablenull|Cicatrization|Finding|false|false||scarring
null|Cicatrix|Finding|false|false||scarringnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|Areas <Spilosomini>|Entity|true|false||areasnull|Area|Modifier|false|false||areasnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Zone|Modifier|false|false||zonenull|Redistribution|Finding|false|false||redistributionnull|Cardiomegaly|Finding|false|false||cardiomegalynull|Pulmonary venous hypertension|Finding|false|false||pulmonary venous hypertensionnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Venous hypertension|Disorder|false|false||venous hypertensionnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Atrial Fibrillation|Disorder|false|false||AFibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||AFibnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Recent|Time|false|false||recentnull|Hospitalization|Procedure|false|false||hospitalizationsnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Last|Modifier|false|false||lastnull|Several|LabModifier|false|false||severalnull|month|Time|false|false||monthsnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Wheezing|Finding|false|false||wheezingnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Steroids|Drug|false|false||steroids
null|Steroids|Drug|false|false||steroidsnull|Pisum sativum (pea) extract|Drug|false|false||PEA
null|null|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|Pisum sativum (pea) extract|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|palmidrol|Drug|false|false||PEAnull|Electromechanical dissociation|Disorder|false|false||PEAnull|area PEa of Pandya|Anatomy|false|false||PEAnull|Pisum sativum|Entity|false|false||PEAnull|Cardiac Arrest|Disorder|false|false||arrestnull|Encounter due to problems related to other legal circumstances - arrest|Finding|false|false||arrestnull|Law enforcement arrest|Event|false|false||arrestnull|Arrested progression|Time|false|false||arrestnull|Thought|Finding|false|false||thought
null|null|Finding|false|false||thoughtnull|Hypoxemia|Finding|false|false||hypoxemia
null|Blood oxygen concentration below reference range (finding)|Finding|false|false||hypoxemianull|Intubation, Intratracheal|Procedure|false|false||endotracheal intubationnull|endotracheal|Modifier|false|false||endotrachealnull|Intubation (procedure)|Procedure|false|false||intubationnull|Mechanical ventilation finding|Finding|false|false||mechanical ventilationnull|Mechanical ventilation|Procedure|false|false||mechanical ventilationnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Ventilation, function (observable entity)|Finding|false|false||ventilation
null|Respiration|Finding|false|false||ventilationnull|Assisted breathing|Procedure|false|false||ventilationnull|Environmental air flow|Phenomenon|false|false||ventilationnull|temporary pacemaker|Device|false|false||temporary pacemakernull|EntityNameUseR2 - temporary|Finding|false|false||temporary
null|Job Status - Temporary|Finding|false|false||temporarynull|Transitory|Time|false|false||temporarynull|null|Finding|false|false||pacemakernull|Artificial cardiac pacemaker|Device|false|false||pacemaker
null|Pacemakers|Device|false|false||pacemakernull|Menstruation|Finding|false|false||periodsnull|Bradycardia by ECG Finding|Finding|false|false||bradycardia
null|Bradycardia|Finding|false|false||bradycardianull|Pisum sativum (pea) extract|Drug|false|false||PEA
null|null|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|Pisum sativum (pea) extract|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|palmidrol|Drug|false|false||PEAnull|Electromechanical dissociation|Disorder|false|false||PEAnull|area PEa of Pandya|Anatomy|false|false||PEAnull|Pisum sativum|Entity|false|false||PEAnull|Cardiac Arrest|Disorder|false|false||arrestnull|Encounter due to problems related to other legal circumstances - arrest|Finding|false|false||arrestnull|Law enforcement arrest|Event|false|false||arrestnull|Arrested progression|Time|false|false||arrestnull|Manifestation of|Modifier|false|false||manifestation ofnull|Manifestation of|Modifier|false|false||manifestationnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Hypoxemia|Finding|false|false||hypoxemia
null|Blood oxygen concentration below reference range (finding)|Finding|false|false||hypoxemianull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Hypercapnia|Finding|false|false||hypercarbianull|Cardiac Arrest|Disorder|false|false||arrestnull|Encounter due to problems related to other legal circumstances - arrest|Finding|false|false||arrestnull|Law enforcement arrest|Event|false|false||arrestnull|Arrested progression|Time|false|false||arrestnull|Cognitive|Finding|false|false||cognitivenull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Unable|Finding|false|false||unablenull|Ventilator - respiratory equipment|Device|false|false||ventilator
null|null|Device|false|false||ventilatornull|Location Equipment - Ventilator|Modifier|false|false||ventilatornull|Capacity|LabModifier|false|false||capacitynull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Intubation (procedure)|Procedure|false|false||intubationnull|Mechanical ventilation finding|Finding|false|false||mechanical ventilationnull|Mechanical ventilation|Procedure|false|false||mechanical ventilationnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Ventilation, function (observable entity)|Finding|false|false||ventilation
null|Respiration|Finding|false|false||ventilationnull|Assisted breathing|Procedure|false|false||ventilationnull|Environmental air flow|Phenomenon|false|false||ventilationnull|Mechanical ventilation finding|Finding|false|false||mechanical ventilationnull|Mechanical ventilation|Procedure|false|false||mechanical ventilationnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Ventilation, function (observable entity)|Finding|false|false||ventilation
null|Respiration|Finding|false|false||ventilationnull|Assisted breathing|Procedure|false|false||ventilationnull|Environmental air flow|Phenomenon|false|false||ventilationnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Ventilation, function (observable entity)|Finding|false|false||ventilation
null|Respiration|Finding|false|false||ventilationnull|Assisted breathing|Procedure|false|false||ventilationnull|Environmental air flow|Phenomenon|false|false||ventilationnull|Extensive|Modifier|false|false||extensivenull|Discussion (procedure)|Procedure|false|false||discussionsnull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|daunorubicin|Drug|false|false||DNR
null|daunorubicin|Drug|false|false||DNRnull|Do-Not-Resuscitate Orders|Finding|false|false||DNR
null|Do not resuscitate status|Finding|false|false||DNRnull|null|Attribute|false|false||DNRnull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|spending|LabModifier|false|false||spendnull|Quality|Modifier|false|false||qualitynull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Morning|Time|false|false||morningnull|null|Finding|false|false||Autopsynull|Autopsy - Consent type|Procedure|false|false||Autopsy
null|Autopsy|Procedure|false|false||Autopsynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Ruta graveolens preparation|Drug|false|false||RUE
null|Ruta graveolens preparation|Drug|false|false||RUEnull|Ruta graveolens|Entity|false|false||RUE
null|Ruta|Entity|false|false||RUEnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Atrial Fibrillation|Disorder|false|false||atrial fibrillationnull|null|Attribute|false|false||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|argatroban|Drug|false|false||argatroban
null|argatroban|Drug|false|false||argatrobannull|Concern|Finding|false|false||concernnull|Heparin-induced thrombocytopenia|Disorder|false|false||HITnull|Hit - database search return|Finding|false|false||HITnull|Hittite Language|Entity|false|false||HITnull|Struck by|Modifier|false|false||HITnull|Platelet Factor 4, human|Drug|false|false||PF4
null|Platelet Factor 4, human|Drug|false|false||PF4
null|Platelet Factor 4|Drug|false|false||PF4
null|Platelet Factor 4|Drug|false|false||PF4null|PF4 gene|Finding|false|false||PF4null|antibodies (medication)|Drug|false|false||antibodies
null|antibodies (medication)|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodiesnull|IPSS-R Risk Category Very Low|Finding|false|false||very low
null|Very low (qualifier value)|Finding|false|false||very lownull|Very|Modifier|false|false||verynull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Unlikely|Finding|false|false||unlikelynull|Unlikely Related to Intervention|Modifier|false|false||unlikelynull|Acute sinusitis|Disorder|false|false||acute sinusitisnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Sinusitis|Disorder|false|false||sinusitisnull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Calcitrate|Drug|false|false||Calcitrate
null|Calcitrate|Drug|false|false||Calcitratenull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|calcium citrate|Drug|false|false||calcium citrate
null|calcium citrate|Drug|false|false||calcium citratenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|citrate|Drug|false|false||citrate
null|citrate|Drug|false|false||citrate
null|Citrates|Drug|false|false||citratenull|Citrate measurement|Procedure|false|false||citratenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|Theophylline SR|Drug|false|false||Theophylline SR
null|Theophylline SR|Drug|false|false||Theophylline SRnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Term (lexical)|Finding|false|false||term
null|Term Birth|Finding|false|false||termnull|Term (temporal)|Time|false|false||termnull|Use of steroids|Finding|false|false||steroid usenull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONE
null|prednisone|Drug|false|false||PredniSONEnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||Insomnianull|Sleeplessness|Finding|false|false||Insomnianull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Vertigo as late effect of cerebrovascular disease|Disorder|false|false||vertigonull|Vertigo|Finding|false|false||vertigonull|Vertigo <Vertiginidae>|Entity|false|false||vertigonull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|Once a day, at bedtime|Time|false|false||QHSnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|Wheezing|Finding|false|false||Wheezingnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|guaifenesin|Drug|false|false||Guaifenesin
null|guaifenesin|Drug|false|false||Guaifenesinnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal dosage form|Drug|false|false||NASALnull|Nasal Route of Administration|Finding|false|false||NASAL
null|Nasal (intended site)|Finding|false|false||NASALnull|null|Anatomy|false|false||NASALnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Hypersensitivity|Finding|false|false||allergiesnull|null|Attribute|false|false||allergiesnull|ferrous sulfate|Drug|false|false||Ferrous Sulfate
null|ferrous sulfate|Drug|false|false||Ferrous Sulfatenull|Ferrous|Drug|false|false||Ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Daily|Time|false|false||DAILYnull|dorzolamide|Drug|false|false||Dorzolamide
null|dorzolamide|Drug|false|false||Dorzolamidenull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Sodium Chloride Nasal Product|Drug|false|false||Sodium Chloride Nasalnull|sodium chloride|Drug|false|false||Sodium Chloridenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Four times daily|Time|false|false||QIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nasal discomfort|Finding|false|false||nasal discomfortnull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Discomfort|Finding|false|false||discomfortnull|morphine sulfate|Drug|false|false||Morphine Sulfate
null|morphine sulfate|Drug|false|false||Morphine Sulfatenull|morphine|Drug|false|false||Morphine
null|morphine|Drug|false|false||Morphinenull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Oral Solution|Drug|false|false||Oral Solutionnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|Kilogram per Cubic Meter|LabModifier|false|false||mg/mLnull|per milliliter|LabModifier|false|false||/mLnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Budesonide Nasal (Brand Name)|Drug|false|false||Budesonide Nasal
null|Budesonide Nasal Product|Drug|false|false||Budesonide Nasalnull|budesonide|Drug|false|false||Budesonide
null|budesonide|Drug|false|false||Budesonidenull|Nasal Inhaler|Device|false|false||Nasal Inhaler
null|Inhalers, Nasal|Device|false|false||Nasal Inhalernull|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal brand of oxymetazoline|Drug|false|false||Nasal
null|Nasal dosage form|Drug|false|false||Nasalnull|Nasal Route of Administration|Finding|false|false||Nasal
null|Nasal (intended site)|Finding|false|false||Nasalnull|null|Anatomy|false|false||Nasalnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Certificate Status - Expired|Finding|false|false||Expired
null|Referral status - Expired|Finding|false|false||Expired
null|Cessation of life|Finding|false|false||Expired
null|Expiration, Respiratory|Finding|false|false||Expired
null|Expiration|Finding|false|false||Expirednull|Specimen Reject Reason - Expired|Modifier|false|false||Expirednull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Pisum sativum (pea) extract|Drug|false|false||PEA
null|null|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|pea allergenic extract|Drug|false|false||PEA
null|Pisum sativum (pea) extract|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|phosphoethanolamine|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|PEA Preparation|Drug|false|false||PEA
null|palmidrol|Drug|false|false||PEAnull|Electromechanical dissociation|Disorder|false|false||PEAnull|area PEa of Pandya|Anatomy|false|false||PEAnull|Pisum sativum|Entity|false|false||PEAnull|Cardiac Arrest|Disorder|false|false||Arrestnull|Encounter due to problems related to other legal circumstances - arrest|Finding|false|false||Arrestnull|Law enforcement arrest|Event|false|false||Arrestnull|Arrested progression|Time|false|false||Arrestnull|Respiratory Failure|Disorder|false|false||Respiratory Failurenull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Sinusitis|Disorder|false|false||Sinusitisnull|Ruta graveolens preparation|Drug|false|false||RUE
null|Ruta graveolens preparation|Drug|false|false||RUEnull|Ruta graveolens|Entity|false|false||RUE
null|Ruta|Entity|false|false||RUEnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis|Procedure|false|false||DIAGNOSESnull|Atrial Fibrillation|Disorder|false|false||Atrial fibrillationnull|null|Attribute|false|false||Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Atrial fibrillationnull|Heart Atrium|Anatomy|false|false||Atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions