CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Plastics|Drug|false|false||PLASTICnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Paxil|Drug|false|false||Paxil
null|Paxil|Drug|false|false||Paxilnull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Craniotomy|Procedure|false|false||craniotomynull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Scalp flap|Anatomy|false|false||scalp flapnull|Scalp structure|Anatomy|false|false||scalpnull|ALOX5AP gene|Finding|false|false||flapnull|Surgical Flaps|Anatomy|false|false||flapnull|Split thickness graft of skin (substance)|Drug|false|false||split thickness skin graftnull|Split thickness skin graft (procedure)|Procedure|false|false||split thickness skin graftnull|Splitting|Finding|false|false||splitnull|Thickness of skin|Finding|false|false||thickness skinnull|Thick|Modifier|false|false||thicknessnull|Skin graft material|Drug|false|false||skin graftnull|skin graft (physical finding)|Finding|false|false||skin graftnull|Skin Transplantation|Procedure|false|false||skin graftnull|Transplanted skin|Anatomy|false|false||skin graftnull|Skin and subcutaneous tissue disorders|Disorder|false|false||skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||VACnull|VAC Regimen (Vincristine-Dactinomycin-Cyclophosphamide)|Procedure|false|false||VAC
null|cyclophosphamide/doxorubicin/vinblastine protocol|Procedure|false|false||VAC
null|cyclophosphamide/dactinomycin/vinblastine protocol|Procedure|false|false||VAC
null|VAC protocol|Procedure|false|false||VACnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Numerous|LabModifier|false|false||multiplenull|null|Time|false|false||priornull|Operative Surgical Procedures|Procedure|false|false||surgeriesnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Chemotherapy Regimen|Procedure|false|false||chemo
null|Chemotherapy|Procedure|false|false||chemonull|Radiation Ionizing Radiotherapy|Procedure|false|false||radiation
null|Radiotherapy Research|Procedure|false|false||radiation
null|Radiation therapy (procedure)|Procedure|false|false||radiationnull|Electromagnetic Radiation|Phenomenon|false|false||radiation
null|Radiation|Phenomenon|false|false||radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Pruritus|Finding|false|false||pruritusnull|sensory perception of itch|Modifier|false|false||pruritusnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|husband|Subject|false|false||husbandnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Metals|Drug|false|false||metalnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Metals|Drug|false|false||metalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Bone flap|Anatomy|true|false||bone flapnull|Specimen Type - Bone|Finding|true|false||bone
null|null|Finding|true|false||bonenull|Skeletal bone|Anatomy|true|false||bone
null|XXX bone|Anatomy|true|false||bonenull|ALOX5AP gene|Finding|true|false||flapnull|Surgical Flaps|Anatomy|true|false||flapnull|Rotational|Modifier|false|false||rotationalnull|ALOX5AP gene|Finding|false|false||flapnull|Surgical Flaps|Anatomy|false|false||flapnull|Skin graft material|Drug|false|false||skin graftnull|skin graft (physical finding)|Finding|false|false||skin graftnull|Skin Transplantation|Procedure|false|false||skin graftnull|Transplanted skin|Anatomy|false|false||skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|coverage - HL7PublishingDomain|Finding|false|false||coverage
null|null|Finding|false|false||coverage
null|coverage - financial contract|Finding|false|false||coveragenull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||Craniotomynull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Craniotomy|Procedure|false|false||craniotomynull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Accutane|Drug|false|false||Accutane
null|Accutane|Drug|false|false||Accutanenull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Disease|Disorder|false|false||diseasenull|Tubal Ligation|Procedure|false|false||tubal ligationnull|Ligation|Procedure|false|false||ligationnull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Acute bronchitis|Disorder|false|false||bronchitis
null|Bronchitis|Disorder|false|false||bronchitisnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Seizures|Finding|false|false||seizuresnull|Apyrexial|Finding|false|false||Afebrilenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Scalp structure|Anatomy|false|false||scalpnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Cleaning (activity)|Event|false|false||cleannull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Body Substance Discharge|Finding|true|false||drainage
null|Body Fluid Discharge|Finding|true|false||drainagenull|Drainage procedure|Procedure|true|false||drainagenull|Hemorrhage|Finding|true|false||bleedingnull|Admission activity|Procedure|true|false||admission
null|Hospital admission|Procedure|true|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Plastic surgery service|Entity|false|false||plastic surgery servicenull|Plastic Surgical Procedures|Procedure|false|false||plastic surgerynull|Plastic Surgery Specialty|Title|false|false||plastic surgerynull|Plastics|Drug|false|false||plasticnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|ALOX5AP gene|Finding|false|false||flapnull|Surgical Flaps|Anatomy|false|false||flapnull|Skin graft material|Drug|false|false||skin graftnull|skin graft (physical finding)|Finding|false|false||skin graftnull|Skin Transplantation|Procedure|false|false||skin graftnull|Transplanted skin|Anatomy|false|false||skin graftnull|Skin and subcutaneous tissue disorders|Disorder|false|false||skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Scalp defect|Disorder|false|false||scalp defectnull|Scalp structure|Anatomy|false|false||scalpnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Pain Relief brand of acetaminophen|Drug|false|false||pain relief
null|Pain Relief brand of acetaminophen|Drug|false|false||pain reliefnull|Pain relief|Procedure|false|false||pain reliefnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Cardiovascular system|Anatomy|false|false||cardiovascular
null|Cardiovascular|Anatomy|false|false||cardiovascularnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Oral intake|Finding|false|false||oral intakenull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Appropriate|Modifier|false|false||appropriatenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Intestines|Anatomy|false|false||bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Defecation|Finding|false|false||bowel movementnull|Intestines|Anatomy|false|false||bowelnull|Movement|Finding|false|false||movementnull|Measuring intake and output|Procedure|false|false||Intake and outputnull|Intake|Finding|false|false||Intakenull|Measurement of fluid intake|Procedure|false|false||Intake
null|Intake (treatment)|Procedure|false|false||Intakenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|On IV|Finding|false|false||on IVnull|cefazolin|Drug|false|false||cefazolin
null|cefazolin|Drug|false|false||cefazolinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|cefadroxil|Drug|false|false||cefadroxil
null|cefadroxil|Drug|false|false||cefadroxilnull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Prophylactic treatment|Procedure|false|false||Prophylaxisnull|prevention & control|Modifier|false|false||Prophylaxisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|subcutaneous heparin|Drug|false|false||subcutaneous heparin
null|subcutaneous heparin|Drug|false|false||subcutaneous heparinnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Ambulate|Finding|false|false||ambulatenull|Early|Time|false|false||earlynull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|null|Finding|true|false||regular dietnull|Regular|Modifier|true|false||regularnull|Diet (animal life circumstance)|Drug|true|false||diet
null|Diet|Drug|true|false||dietnull|diet - supply|Finding|true|false||dietnull|Diet therapy|Procedure|true|false||dietnull|Urination|Finding|true|false||voiding
null|Voids|Finding|true|false||voidingnull|Helping Behavior|Finding|true|false||assistancenull|Assisted (qualifier value)|Modifier|true|false||assistancenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Scalp structure|Anatomy|false|false||scalpnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Cleaning (activity)|Event|false|false||cleannull|Pink color|Modifier|false|false||pinknull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Entity|Entity|false|false||thingnull|Donor graft|Drug|false|false||graft donornull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|Donor site|Anatomy|false|false||donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Original|Modifier|false|false||originalnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|Ability to dress|Finding|false|false||dressing
null|null|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Pentasa|Drug|false|false||Pentasa
null|Pentasa|Drug|false|false||Pentasanull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|zolpidem|Drug|false|false||zolpidem
null|zolpidem|Drug|false|false||zolpidemnull|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl er
null|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl ernull|venlafaxine hydrochloride|Drug|false|false||venlafaxine hcl
null|venlafaxine hydrochloride|Drug|false|false||venlafaxine hclnull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|Flinders medical centre-7 marker|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hclnull|Hairy Cell Leukemia|Disorder|false|false||hclnull|promethazine|Drug|false|false||promethazine
null|promethazine|Drug|false|false||promethazinenull|Keflex|Drug|false|false||keflex
null|Keflex|Drug|false|false||keflexnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|dicyclomine|Drug|false|false||dicyclomine
null|dicyclomine|Drug|false|false||dicyclominenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Every eight hours|Time|false|false||Q8Hnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false||Disknull|Disc - Body Part|Anatomy|false|false||Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|mesalamine|Drug|false|false||mesalamine
null|mesalamine|Drug|false|false||mesalaminenull|Extended Release Oral Capsule|Drug|false|false||Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Extended Release Oral Capsule|Drug|false|false||Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Four times daily|Time|false|false||QIDnull|4 times|Finding|false|false||4 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false||Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|propylthiouracil|Drug|false|false||propylthiouracil
null|propylthiouracil|Drug|false|false||propylthiouracilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every eight hours|Time|false|false||Q8Hnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|bacitracin zinc|Drug|false|false||bacitracin zinc
null|bacitracin zinc|Drug|false|false||bacitracin zincnull|bacitracin|Drug|false|false||bacitracin
null|bacitracin|Drug|false|false||bacitracinnull|Zinc Supplements|Drug|false|false||zinc
null|Zinc Drug Class|Drug|false|false||zinc
null|Dietary Zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zincnull|Zinc measurement|Procedure|false|false||zincnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Ointments|Drug|false|false||Ointmentnull|APPL1 gene|Finding|false|false||Applnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|refill|Finding|false|false||Refillsnull|cefadroxil|Drug|false|false||cefadroxil
null|cefadroxil|Drug|false|false||cefadroxilnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|MAX protein, human|Drug|false|false||Max
null|MAX protein, human|Drug|false|false||Maxnull|Max (cigarettes)|Finding|false|false||Max
null|Oncogene MAX|Finding|false|false||Max
null|MAX gene|Finding|false|false||Maxnull|Maximum|LabModifier|false|false||Maxnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Craniotomy|Procedure|false|false||craniotomynull|Wound status|Finding|false|false||wound Statusnull|null|Attribute|false|false||wound Statusnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Hardware Removal|Procedure|false|false||hardware removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Splitting|Finding|false|false||splitnull|Thickness of skin|Finding|false|false||thickness skinnull|Thick|Modifier|false|false||thicknessnull|Skin graft material|Drug|false|false||skin graftnull|skin graft (physical finding)|Finding|false|false||skin graftnull|Skin Transplantation|Procedure|false|false||skin graftnull|Transplanted skin|Anatomy|false|false||skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|HL7 Version 2.5 - Application|Finding|false|false||application
null|Application Document|Finding|false|false||application
null|Computer Application|Finding|false|false||application
null|Regulatory Application|Finding|false|false||application
null|Apply|Finding|false|false||applicationnull|Application procedure|Procedure|false|false||applicationnull|Application - unit of product usage|LabModifier|false|false||applicationnull|Scalp structure|Anatomy|false|false||scalpnull|Donor site|Anatomy|false|false||donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Always - AcknowledgementCondition|Finding|false|false||always
null|All of the Time|Finding|false|false||alwaysnull|Always (frequency)|Time|false|false||alwaysnull|Apply (administration method)|Finding|false|false||apply
null|Apply (instruction)|Finding|false|false||apply
null|null|Finding|false|false||apply
null|Apply|Finding|false|false||applynull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Suction drainage|Procedure|false|false||suctionnull|Location Equipment - Suction|Modifier|false|false||suctionnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Suction drainage|Procedure|true|false||suctionnull|Location Equipment - Suction|Modifier|true|false||suctionnull|Skin graft material|Drug|false|false||skin graftnull|skin graft (physical finding)|Finding|false|false||skin graftnull|Skin Transplantation|Procedure|false|false||skin graftnull|Transplanted skin|Anatomy|false|false||skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Graft Dosage Form|Drug|false|false||graft
null|Graft material|Drug|false|false||graftnull|Graft - Specimen Source Codes|Finding|false|false||graftnull|Graft Procedures on the Head|Procedure|false|false||graft
null|Grafting procedure|Procedure|false|false||graftnull|Transplanted tissue|Anatomy|false|false||graftnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Scalp structure|Anatomy|false|false||scalpnull|Xeroform|Drug|false|false||Xeroform
null|Xeroform|Drug|false|false||Xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|null|Drug|false|false||bacitracin ointmentnull|bacitracin|Drug|false|false||bacitracin
null|bacitracin|Drug|false|false||bacitracinnull|Ointments|Drug|false|false||ointmentnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Warning - AcknowledgementDetailType|Finding|false|false||WARNING
null|Cautionary Warning|Finding|false|false||WARNING
null|System Alert|Finding|false|false||WARNING
null|Warning - Error severity|Finding|false|false||WARNING
null|Warning - EquipmentAlertLevel|Finding|false|false||WARNINGnull|Warning - Alert level|Modifier|false|false||WARNINGnull|Xeroform|Drug|true|false||xeroform
null|Xeroform|Drug|true|false||xeroformnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Skin graft material|Drug|true|false||skin graftnull|skin graft (physical finding)|Finding|true|false||skin graftnull|Skin Transplantation|Procedure|true|false||skin graftnull|Transplanted skin|Anatomy|true|false||skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|true|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|true|false||skinnull|Skin Specimen Source Code|Finding|true|false||skin
null|Skin Specimen|Finding|true|false||skinnull|Skin, Human|Anatomy|true|false||skin
null|Skin|Anatomy|true|false||skinnull|Graft Dosage Form|Drug|true|false||graft
null|Graft material|Drug|true|false||graftnull|Graft - Specimen Source Codes|Finding|true|false||graftnull|Graft Procedures on the Head|Procedure|true|false||graft
null|Grafting procedure|Procedure|true|false||graftnull|Transplanted tissue|Anatomy|true|false||graftnull|null|Finding|true|false||sitenull|Anatomic Site|Anatomy|true|false||sitenull|Study Site|Modifier|true|false||site
null|Site|Modifier|true|false||sitenull|Free of (attribute)|Finding|true|false||free ofnull|Free of (attribute)|Finding|true|false||freenull|Empty (qualifier)|Modifier|true|false||freenull|Pressure (finding)|Finding|true|false||pressure
null|null|Finding|true|false||pressure
null|Baresthesia|Finding|true|false||pressurenull|null|Phenomenon|true|false||pressurenull|Pressure (property)|LabModifier|true|false||pressurenull|Temperature extreme|Phenomenon|true|false||extreme temperaturesnull|Extreme Response|Finding|true|false||extremenull|Extreme|Modifier|true|false||extremenull|Temperature|LabModifier|true|false||temperaturesnull|null|Finding|true|false||covernull|Cover (physical object)|Device|true|false||cover
null|Cover Device|Device|true|false||covernull|Loose|Modifier|true|false||loosenull|Graft Dosage Form|Drug|true|false||graft
null|Graft material|Drug|true|false||graftnull|Graft - Specimen Source Codes|Finding|true|false||graftnull|Graft Procedures on the Head|Procedure|true|false||graft
null|Grafting procedure|Procedure|true|false||graftnull|Transplanted tissue|Anatomy|true|false||graftnull|null|Finding|true|false||sitenull|Anatomic Site|Anatomy|true|false||sitenull|Study Site|Modifier|true|false||site
null|Site|Modifier|true|false||sitenull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Water running|Procedure|true|false||water runnull|Running water|Phenomenon|true|false||water runnull|Water Specimen|Drug|true|false||water
null|water|Drug|true|false||water
null|water|Drug|true|false||waternull|Water - Specimen Source Codes|Finding|true|false||waternull|Hydrotherapy|Procedure|true|false||waternull|Does run (finding)|Finding|true|false||run
null|Running (physical activity)|Finding|true|false||run
null|Go Jogging or Running Question|Finding|true|false||run
null|Run action|Finding|true|false||runnull|Rundi language|Entity|true|false||runnull|Problems with head|Disorder|true|false||headnull|Procedure on head|Procedure|true|false||headnull|Structure of head of caudate nucleus|Anatomy|true|false||head
null|Head|Anatomy|true|false||headnull|Head Device|Device|true|false||headnull|Scalp structure|Anatomy|false|false||scalpnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Donor site|Anatomy|false|false||donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Old|Time|false|false||oldnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Own|Finding|false|false||ownnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Plastics|Drug|false|false||Plasticnull|Free of (attribute)|Finding|false|false||free ofnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Shower (physical object)|Device|false|false||showernull|Plastics|Drug|false|false||plasticnull|Leave from Employment|Finding|false|false||leavenull|null|Event|false|false||leavenull|Donor site|Anatomy|false|false||donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Decompression Sickness|Disorder|true|false||bendnull|Does bend|Finding|true|false||bendnull|Heavy (weight) (qualifier value)|Modifier|true|false||heavy
null|Heavy (amount)|Modifier|true|false||heavynull|Lifting|Event|true|false||liftingnull|Strenuous Exercise|Finding|true|false||strenuous activitynull|Strenuous|Modifier|true|false||strenuousnull|Activity (animal life circumstance)|Finding|true|false||activity
null|Physical activity|Finding|true|false||activitynull|Activities|Event|true|false||activitynull|null|Modifier|true|false||activitynull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Regular|Modifier|false|false||regularnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenol
null|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenolnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Mild pain|Finding|false|false||mild pain
null|Neck Pain Score 2|Finding|false|false||mild painnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Packaging Materials|Device|false|false||packaging
null|Drug Packaging|Device|false|false||packagingnull|Packaging|Phenomenon|false|false||packagingnull|Packing (action)|Event|false|false||packagingnull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|Vicodin|Drug|false|false||Vicodin
null|Vicodin|Drug|false|false||Vicodinnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Active ingredient|Drug|true|false||active ingredientnull|Has active ingredient|Modifier|true|false||active ingredientnull|Ingredient|Drug|true|false||ingredientnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Additional|Finding|true|false||additionalnull|Tylenol|Drug|true|false||Tylenol
null|Tylenol|Drug|true|false||Tylenolnull|prescription document|Finding|true|false||prescriptionnull|Prescription (procedure)|Procedure|true|false||prescriptionnull|Prescription (attribute)|Attribute|true|false||prescriptionnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Tylenol|Drug|true|false||tylenol
null|Tylenol|Drug|true|false||tylenolnull|Antibiotics|Drug|false|false||antibioticnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|2 times per day|Finding|false|false||2 times per daynull|2 times|Finding|false|false||2 timesnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Different|Modifier|false|false||differentnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|heavy machinery|Device|true|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|true|false||heavy
null|Heavy (amount)|Modifier|true|false||heavynull|Contact with machinery|Disorder|true|false||machinerynull|Industrial machine|Device|true|false||machinerynull|Narcotics|Drug|true|false||narcotic
null|Narcotics|Drug|true|false||narcoticnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Have Constipation|Finding|false|false||have constipationnull|Constipation|Finding|false|false||constipationnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Etc.|Finding|false|false||etcnull|Drinking (function)|Finding|false|false||drinking
null|Alcohol consumption|Finding|false|false||drinkingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Stool Softener|Drug|false|false||stool softenersnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Food|Drug|false|false||foodsnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Fiber brand of calcium polycarbophil|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false||fibernull|Tissue fiber|Anatomy|false|false||fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Pharmaceutical Preparations|Drug|true|false||medicinesnull|Motrin|Drug|true|false||Motrin
null|Motrin|Drug|true|false||Motrinnull|aspirin|Drug|true|false||Aspirin
null|aspirin|Drug|true|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Etc.|Finding|false|false||etcnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Following|Time|true|false||following
null|Status post|Time|true|false||followingnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Fever with chills|Finding|false|false||fever with chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Physiologic warmth|Finding|false|false||warmth
null|Social warmth|Finding|false|false||warmthnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Unusual|Modifier|false|false||unusualnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Large amount|LabModifier|false|false||large amountnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Hemorrhage|Finding|false|false||bleedingnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than|LabModifier|true|false||greater thannull|Greater|LabModifier|false|false||greaternull|Severe Extremity Pain|Finding|true|false||Severe pain
null|Severe pain|Finding|true|false||Severe pain
null|Neck Pain Score 6|Finding|true|false||Severe painnull|Severe - Severity of Illness Code|Finding|true|false||Severe
null|Intensity and Distress 5|Finding|true|false||Severe
null|Severe - Triage Code|Finding|true|false||Severe
null|Severe (severity modifier)|Finding|true|false||Severe
null|Allergy Severity - Severe|Finding|true|false||Severenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Vomiting|Finding|true|false||vomitingnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Else|Finding|false|false||elsenull|Equipment Alert Level - Serious|Finding|true|false||serious
null|Device Alert Level - Serious|Finding|true|false||serious
null|Alert level - Serious|Finding|true|false||seriousnull|Serious|Modifier|true|false||seriousnull|Changing|Finding|true|false||change innull|Changed status|LabModifier|true|false||change innull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Concern|Finding|true|false||concernnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions