 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
F|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
SURGERY|159,166
<EOL>|166,167
<EOL>|168,169
Patient|181,188
recorded|189,197
as|198,200
having|201,207
No|208,210
Known|211,216
Allergies|217,226
to|227,229
Drugs|230,235
<EOL>|235,236
<EOL>|237,238
Attending|238,247
:|247,248
_|249,250
_|250,251
_|251,252
.|252,253
<EOL>|253,254
<EOL>|255,256
diverticulitis|273,287
<EOL>|287,288
<EOL>|289,290
Major|290,295
Surgical|296,304
or|305,307
Invasive|308,316
Procedure|317,326
:|326,327
<EOL>|327,328
s|328,329
/|329,330
p|330,331
laparoscopic|332,344
sigmoid|345,352
colectomy|353,362
<EOL>|363,364
<EOL>|364,365
<EOL>|366,367
Mrs.|395,399
_|400,401
_|401,402
_|402,403
is|404,406
a|407,408
_|409,410
_|410,411
_|411,412
F|413,414
with|415,419
history|420,427
of|428,430
recurrent|431,440
diverticulitis|441,455
,|455,456
<EOL>|457,458
originally|458,468
<EOL>|468,469
diagnosed|469,478
_|479,480
_|480,481
_|481,482
_|483,484
_|484,485
_|485,486
.|486,487
Pt|488,490
reports|491,498
a|499,500
one|501,504
month|505,510
history|511,518
of|519,521
<EOL>|522,523
LLQ|523,526
<EOL>|526,527
pain|527,531
varying|532,539
_|540,541
_|541,542
_|542,543
intensity|544,553
.|553,554
Pt|555,557
was|558,561
prescribed|562,572
a|573,574
10|575,577
day|578,581
course|582,588
of|589,591
<EOL>|591,592
Cipro|592,597
/|597,598
Flagyl|598,604
PO|605,607
which|608,613
she|614,617
completed|618,627
on|628,630
_|631,632
_|632,633
_|633,634
.|634,635
Pt|636,638
was|639,642
doing|643,648
<EOL>|649,650
well|650,654
<EOL>|654,655
until|655,660
abdominal|661,670
pain|671,675
returned|676,684
_|685,686
_|686,687
_|687,688
,|688,689
one|690,693
week|694,698
after|699,704
finishing|705,714
<EOL>|714,715
antibiotic|715,725
course|726,732
.|732,733
Pt|734,736
reports|737,744
no|745,747
nausea|748,754
or|755,757
vomiting|758,766
,|766,767
pt|768,770
has|771,774
been|775,779
<EOL>|779,780
able|780,784
to|785,787
maintain|788,796
hydration|797,806
with|807,811
regular|812,819
PO|820,822
intake|823,829
although|830,838
<EOL>|838,839
appetite|839,847
has|848,851
been|852,856
somewhat|857,865
decreased|866,875
.|875,876
Pt|877,879
has|880,883
been|884,888
having|889,895
<EOL>|896,897
regular|897,904
,|904,905
<EOL>|905,906
non-bloody|906,916
bowel|917,922
movements|923,932
,|932,933
pt|934,936
reports|937,944
several|945,952
small|953,958
,|958,959
soft|960,964
-|964,965
brown|965,970
<EOL>|970,971
bowel|971,976
movements|977,986
today|987,992
.|992,993
No|994,996
diarrhea|997,1005
.|1005,1006
Pt|1007,1009
presents|1010,1018
to|1019,1021
_|1022,1023
_|1023,1024
_|1024,1025
today|1026,1031
<EOL>|1032,1033
as|1033,1035
<EOL>|1035,1036
a|1036,1037
direct|1038,1044
admission|1045,1054
for|1055,1058
refractory|1059,1069
LLQ|1070,1073
pain|1074,1078
.|1078,1079
<EOL>|1079,1080
<EOL>|1080,1081
<EOL>|1082,1083
diverticulitis|1105,1119
<EOL>|1119,1120
Migraines|1120,1129
<EOL>|1129,1130
Left|1130,1134
finger|1135,1141
cellulitis|1142,1152
<EOL>|1152,1153
<EOL>|1154,1155
:|1169,1170
<EOL>|1170,1171
_|1171,1172
_|1172,1173
_|1173,1174
<EOL>|1174,1175
:|1189,1190
<EOL>|1190,1191
father|1191,1197
with|1198,1202
h|1203,1204
/|1204,1205
o|1205,1206
colitis|1207,1214
<EOL>|1214,1215
<EOL>|1216,1217
Crimson|1232,1239
Admission|1240,1249
<EOL>|1249,1250
Temp|1250,1254
98.6|1255,1259
,|1259,1260
HR|1261,1263
70|1264,1266
,|1266,1267
BP|1268,1270
110|1271,1274
/|1274,1275
70|1275,1277
,|1277,1278
RR|1279,1281
18|1282,1284
,|1284,1285
96|1286,1288
%|1288,1289
RA|1290,1292
<EOL>|1292,1293
Gen|1293,1296
:|1296,1297
well|1298,1302
,|1302,1303
NAD|1304,1307
,|1307,1308
A|1309,1310
&|1310,1311
O|1311,1312
<EOL>|1312,1313
CV|1313,1315
:|1315,1316
RRR|1317,1320
,|1320,1321
No|1322,1324
R|1325,1326
/|1326,1327
G|1327,1328
/|1328,1329
M|1329,1330
<EOL>|1330,1331
RESP|1331,1335
:|1335,1336
CTAB|1337,1341
<EOL>|1341,1342
ABD|1342,1345
:|1345,1346
Focal|1347,1352
tenderness|1353,1363
LLQ|1364,1367
inferolateral|1368,1381
to|1382,1384
umbilicus|1385,1394
,|1394,1395
otherwise|1396,1405
<EOL>|1405,1406
NT|1406,1408
,|1408,1409
ND|1410,1412
,|1412,1413
no|1414,1416
guarding|1417,1425
or|1426,1428
rebound|1429,1436
<EOL>|1436,1437
EXT|1437,1440
:|1440,1441
No|1442,1444
edema|1445,1450
<EOL>|1450,1451
<EOL>|1451,1452
<EOL>|1453,1454
Pertinent|1454,1463
Results|1464,1471
:|1471,1472
<EOL>|1472,1473
RADIOLOGY|1473,1482
Final|1484,1489
Report|1490,1496
<EOL>|1496,1497
CT|1497,1499
PELVIS|1500,1506
W|1507,1508
/|1508,1509
CONTRAST|1509,1517
_|1519,1520
_|1520,1521
_|1521,1522
2|1523,1524
:|1524,1525
58|1525,1527
AM|1528,1530
<EOL>|1530,1531
UNDERLYING|1531,1541
MEDICAL|1542,1549
CONDITION|1550,1559
:|1559,1560
<EOL>|1560,1561
_|1561,1562
_|1562,1563
_|1563,1564
year|1565,1569
old|1570,1573
woman|1574,1579
with|1580,1584
diverticulitis|1585,1599
,|1599,1600
increasing|1601,1611
RLQ|1612,1615
pain|1616,1620
<EOL>|1621,1622
IMPRESSION|1622,1632
:|1632,1633
Moderate|1634,1642
uncomplicated|1643,1656
diverticulitis|1657,1671
at|1672,1674
the|1675,1678
<EOL>|1679,1680
junction|1680,1688
of|1689,1691
the|1692,1695
descending|1696,1706
colon|1707,1712
and|1713,1716
sigmoid|1717,1724
colon|1725,1730
.|1730,1731
Stable|1732,1738
<EOL>|1739,1740
mildly|1740,1746
enlarged|1747,1755
retroperitoneal|1756,1771
lymph|1772,1777
nodes|1778,1783
may|1784,1787
be|1788,1790
reactive|1791,1799
_|1800,1801
_|1801,1802
_|1802,1803
<EOL>|1804,1805
nature|1805,1811
.|1811,1812
If|1813,1815
surgery|1816,1823
has|1824,1827
not|1828,1831
been|1832,1836
contemplated|1837,1849
,|1849,1850
a|1851,1852
followup|1853,1861
is|1862,1864
<EOL>|1865,1866
recommended|1866,1877
_|1878,1879
_|1879,1880
_|1880,1881
six|1882,1885
weeks|1886,1891
,|1891,1892
to|1893,1895
assess|1896,1902
for|1903,1906
complete|1907,1915
resolution|1916,1926
of|1927,1929
<EOL>|1930,1931
these|1931,1936
findings|1937,1945
.|1945,1946
<EOL>|1946,1947
.|1947,1948
<EOL>|1948,1949
_|1949,1950
_|1950,1951
_|1951,1952
06|1953,1955
:|1955,1956
05AM|1956,1960
BLOOD|1961,1966
WBC|1967,1970
-|1970,1971
9.9|1971,1974
RBC|1975,1978
-|1978,1979
2|1979,1980
.|1980,1981
85|1981,1983
*|1983,1984
Hgb|1985,1988
-|1988,1989
8|1989,1990
.|1990,1991
9|1991,1992
*|1992,1993
Hct|1994,1997
-|1997,1998
25|1998,2000
.|2000,2001
9|2001,2002
*|2002,2003
<EOL>|2004,2005
MCV|2005,2008
-|2008,2009
91|2009,2011
MCH|2012,2015
-|2015,2016
31.3|2016,2020
MCHC|2021,2025
-|2025,2026
34.4|2026,2030
RDW|2031,2034
-|2034,2035
13.0|2035,2039
Plt|2040,2043
_|2044,2045
_|2045,2046
_|2046,2047
<EOL>|2047,2048
_|2048,2049
_|2049,2050
_|2050,2051
09|2052,2054
:|2054,2055
10AM|2055,2059
BLOOD|2060,2065
WBC|2066,2069
-|2069,2070
23|2070,2072
.|2072,2073
2|2073,2074
*|2074,2075
#|2075,2076
RBC|2077,2080
-|2080,2081
3|2081,2082
.|2082,2083
73|2083,2085
*|2085,2086
Hgb|2087,2090
-|2090,2091
11|2091,2093
.|2093,2094
6|2094,2095
*|2095,2096
Hct|2097,2100
-|2100,2101
33|2101,2103
.|2103,2104
5|2104,2105
*|2105,2106
<EOL>|2107,2108
MCV|2108,2111
-|2111,2112
90|2112,2114
MCH|2115,2118
-|2118,2119
31.0|2119,2123
MCHC|2124,2128
-|2128,2129
34.5|2129,2133
RDW|2134,2137
-|2137,2138
13.0|2138,2142
Plt|2143,2146
_|2147,2148
_|2148,2149
_|2149,2150
<EOL>|2150,2151
_|2151,2152
_|2152,2153
_|2153,2154
05|2155,2157
:|2157,2158
25AM|2158,2162
BLOOD|2163,2168
WBC|2169,2172
-|2172,2173
10.5|2173,2177
RBC|2178,2181
-|2181,2182
3|2182,2183
.|2183,2184
98|2184,2186
*|2186,2187
Hgb|2188,2191
-|2191,2192
12.7|2192,2196
Hct|2197,2200
-|2200,2201
34|2201,2203
.|2203,2204
4|2204,2205
*|2205,2206
<EOL>|2207,2208
MCV|2208,2211
-|2211,2212
87|2212,2214
MCH|2215,2218
-|2218,2219
32.0|2219,2223
MCHC|2224,2228
-|2228,2229
37|2229,2231
.|2231,2232
0|2232,2233
*|2233,2234
RDW|2235,2238
-|2238,2239
12.8|2239,2243
Plt|2244,2247
_|2248,2249
_|2249,2250
_|2250,2251
<EOL>|2251,2252
_|2252,2253
_|2253,2254
_|2254,2255
06|2256,2258
:|2258,2259
05AM|2259,2263
BLOOD|2264,2269
Plt|2270,2273
_|2274,2275
_|2275,2276
_|2276,2277
<EOL>|2277,2278
_|2278,2279
_|2279,2280
_|2280,2281
05|2282,2284
:|2284,2285
15AM|2285,2289
BLOOD|2290,2295
_|2296,2297
_|2297,2298
_|2298,2299
PTT|2300,2303
-|2303,2304
28.3|2304,2308
_|2309,2310
_|2310,2311
_|2311,2312
<EOL>|2312,2313
_|2313,2314
_|2314,2315
_|2315,2316
05|2317,2319
:|2319,2320
25AM|2320,2324
BLOOD|2325,2330
_|2331,2332
_|2332,2333
_|2333,2334
PTT|2335,2338
-|2338,2339
28.4|2339,2343
_|2344,2345
_|2345,2346
_|2346,2347
<EOL>|2347,2348
_|2348,2349
_|2349,2350
_|2350,2351
06|2352,2354
:|2354,2355
05AM|2355,2359
BLOOD|2360,2365
Glucose|2366,2373
-|2373,2374
109|2374,2377
*|2377,2378
UreaN|2379,2384
-|2384,2385
9|2385,2386
Creat|2387,2392
-|2392,2393
1|2393,2394
.|2394,2395
9|2395,2396
*|2396,2397
Na|2398,2400
-|2400,2401
138|2401,2404
<EOL>|2405,2406
K|2406,2407
-|2407,2408
3|2408,2409
.|2409,2410
2|2410,2411
*|2411,2412
Cl|2413,2415
-|2415,2416
100|2416,2419
HCO3|2420,2424
-|2424,2425
30|2425,2427
AnGap|2428,2433
-|2433,2434
11|2434,2436
<EOL>|2436,2437
_|2437,2438
_|2438,2439
_|2439,2440
05|2441,2443
:|2443,2444
25AM|2444,2448
BLOOD|2449,2454
Glucose|2455,2462
-|2462,2463
127|2463,2466
*|2466,2467
UreaN|2468,2473
-|2473,2474
5|2474,2475
*|2475,2476
Creat|2477,2482
-|2482,2483
0.6|2483,2486
Na|2487,2489
-|2489,2490
138|2490,2493
<EOL>|2494,2495
K|2495,2496
-|2496,2497
4.0|2497,2500
Cl|2501,2503
-|2503,2504
102|2504,2507
HCO3|2508,2512
-|2512,2513
27|2513,2515
AnGap|2516,2521
-|2521,2522
13|2522,2524
<EOL>|2524,2525
_|2525,2526
_|2526,2527
_|2527,2528
06|2529,2531
:|2531,2532
05AM|2532,2536
BLOOD|2537,2542
ALT|2543,2546
-|2546,2547
85|2547,2549
*|2549,2550
AST|2551,2554
-|2554,2555
49|2555,2557
*|2557,2558
LD|2559,2561
(|2561,2562
LDH|2562,2565
)|2565,2566
-|2566,2567
204|2567,2570
AlkPhos|2571,2578
-|2578,2579
208|2579,2582
*|2582,2583
<EOL>|2584,2585
TotBili|2585,2592
-|2592,2593
0.7|2593,2596
<EOL>|2596,2597
_|2597,2598
_|2598,2599
_|2599,2600
05|2601,2603
:|2603,2604
25AM|2604,2608
BLOOD|2609,2614
ALT|2615,2618
-|2618,2619
15|2619,2621
AST|2622,2625
-|2625,2626
14|2626,2628
LD|2629,2631
(|2631,2632
LDH|2632,2635
)|2635,2636
-|2636,2637
149|2637,2640
AlkPhos|2641,2648
-|2648,2649
47|2649,2651
<EOL>|2652,2653
Amylase|2653,2660
-|2660,2661
42|2661,2663
TotBili|2664,2671
-|2671,2672
1|2672,2673
.|2673,2674
7|2674,2675
*|2675,2676
<EOL>|2676,2677
_|2677,2678
_|2678,2679
_|2679,2680
06|2681,2683
:|2683,2684
05AM|2684,2688
BLOOD|2689,2694
Albumin|2695,2702
-|2702,2703
2|2703,2704
.|2704,2705
8|2705,2706
*|2706,2707
Calcium|2708,2715
-|2715,2716
8|2716,2717
.|2717,2718
2|2718,2719
*|2719,2720
Phos|2721,2725
-|2725,2726
2.8|2726,2729
Mg|2730,2732
-|2732,2733
2.4|2733,2736
<EOL>|2736,2737
_|2737,2738
_|2738,2739
_|2739,2740
05|2741,2743
:|2743,2744
25AM|2744,2748
BLOOD|2749,2754
Albumin|2755,2762
-|2762,2763
4.0|2763,2766
Calcium|2767,2774
-|2774,2775
8.9|2775,2778
Phos|2779,2783
-|2783,2784
3.5|2784,2787
Mg|2788,2790
-|2790,2791
2.0|2791,2794
<EOL>|2794,2795
_|2795,2796
_|2796,2797
_|2797,2798
05|2799,2801
:|2801,2802
15AM|2802,2806
BLOOD|2807,2812
Vanco|2813,2818
-|2818,2819
25.0|2819,2823
*|2823,2824
<EOL>|2824,2825
.|2825,2826
<EOL>|2826,2827
_|2827,2828
_|2828,2829
_|2829,2830
12|2831,2833
:|2833,2834
23|2834,2836
pm|2837,2839
SWAB|2840,2844
Site|2849,2853
:|2853,2854
ABDOMEN|2855,2862
<EOL>|2862,2863
Fluid|2869,2874
should|2875,2881
not|2882,2885
be|2886,2888
sent|2889,2893
_|2894,2895
_|2895,2896
_|2896,2897
swab|2898,2902
transport|2903,2912
media|2913,2918
.|2918,2919
Submit|2921,2927
<EOL>|2928,2929
fluids|2929,2935
_|2936,2937
_|2937,2938
_|2938,2939
a|2940,2941
<EOL>|2941,2942
capped|2948,2954
syringe|2955,2962
(|2963,2964
no|2964,2966
needle|2967,2973
)|2973,2974
,|2974,2975
red|2976,2979
top|2980,2983
tube|2984,2988
,|2988,2989
or|2990,2992
sterile|2993,3000
cup|3001,3004
.|3004,3005
<EOL>|3006,3007
GRAM|3010,3014
STAIN|3015,3020
(|3021,3022
Final|3022,3027
_|3028,3029
_|3029,3030
_|3030,3031
:|3031,3032
<EOL>|3033,3034
1|3040,3041
+|3041,3042
(|3046,3047
<|3047,3048
1|3048,3049
per|3050,3053
1000X|3054,3059
FIELD|3060,3065
)|3065,3066
:|3066,3067
POLYMORPHONUCLEAR|3070,3087
<EOL>|3088,3089
LEUKOCYTES|3089,3099
.|3099,3100
<EOL>|3101,3102
4|3108,3109
+|3109,3110
(|3113,3114
>|3114,3115
10|3115,3117
per|3118,3121
1000X|3122,3127
FIELD|3128,3133
)|3133,3134
:|3134,3135
GRAM|3138,3142
POSITIVE|3143,3151
COCCI|3152,3157
.|3157,3158
<EOL>|3159,3160
_|3194,3195
_|3195,3196
_|3196,3197
PAIRS|3198,3203
,|3203,3204
CHAINS|3205,3211
,|3211,3212
AND|3213,3216
CLUSTERS|3217,3225
<EOL>|3225,3226
FLUID|3229,3234
CULTURE|3235,3242
(|3243,3244
Final|3244,3249
_|3250,3251
_|3251,3252
_|3252,3253
:|3253,3254
<EOL>|3255,3256
STAPH|3262,3267
AUREUS|3268,3274
COAG|3275,3279
+|3280,3281
.|3281,3282
MODERATE|3286,3294
GROWTH|3295,3301
.|3301,3302
CLINDAMYCIN|3304,3315
PER|3316,3319
<EOL>|3320,3321
ID|3321,3323
.|3323,3324
.|3324,3325
<EOL>|3326,3327
This|3336,3340
isolate|3341,3348
is|3349,3351
presumed|3352,3360
to|3361,3363
be|3364,3366
resistant|3367,3376
to|3377,3379
clindamycin|3380,3391
<EOL>|3392,3393
based|3393,3398
on|3399,3401
<EOL>|3401,3402
the|3411,3414
detection|3415,3424
of|3425,3427
inducible|3428,3437
resistance|3438,3448
.|3449,3450
<EOL>|3450,3451
ANAEROBIC|3454,3463
CULTURE|3464,3471
(|3472,3473
Preliminary|3473,3484
)|3484,3485
:|3485,3486
NO|3490,3492
ANAEROBES|3493,3502
ISOLATED|3503,3511
.|3511,3512
<EOL>|3513,3514
ACID|3517,3521
FAST|3522,3526
SMEAR|3527,3532
(|3533,3534
Final|3534,3539
_|3540,3541
_|3541,3542
_|3542,3543
:|3543,3544
<EOL>|3545,3546
NO|3552,3554
ACID|3555,3559
FAST|3560,3564
BACILLI|3565,3572
SEEN|3573,3577
ON|3578,3580
DIRECT|3581,3587
SMEAR|3588,3593
.|3593,3594
<EOL>|3595,3596
ACID|3599,3603
FAST|3604,3608
CULTURE|3609,3616
(|3617,3618
Preliminary|3618,3629
)|3629,3630
:|3630,3631
<EOL>|3632,3633
A|3639,3640
swab|3641,3645
is|3646,3648
not|3649,3652
the|3653,3656
optimal|3657,3664
specimen|3665,3673
for|3674,3677
recovery|3678,3686
of|3687,3689
<EOL>|3690,3691
mycobacteria|3691,3703
or|3704,3706
<EOL>|3706,3707
filamentous|3713,3724
fungi|3725,3730
.|3730,3731
A|3733,3734
negative|3735,3743
result|3744,3750
should|3751,3757
be|3758,3760
<EOL>|3761,3762
interpreted|3762,3773
with|3774,3778
<EOL>|3778,3779
caution|3785,3792
.|3792,3793
Whenever|3795,3803
possible|3804,3812
tissue|3813,3819
biopsy|3820,3826
or|3827,3829
aspirated|3830,3839
<EOL>|3840,3841
fluid|3841,3846
should|3847,3853
<EOL>|3853,3854
be|3860,3862
submitted|3863,3872
.|3872,3873
<EOL>|3874,3875
FUNGAL|3878,3884
CULTURE|3885,3892
(|3893,3894
Preliminary|3894,3905
)|3905,3906
:|3906,3907
<EOL>|3908,3909
NO|3915,3917
FUNGUS|3918,3924
ISOLATED|3925,3933
.|3933,3934
<EOL>|3935,3936
A|3942,3943
swab|3944,3948
is|3949,3951
not|3952,3955
the|3956,3959
optimal|3960,3967
specimen|3968,3976
for|3977,3980
recovery|3981,3989
of|3990,3992
<EOL>|3993,3994
mycobacteria|3994,4006
or|4007,4009
<EOL>|4009,4010
filamentous|4016,4027
fungi|4028,4033
.|4033,4034
A|4036,4037
negative|4038,4046
result|4047,4053
should|4054,4060
be|4061,4063
<EOL>|4064,4065
interpreted|4065,4076
with|4077,4081
<EOL>|4081,4082
caution|4088,4095
.|4095,4096
Whenever|4098,4106
possible|4107,4115
tissue|4116,4122
biopsy|4123,4129
or|4130,4132
aspirated|4133,4142
<EOL>|4143,4144
fluid|4144,4149
should|4150,4156
<EOL>|4156,4157
be|4163,4165
submitted|4166,4175
.|4175,4176
<EOL>|4177,4178
.|4178,4179
<EOL>|4179,4180
Pathology|4180,4189
Examination|4190,4201
<EOL>|4202,4203
SPECIMEN|4203,4211
SUBMITTED|4212,4221
:|4221,4222
sigmoid|4223,4230
colon|4231,4236
.|4236,4237
<EOL>|4237,4238
Procedure|4238,4247
date|4248,4252
_|4257,4258
_|4258,4259
_|4259,4260
<EOL>|4261,4262
Sigmoid|4275,4282
colon|4283,4288
,|4288,4289
segmental|4290,4299
resection|4300,4309
:|4309,4310
<EOL>|4311,4312
Colonic|4312,4319
segment|4320,4327
with|4328,4332
organizing|4333,4343
pericolic|4344,4353
abscess|4354,4361
,|4361,4362
consistent|4363,4373
<EOL>|4374,4375
with|4375,4379
ruptured|4380,4388
diverticulum|4389,4401
.|4401,4402
<EOL>|4403,4404
Unremarkable|4404,4416
regional|4417,4425
lymph|4426,4431
nodes|4432,4437
.|4437,4438
<EOL>|4439,4440
No|4440,4442
intrinsic|4443,4452
mucosal|4453,4460
abnormalities|4461,4474
seen|4475,4479
.|4479,4480
<EOL>|4480,4481
Clinical|4481,4489
:|4489,4490
Diverticulitis|4491,4505
.|4505,4506
<EOL>|4506,4507
.|4507,4508
<EOL>|4508,4509
RADIOLOGY|4509,4518
Final|4520,4525
Report|4526,4532
<EOL>|4532,4533
CT|4533,4535
ABDOMEN|4536,4543
W|4544,4545
/|4545,4546
CONTRAST|4546,4554
_|4556,4557
_|4557,4558
_|4558,4559
10|4560,4562
:|4562,4563
22|4563,4565
AM|4566,4568
<EOL>|4568,4569
Reason|4569,4575
:|4575,4576
Rule|4577,4581
out|4582,4585
subcutaneous|4586,4598
air|4599,4602
or|4603,4605
fluid|4606,4611
.|4611,4612
IV|4613,4615
contrast|4616,4624
ONLY|4625,4629
.|4629,4630
<EOL>|4631,4632
HISTORY|4632,4639
:|4639,4640
_|4641,4642
_|4642,4643
_|4643,4644
female|4645,4651
with|4652,4656
recurrent|4657,4666
diverticulitis|4667,4681
,|4681,4682
<EOL>|4683,4684
status|4684,4690
post|4691,4695
laparoscopic|4696,4708
sigmoid|4709,4716
colectomy|4717,4726
,|4726,4727
now|4728,4731
with|4732,4736
incisional|4737,4747
<EOL>|4748,4749
erythema|4749,4757
.|4757,4758
Rule|4759,4763
out|4764,4767
subcutaneous|4768,4780
air|4781,4784
or|4785,4787
fluid|4788,4793
.|4793,4794
<EOL>|4794,4795
1.|4807,4809
Status|4810,4816
post|4817,4821
sigmoid|4822,4829
colectomy|4830,4839
with|4840,4844
a|4845,4846
small|4847,4852
amount|4853,4859
of|4860,4862
<EOL>|4863,4864
post-operative|4864,4878
free|4879,4883
intraperitoneal|4884,4899
air|4900,4903
and|4904,4907
fluid|4908,4913
within|4914,4920
the|4921,4924
<EOL>|4925,4926
pelvis|4926,4932
.|4932,4933
<EOL>|4933,4934
2.|4934,4936
Small|4937,4942
amount|4943,4949
of|4950,4952
scattered|4953,4962
subcutaneous|4963,4975
air|4976,4979
_|4980,4981
_|4981,4982
_|4982,4983
the|4984,4987
mid|4988,4991
and|4992,4995
<EOL>|4996,4997
lower|4997,5002
anterior|5003,5011
abdominal|5012,5021
wall|5022,5026
consistent|5027,5037
with|5038,5042
postsurgical|5043,5055
<EOL>|5056,5057
change|5057,5063
,|5063,5064
without|5065,5072
evidence|5073,5081
of|5082,5084
discrete|5085,5093
fluid|5094,5099
collection|5100,5110
.|5110,5111
<EOL>|5111,5112
<EOL>|5112,5113
<EOL>|5114,5115
Mrs.|5138,5142
_|5143,5144
_|5144,5145
_|5145,5146
was|5147,5150
directly|5151,5159
admitted|5160,5168
to|5169,5171
_|5172,5173
_|5173,5174
_|5174,5175
from|5176,5180
Dr.|5181,5184
_|5185,5186
_|5186,5187
_|5187,5188
<EOL>|5189,5190
office|5190,5196
with|5197,5201
persistent|5202,5212
abdominal|5213,5222
pain|5223,5227
likely|5228,5234
related|5235,5242
to|5243,5245
<EOL>|5246,5247
diverticulitis|5247,5261
flare|5262,5267
.|5267,5268
Her|5269,5272
vitals|5273,5279
signs|5280,5285
and|5286,5289
labwork|5290,5297
remained|5298,5306
<EOL>|5307,5308
stable|5308,5314
excluding|5315,5324
a|5325,5326
slightly|5327,5335
decreased|5336,5345
hematocrit|5346,5356
.|5356,5357
She|5358,5361
was|5362,5365
<EOL>|5366,5367
started|5367,5374
on|5375,5377
IV|5378,5380
Cipro|5381,5386
&|5387,5388
Flagyl|5389,5395
,|5395,5396
made|5397,5401
NPO|5402,5405
with|5406,5410
IVF|5411,5414
hydration|5415,5424
,|5424,5425
pain|5426,5430
<EOL>|5431,5432
managment|5432,5441
,|5441,5442
and|5443,5446
serial|5447,5453
abdominal|5454,5463
exams|5464,5469
.|5469,5470
<EOL>|5471,5472
.|5472,5473
<EOL>|5473,5474
HD2|5474,5477
-|5477,5478
HD7|5478,5481
-|5481,5482
She|5482,5485
underwent|5486,5495
a|5496,5497
abd|5498,5501
CT|5502,5504
scan|5505,5509
which|5510,5515
revealed|5516,5524
uncomplicated|5525,5538
<EOL>|5539,5540
diverticulitis|5540,5554
.|5554,5555
She|5556,5559
continued|5560,5569
with|5570,5574
the|5575,5578
above|5579,5584
mentioned|5585,5594
treatment|5595,5604
<EOL>|5605,5606
regimen|5606,5613
.|5613,5614
Her|5615,5618
abdominal|5619,5628
pain|5629,5633
responded|5634,5643
well|5644,5648
to|5649,5651
IV|5652,5654
Dilaudid|5655,5663
.|5663,5664
She|5665,5668
<EOL>|5669,5670
had|5670,5673
multiple|5674,5682
non-bloody|5683,5693
stools|5694,5700
.|5700,5701
She|5702,5705
continued|5706,5715
to|5716,5718
ambulate|5719,5727
<EOL>|5728,5729
without|5729,5736
difficulty|5737,5747
,|5747,5748
and|5749,5752
refused|5753,5760
SC|5761,5763
Heparing|5764,5772
injections|5773,5783
.|5783,5784
Surgical|5785,5793
<EOL>|5794,5795
options|5795,5802
were|5803,5807
discussed|5808,5817
b|5818,5819
/|5819,5820
w|5820,5821
patient|5822,5829
and|5830,5833
Dr.|5834,5837
_|5838,5839
_|5839,5840
_|5840,5841
.|5841,5842
Surgery|5843,5850
<EOL>|5851,5852
planned|5852,5859
for|5860,5863
_|5864,5865
_|5865,5866
_|5866,5867
.|5867,5868
TPN|5869,5872
&|5873,5874
PICC|5875,5879
was|5880,5883
not|5884,5887
indicated|5888,5897
.|5897,5898
She|5899,5902
was|5903,5906
<EOL>|5907,5908
started|5908,5915
on|5916,5918
Ensure|5919,5925
supplements|5926,5937
.|5937,5938
Operative|5939,5948
consent|5949,5956
,|5956,5957
labwork|5958,5965
,|5965,5966
CXR|5967,5970
,|5970,5971
<EOL>|5972,5973
&|5973,5974
EKG|5975,5978
were|5979,5983
collected|5984,5993
.|5993,5994
<EOL>|5994,5995
.|5995,5996
<EOL>|5996,5997
HD8|5997,6000
-|6000,6001
She|6001,6004
was|6005,6008
made|6009,6013
NPO|6014,6017
overnight|6018,6027
for|6028,6031
surgery|6032,6039
.|6039,6040
Continue|6041,6049
with|6050,6054
IVF|6055,6058
.|6058,6059
<EOL>|6060,6061
Surgery|6061,6068
was|6069,6072
performed|6073,6082
on|6083,6085
_|6086,6087
_|6087,6088
_|6088,6089
.|6089,6090
Her|6091,6094
operative|6095,6104
course|6105,6111
was|6112,6115
<EOL>|6116,6117
uncomplicated|6117,6130
.|6130,6131
Routinely|6132,6141
observed|6142,6150
_|6151,6152
_|6152,6153
_|6153,6154
PACU|6155,6159
,|6159,6160
and|6161,6164
transferred|6165,6176
to|6177,6179
<EOL>|6180,6181
_|6181,6182
_|6182,6183
_|6183,6184
.|6184,6185
<EOL>|6186,6187
.|6187,6188
<EOL>|6188,6189
POD1|6189,6193
-|6193,6194
Continued|6194,6203
with|6204,6208
IVF|6209,6212
,|6212,6213
NPO|6214,6217
,|6217,6218
and|6219,6222
foley|6223,6228
.|6228,6229
PCA|6230,6233
for|6234,6237
pain|6238,6242
management|6243,6253
<EOL>|6254,6255
with|6255,6259
adequate|6260,6268
relief|6269,6275
.|6275,6276
<EOL>|6277,6278
.|6278,6279
<EOL>|6279,6280
POD2|6280,6284
-|6284,6285
3|6285,6286
-|6286,6287
Reported|6287,6295
flatus|6296,6302
and|6303,6306
had|6307,6310
a|6311,6312
small|6313,6318
BM|6319,6321
.|6321,6322
Abdomen|6323,6330
appropriately|6331,6344
<EOL>|6345,6346
TTP|6346,6349
/|6349,6350
ND|6350,6352
with|6353,6357
active|6358,6364
bowel|6365,6370
sounds|6371,6377
.|6377,6378
Ffanesstial|6379,6390
incision|6391,6399
with|6400,6404
<EOL>|6405,6406
increased|6406,6415
erythema|6416,6424
extending|6425,6434
to|6435,6437
right|6438,6443
.|6443,6444
IV|6445,6447
Vancomycin|6448,6458
started|6459,6466
.|6466,6467
No|6468,6470
<EOL>|6471,6472
improvement|6472,6483
_|6484,6485
_|6485,6486
_|6486,6487
wound|6488,6493
x|6494,6495
24|6496,6498
hrs|6499,6502
.|6502,6503
Zosyn|6504,6509
added|6510,6515
to|6516,6518
regimen|6519,6526
.|6526,6527
Pain|6528,6532
<EOL>|6533,6534
medication|6534,6544
switched|6545,6553
to|6554,6556
PO|6557,6559
medication|6560,6570
.|6570,6571
_|6572,6573
_|6573,6574
_|6574,6575
pump|6576,6580
removed|6581,6588
.|6588,6589
<EOL>|6589,6590
.|6590,6591
<EOL>|6591,6592
POD4|6592,6596
-|6596,6597
5|6597,6598
-|6598,6599
Temp|6599,6603
spike|6604,6609
to|6610,6612
102.5|6613,6618
,|6618,6619
IV|6620,6622
antibiotics|6623,6634
started|6635,6642
.|6642,6643
WBC|6644,6647
spike|6648,6653
to|6654,6656
<EOL>|6657,6658
23|6658,6660
from|6661,6665
8|6666,6667
with|6668,6672
10|6673,6675
%|6675,6676
bands|6677,6682
.|6682,6683
Reports|6684,6691
of|6692,6694
persistent|6695,6705
nausea|6706,6712
-|6712,6713
zofran|6713,6719
<EOL>|6720,6721
mildly|6721,6727
effective|6728,6737
.|6737,6738
Compazine|6739,6748
added|6749,6754
to|6755,6757
regimen|6758,6765
with|6766,6770
improved|6771,6779
<EOL>|6780,6781
effects|6781,6788
.|6788,6789
IVF|6790,6793
continued|6794,6803
.|6803,6804
ID|6805,6807
team|6808,6812
consulted|6813,6822
regarding|6823,6832
antibiotic|6833,6843
<EOL>|6844,6845
regimen|6845,6852
.|6852,6853
Underwent|6854,6863
CT|6864,6866
scan|6867,6871
of|6872,6874
abd|6875,6878
with|6879,6883
no|6884,6886
significatn|6887,6898
intra-abd|6899,6908
<EOL>|6909,6910
.|6918,6919
Wound|6920,6925
opened|6926,6932
at|6933,6935
bedside|6936,6943
on|6944,6946
_|6947,6948
_|6948,6949
_|6949,6950
.|6950,6951
Cultures|6952,6960
of|6961,6963
serous|6964,6970
<EOL>|6971,6972
fluid|6972,6977
sent|6978,6982
to|6983,6985
_|6986,6987
_|6987,6988
_|6988,6989
.|6989,6990
Site|6991,6995
packed|6996,7002
with|7003,7007
w|7008,7009
-|7009,7010
d|7010,7011
dressing|7012,7020
.|7020,7021
Infectious|7022,7032
<EOL>|7033,7034
reaction|7034,7042
likely|7043,7049
r|7050,7051
/|7051,7052
t|7052,7053
GAS|7054,7057
or|7058,7060
staphylococcus|7061,7075
aureus|7076,7082
.|7082,7083
Nasal|7084,7089
swab|7090,7094
for|7095,7098
<EOL>|7099,7100
staphy|7100,7106
collected|7107,7116
&|7117,7118
sent|7119,7123
to|7124,7126
Micro|7127,7132
.|7132,7133
Clindamycin|7134,7145
IV|7146,7148
added|7149,7154
to|7155,7157
<EOL>|7158,7159
regimen|7159,7166
.|7166,7167
Cultures|7168,7176
were|7177,7181
followed|7182,7190
,|7190,7191
and|7192,7195
wound|7196,7201
checked|7202,7209
serially|7210,7218
.|7218,7219
<EOL>|7220,7221
T|7221,7222
-|7222,7223
max|7223,7226
100.7|7227,7232
.|7232,7233
Bump|7234,7238
_|7239,7240
_|7240,7241
_|7241,7242
creatinine|7243,7253
noted|7254,7259
0.6|7260,7263
to|7264,7266
1.7|7267,7270
.|7270,7271
<EOL>|7271,7272
.|7272,7273
<EOL>|7273,7274
POD6|7274,7278
-|7278,7279
wound|7279,7284
culture|7285,7292
positive|7293,7301
for|7302,7305
MSSA|7306,7310
.|7310,7311
IV|7312,7314
Nafcillin|7315,7324
added|7325,7330
with|7331,7335
<EOL>|7336,7337
continued|7337,7346
Clinda.|7347,7354
IV|7355,7357
Vanco|7358,7363
&|7364,7365
Zosyn|7366,7371
discontinued|7372,7384
.|7384,7385
CDIFF|7386,7391
cultures|7392,7400
<EOL>|7401,7402
negative|7402,7410
x|7411,7412
3.|7413,7415
Nasal|7416,7421
swab|7422,7426
for|7427,7430
Staph|7431,7436
cultured|7437,7445
collected|7446,7455
.|7455,7456
Patient|7457,7464
<EOL>|7465,7466
reports|7466,7473
nausea|7474,7480
still|7481,7486
present|7487,7494
,|7494,7495
but|7496,7499
better|7500,7506
.|7506,7507
Has|7508,7511
been|7512,7516
eating|7517,7523
small|7524,7529
<EOL>|7530,7531
amount|7531,7537
of|7538,7540
regular|7541,7548
food|7549,7553
with|7554,7558
continued|7559,7568
flatus|7569,7575
and|7576,7579
liquid|7580,7586
stool|7587,7592
<EOL>|7593,7594
production|7594,7604
.|7604,7605
Continues|7606,7615
with|7616,7620
IVF|7621,7624
due|7625,7628
to|7629,7631
elevated|7632,7640
Creatinine|7641,7651
to|7652,7654
<EOL>|7655,7656
1.9|7656,7659
.|7659,7660
Adequate|7661,7669
urine|7670,7675
output|7676,7682
.|7682,7683
Ambulating|7684,7694
independently|7695,7708
.|7708,7709
LFT|7710,7713
's|7713,7715
<EOL>|7716,7717
slightly|7717,7725
elevated|7726,7734
as|7735,7737
well|7738,7742
.|7742,7743
<EOL>|7743,7744
.|7744,7745
<EOL>|7745,7746
POD7|7746,7750
-|7750,7751
IV|7751,7753
Clindamycin|7754,7765
discontinued|7766,7778
due|7779,7782
to|7783,7785
culture|7786,7793
resistance|7794,7804
.|7804,7805
<EOL>|7806,7807
Nafcillin|7807,7816
continued|7817,7826
.|7826,7827
Patient|7828,7835
's|7835,7837
status|7838,7844
contiues|7845,7853
to|7854,7856
improve|7857,7864
.|7864,7865
<EOL>|7866,7867
Remains|7867,7874
afebrile|7875,7883
,|7883,7884
decreased|7885,7894
WBC|7895,7898
,|7898,7899
and|7900,7903
improved|7904,7912
appearance|7913,7923
of|7924,7926
<EOL>|7927,7928
wound|7928,7933
including|7934,7943
erythema|7944,7952
.|7952,7953
IVF|7954,7957
switched|7958,7966
to|7967,7969
maintenance|7970,7981
.|7981,7982
<EOL>|7982,7983
.|7983,7984
<EOL>|7984,7985
POD8|7985,7989
-|7989,7990
Nasal|7990,7995
swab|7996,8000
-|8000,8001
no|8001,8003
growth|8004,8010
.|8010,8011
Continues|8012,8021
IVF|8022,8025
&|8026,8027
Nafcillin|8028,8037
.|8037,8038
Improved|8039,8047
<EOL>|8048,8049
PO|8049,8051
intake|8052,8058
.|8058,8059
Continues|8060,8069
with|8070,8074
complaints|8075,8085
of|8086,8088
intermittent|8089,8101
nausea|8102,8108
,|8108,8109
<EOL>|8110,8111
improving|8111,8120
slowly|8121,8127
,|8127,8128
&|8129,8130
responsive|8131,8141
to|8142,8144
Compazine|8145,8154
.|8154,8155
Ambulating|8156,8166
<EOL>|8167,8168
independently|8168,8181
.|8181,8182
Remains|8183,8190
afebrile|8191,8199
.|8199,8200
<EOL>|8200,8201
<EOL>|8201,8202
POD9|8202,8206
-|8206,8207
Discharge|8207,8216
day|8217,8220
:|8220,8221
Creatinine|8222,8232
continued|8233,8242
to|8243,8245
decrease|8246,8254
.|8254,8255
Currently|8256,8265
<EOL>|8266,8267
1.4|8267,8270
.|8270,8271
Creatinine|8272,8282
level|8283,8288
will|8289,8293
be|8294,8296
collected|8297,8306
per|8307,8310
Home|8311,8315
_|8316,8317
_|8317,8318
_|8318,8319
on|8320,8322
_|8323,8324
_|8324,8325
_|8325,8326
<EOL>|8327,8328
_|8328,8329
_|8329,8330
_|8330,8331
,|8331,8332
and|8333,8336
called|8337,8343
into|8344,8348
PCP|8349,8352
/|8352,8353
Dr|8353,8355
.|8355,8356
_|8357,8358
_|8358,8359
_|8359,8360
.|8360,8361
Continued|8362,8371
to|8372,8374
<EOL>|8375,8376
tolerate|8376,8384
food|8385,8389
with|8390,8394
intermittent|8395,8407
nausea|8408,8414
,|8414,8415
improved|8416,8424
with|8425,8429
eating|8430,8436
.|8436,8437
<EOL>|8438,8439
All|8439,8442
PO|8443,8445
narcotics|8446,8455
discontinued|8456,8468
,|8468,8469
and|8470,8473
Keflex|8474,8480
switched|8481,8489
to|8490,8492
suspension|8493,8503
<EOL>|8504,8505
which|8505,8510
patient|8511,8518
was|8519,8522
better|8523,8529
able|8530,8534
to|8535,8537
tolerate|8538,8546
.|8546,8547
_|8548,8549
_|8549,8550
_|8550,8551
was|8552,8555
set|8556,8559
up|8560,8562
for|8563,8566
<EOL>|8567,8568
wound|8568,8573
care|8574,8578
.|8578,8579
<EOL>|8580,8581
<EOL>|8582,8583
Medications|8583,8594
on|8595,8597
Admission|8598,8607
:|8607,8608
<EOL>|8608,8609
Lexapro|8609,8616
10|8617,8619
,|8619,8620
nasonex|8621,8628
<EOL>|8629,8630
<EOL>|8631,8632
Discharge|8632,8641
Medications|8642,8653
:|8653,8654
<EOL>|8654,8655
1.|8655,8657
Escitalopram|8658,8670
10|8671,8673
mg|8674,8676
Tablet|8677,8683
Sig|8684,8687
:|8687,8688
One|8689,8692
(|8693,8694
1|8694,8695
)|8695,8696
Tablet|8697,8703
PO|8704,8706
DAILY|8707,8712
<EOL>|8713,8714
(|8714,8715
Daily|8715,8720
)|8720,8721
.|8721,8722
<EOL>|8724,8725
2.|8725,8727
Fluticasone|8728,8739
50|8740,8742
mcg|8743,8746
/|8746,8747
Actuation|8747,8756
Spray|8757,8762
,|8762,8763
Suspension|8764,8774
Sig|8775,8778
:|8778,8779
One|8780,8783
(|8784,8785
1|8785,8786
)|8786,8787
<EOL>|8788,8789
Spray|8789,8794
Nasal|8795,8800
DAILY|8801,8806
(|8807,8808
Daily|8808,8813
)|8813,8814
.|8814,8815
<EOL>|8817,8818
3.|8818,8820
Colace|8821,8827
100|8828,8831
mg|8832,8834
Capsule|8835,8842
Sig|8843,8846
:|8846,8847
One|8848,8851
(|8852,8853
1|8853,8854
)|8854,8855
Capsule|8856,8863
PO|8864,8866
twice|8867,8872
a|8873,8874
day|8875,8878
as|8879,8881
<EOL>|8882,8883
needed|8883,8889
for|8890,8893
constipation|8894,8906
for|8907,8910
1|8911,8912
months|8913,8919
.|8919,8920
<EOL>|8920,8921
Disp|8921,8925
:|8925,8926
*|8926,8927
60|8927,8929
Capsule|8930,8937
(|8937,8938
s|8938,8939
)|8939,8940
*|8940,8941
Refills|8942,8949
:|8949,8950
*|8950,8951
0|8951,8952
*|8952,8953
<EOL>|8953,8954
4.|8954,8956
Lorazepam|8957,8966
0.5|8967,8970
mg|8971,8973
Tablet|8974,8980
Sig|8981,8984
:|8984,8985
One|8986,8989
(|8990,8991
1|8991,8992
)|8992,8993
Tablet|8994,9000
PO|9001,9003
Q8H|9004,9007
(|9008,9009
every|9009,9014
8|9015,9016
<EOL>|9017,9018
hours|9018,9023
)|9023,9024
as|9025,9027
needed|9028,9034
for|9035,9038
anxiety|9039,9046
.|9046,9047
<EOL>|9049,9050
5.|9050,9052
Hydrocortisone|9053,9067
2.5|9068,9071
%|9072,9073
Cream|9074,9079
Sig|9080,9083
:|9083,9084
One|9085,9088
(|9089,9090
1|9090,9091
)|9091,9092
Appl|9093,9097
Rectal|9098,9104
TID|9105,9108
(|9109,9110
3|9110,9111
<EOL>|9112,9113
times|9113,9118
a|9119,9120
day|9121,9124
)|9124,9125
as|9126,9128
needed|9129,9135
for|9136,9139
hemorrhoids|9140,9151
.|9151,9152
<EOL>|9154,9155
6.|9155,9157
Cephalexin|9158,9168
250|9169,9172
mg|9173,9175
/|9175,9176
5|9176,9177
mL|9178,9180
Suspension|9181,9191
for|9192,9195
Reconstitution|9196,9210
Sig|9211,9214
:|9214,9215
Two|9216,9219
<EOL>|9220,9221
(|9221,9222
2|9222,9223
)|9223,9224
PO|9226,9228
q12hrs|9229,9235
(|9236,9237
)|9237,9238
for|9239,9242
5|9243,9244
days|9245,9249
.|9249,9250
<EOL>|9250,9251
Disp|9251,9255
:|9255,9256
*|9256,9257
qs|9257,9259
*|9260,9261
Refills|9262,9269
:|9269,9270
*|9270,9271
0|9271,9272
*|9272,9273
<EOL>|9273,9274
7.|9274,9276
Tylenol|9277,9284
_|9285,9286
_|9286,9287
_|9287,9288
mg|9289,9291
Tablet|9292,9298
Sig|9299,9302
:|9302,9303
Two|9304,9307
(|9308,9309
2|9309,9310
)|9310,9311
Tablet|9312,9318
PO|9319,9321
every|9322,9327
_|9328,9329
_|9329,9330
_|9330,9331
hours|9332,9337
<EOL>|9338,9339
as|9339,9341
needed|9342,9348
for|9349,9352
fever|9353,9358
or|9359,9361
pain|9362,9366
.|9366,9367
<EOL>|9369,9370
8.|9370,9372
Outpatient|9373,9383
Lab|9384,9387
Work|9388,9392
<EOL>|9392,9393
Please|9393,9399
check|9400,9405
serum|9406,9411
Creatinine|9412,9422
on|9423,9425
_|9426,9427
_|9427,9428
_|9428,9429
.|9429,9430
<EOL>|9430,9431
<EOL>|9431,9432
*|9432,9433
*|9433,9434
Call|9434,9438
result|9439,9445
to|9446,9448
PCP|9449,9452
and|9453,9456
Dr.|9457,9460
_|9461,9462
_|9462,9463
_|9463,9464
<EOL>|9464,9465
<EOL>|9465,9466
<EOL>|9467,9468
_|9468,9469
_|9469,9470
_|9470,9471
Disposition|9472,9483
:|9483,9484
<EOL>|9484,9485
Home|9485,9489
With|9490,9494
Service|9495,9502
<EOL>|9502,9503
<EOL>|9504,9505
Facility|9505,9513
:|9513,9514
<EOL>|9514,9515
_|9515,9516
_|9516,9517
_|9517,9518
<EOL>|9518,9519
<EOL>|9520,9521
Discharge|9521,9530
Diagnosis|9531,9540
:|9540,9541
<EOL>|9541,9542
Primary|9542,9549
:|9549,9550
<EOL>|9550,9551
Recurrent|9551,9560
Diverticulitis|9561,9575
<EOL>|9575,9576
Post-op|9576,9583
wound|9584,9589
cellulitis|9590,9600
<EOL>|9600,9601
Post-op|9601,9608
hypovolemia|9609,9620
<EOL>|9620,9621
Post-op|9621,9628
fever|9629,9634
<EOL>|9634,9635
.|9635,9636
<EOL>|9636,9637
Secondary|9637,9646
:|9646,9647
<EOL>|9647,9648
Anxiety|9648,9655
<EOL>|9655,9656
diverticulosis|9656,9670
<EOL>|9670,9671
<EOL>|9671,9672
<EOL>|9673,9674
Stable|9695,9701
<EOL>|9701,9702
Tolerating|9702,9712
a|9713,9714
regular|9715,9722
,|9722,9723
low|9724,9727
-|9727,9728
residue|9728,9735
diet|9736,9740
<EOL>|9740,9741
Adequate|9741,9749
pain|9750,9754
control|9755,9762
with|9763,9767
oral|9768,9772
medication|9773,9783
<EOL>|9783,9784
<EOL>|9784,9785
<EOL>|9786,9787
Please|9811,9817
call|9818,9822
your|9823,9827
doctor|9828,9834
or|9835,9837
return|9838,9844
to|9845,9847
the|9848,9851
ER|9852,9854
for|9855,9858
any|9859,9862
of|9863,9865
the|9866,9869
<EOL>|9870,9871
following|9871,9880
:|9880,9881
<EOL>|9881,9882
*|9882,9883
You|9884,9887
experience|9888,9898
new|9899,9902
chest|9903,9908
pain|9909,9913
,|9913,9914
pressure|9915,9923
,|9923,9924
squeezing|9925,9934
or|9935,9937
<EOL>|9938,9939
tightness|9939,9948
.|9948,9949
<EOL>|9949,9950
*|9950,9951
New|9952,9955
or|9956,9958
worsening|9959,9968
cough|9969,9974
or|9975,9977
wheezing|9978,9986
.|9986,9987
<EOL>|9987,9988
*|9988,9989
If|9990,9992
you|9993,9996
are|9997,10000
vomiting|10001,10009
and|10010,10013
can|10014,10017
not|10017,10020
keep|10021,10025
_|10026,10027
_|10027,10028
_|10028,10029
fluids|10030,10036
or|10037,10039
your|10040,10044
<EOL>|10045,10046
medications|10046,10057
.|10057,10058
<EOL>|10058,10059
*|10059,10060
You|10061,10064
are|10065,10068
getting|10069,10076
dehydrated|10077,10087
due|10088,10091
to|10092,10094
continued|10095,10104
vomiting|10105,10113
,|10113,10114
<EOL>|10115,10116
diarrhea|10116,10124
or|10125,10127
other|10128,10133
reasons|10134,10141
.|10141,10142
Signs|10143,10148
of|10149,10151
dehydration|10152,10163
include|10164,10171
dry|10172,10175
<EOL>|10176,10177
mouth|10177,10182
,|10182,10183
rapid|10184,10189
heartbeat|10190,10199
or|10200,10202
feeling|10203,10210
dizzy|10211,10216
or|10217,10219
faint|10220,10225
when|10226,10230
standing|10231,10239
.|10239,10240
<EOL>|10240,10241
*|10241,10242
You|10243,10246
see|10247,10250
blood|10251,10256
or|10257,10259
dark|10260,10264
/|10264,10265
black|10265,10270
material|10271,10279
when|10280,10284
you|10285,10288
vomit|10289,10294
or|10295,10297
have|10298,10302
a|10303,10304
<EOL>|10305,10306
bowel|10306,10311
movement|10312,10320
.|10320,10321
<EOL>|10321,10322
*|10322,10323
Your|10324,10328
pain|10329,10333
is|10334,10336
not|10337,10340
improving|10341,10350
within|10351,10357
_|10358,10359
_|10359,10360
_|10360,10361
hours|10362,10367
or|10368,10370
not|10371,10374
gone|10375,10379
<EOL>|10380,10381
within|10381,10387
24|10388,10390
hours|10391,10396
.|10396,10397
Call|10398,10402
or|10403,10405
return|10406,10412
immediately|10413,10424
if|10425,10427
your|10428,10432
pain|10433,10437
is|10438,10440
<EOL>|10441,10442
getting|10442,10449
worse|10450,10455
or|10456,10458
is|10459,10461
changing|10462,10470
location|10471,10479
or|10480,10482
moving|10483,10489
to|10490,10492
your|10493,10497
chest|10498,10503
or|10504,10506
<EOL>|10507,10508
<EOL>|10508,10509
back|10509,10513
.|10513,10514
<EOL>|10514,10515
*|10515,10516
Avoid|10516,10521
driving|10522,10529
or|10530,10532
operating|10533,10542
heavy|10543,10548
machinery|10549,10558
while|10559,10564
taking|10565,10571
pain|10572,10576
<EOL>|10577,10578
medications|10578,10589
.|10589,10590
<EOL>|10590,10591
*|10591,10592
You|10593,10596
have|10597,10601
shaking|10602,10609
chills|10610,10616
,|10616,10617
or|10618,10620
a|10621,10622
fever|10623,10628
greater|10629,10636
than|10637,10641
101.5|10642,10647
(|10648,10649
F|10649,10650
)|10650,10651
<EOL>|10652,10653
degrees|10653,10660
or|10661,10663
38|10664,10666
(|10666,10667
C|10667,10668
)|10668,10669
degrees|10670,10677
.|10677,10678
<EOL>|10678,10679
*|10679,10680
Any|10681,10684
serious|10685,10692
change|10693,10699
_|10700,10701
_|10701,10702
_|10702,10703
your|10704,10708
symptoms|10709,10717
,|10717,10718
or|10719,10721
any|10722,10725
new|10726,10729
symptoms|10730,10738
that|10739,10743
<EOL>|10744,10745
concern|10745,10752
you|10753,10756
.|10756,10757
<EOL>|10758,10759
*|10759,10760
Please|10761,10767
resume|10768,10774
all|10775,10778
regular|10779,10786
home|10787,10791
medications|10792,10803
and|10804,10807
take|10808,10812
any|10813,10816
new|10817,10820
<EOL>|10821,10822
meds|10822,10826
<EOL>|10827,10828
as|10828,10830
ordered|10831,10838
.|10838,10839
<EOL>|10840,10841
*|10841,10842
Continue|10843,10851
to|10852,10854
ambulate|10855,10863
several|10864,10871
times|10872,10877
per|10878,10881
day|10882,10885
.|10885,10886
<EOL>|10886,10887
.|10887,10888
<EOL>|10888,10889
WOUND|10889,10894
CARE|10895,10899
:|10899,10900
<EOL>|10900,10901
*|10901,10902
Assess|10902,10908
surgical|10909,10917
wound|10918,10923
site|10924,10928
daily|10929,10934
.|10934,10935
<EOL>|10935,10936
*|10936,10937
Change|10937,10943
packing|10944,10951
at|10952,10954
least|10955,10960
once|10961,10965
per|10966,10969
day|10970,10973
,|10973,10974
and|10975,10978
as|10979,10981
needed|10982,10988
.|10988,10989
<EOL>|10989,10990
*|10990,10991
Pack|10991,10995
with|10996,11000
moistened|11001,11010
gauze|11011,11016
(|11017,11018
Normal|11018,11024
Saline|11025,11031
)|11031,11032
into|11033,11037
incisional|11038,11048
<EOL>|11049,11050
cavity|11050,11056
.|11056,11057
Apply|11058,11063
dry|11064,11067
gauze|11068,11073
on|11074,11076
top|11077,11080
,|11080,11081
and|11082,11085
adhere|11086,11092
with|11093,11097
paper|11098,11103
tape|11104,11108
.|11108,11109
<EOL>|11109,11110
*|11110,11111
*|11111,11112
Changed|11112,11119
top|11120,11123
(|11124,11125
dry|11125,11128
gauze|11129,11134
)|11134,11135
if|11136,11138
saturated|11139,11148
to|11149,11151
prevent|11152,11159
irritation|11160,11170
to|11171,11173
<EOL>|11174,11175
surrounding|11175,11186
skin|11187,11191
.|11191,11192
<EOL>|11192,11193
*|11193,11194
*|11194,11195
If|11195,11197
wound|11198,11203
continues|11204,11213
to|11214,11216
weep|11217,11221
,|11221,11222
pack|11223,11227
with|11228,11232
Aquacel|11234,11241
or|11242,11244
DSD|11245,11248
.|11248,11249
<EOL>|11249,11250
-|11250,11251
You|11251,11254
may|11255,11258
shower|11259,11265
briefly|11266,11273
,|11273,11274
and|11275,11278
wash|11279,11283
around|11284,11290
surgical|11291,11299
incisions|11300,11309
.|11309,11310
<EOL>|11310,11311
-|11311,11312
Avoid|11312,11317
swimming|11318,11326
and|11327,11330
tub|11331,11334
baths|11335,11340
until|11341,11346
wound|11347,11352
completely|11353,11363
healed|11364,11370
<EOL>|11370,11371
-|11371,11372
Please|11372,11378
call|11379,11383
the|11384,11387
doctor|11388,11394
if|11395,11397
you|11398,11401
have|11402,11406
increased|11407,11416
pain|11417,11421
,|11421,11422
swelling|11423,11431
,|11431,11432
<EOL>|11433,11434
redness|11434,11441
,|11441,11442
or|11443,11445
drainage|11446,11454
from|11455,11459
the|11460,11463
incision|11464,11472
sites|11473,11478
.|11478,11479
<EOL>|11479,11480
.|11480,11481
<EOL>|11481,11482
CREATININE|11482,11492
:|11492,11493
<EOL>|11493,11494
*|11494,11495
Please|11495,11501
have|11502,11506
the|11507,11510
_|11511,11512
_|11512,11513
_|11513,11514
check|11515,11520
your|11521,11525
creatinine|11526,11536
on|11537,11539
_|11540,11541
_|11541,11542
_|11542,11543
.|11543,11544
Please|11545,11551
<EOL>|11552,11553
call|11553,11557
Dr.|11558,11561
_|11562,11563
_|11563,11564
_|11564,11565
and|11566,11569
/|11569,11570
or|11570,11572
your|11573,11577
PCP|11578,11581
's|11581,11583
office|11584,11590
with|11591,11595
the|11596,11599
<EOL>|11600,11601
result|11601,11607
.|11607,11608
<EOL>|11608,11609
<EOL>|11609,11610
<EOL>|11611,11612
Followup|11612,11620
Instructions|11621,11633
:|11633,11634
<EOL>|11634,11635
_|11635,11636
_|11636,11637
_|11637,11638
<EOL>|11638,11639

